library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LUT is
port (
	address : in integer range 0 to 65535;
	data_val : out std_logic_vector(15 downto 0)
	);
end LUT;

architecture archLUT of LUT is
	type lut_array is array (0 to 65535) of std_logic_vector(15 downto 0);
   constant lut_data : lut_array := (
0 => "0000000000010101",
1 => "0000000000010101",
2 => "0000000000010101",
3 => "0000000000010101",
4 => "0000000000010101",
5 => "0000000000010110",
6 => "0000000000010110",
7 => "0000000000010110",
8 => "0000000000010110",
9 => "0000000000010110",
10 => "0000000000010110",
11 => "0000000000010110",
12 => "0000000000010110",
13 => "0000000000010110",
14 => "0000000000010110",
15 => "0000000000010110",
16 => "0000000000010110",
17 => "0000000000010110",
18 => "0000000000010110",
19 => "0000000000010110",
20 => "0000000000010110",
21 => "0000000000010110",
22 => "0000000000010110",
23 => "0000000000010110",
24 => "0000000000010110",
25 => "0000000000010110",
26 => "0000000000010110",
27 => "0000000000010110",
28 => "0000000000010110",
29 => "0000000000010110",
30 => "0000000000010110",
31 => "0000000000010110",
32 => "0000000000010110",
33 => "0000000000010110",
34 => "0000000000010110",
35 => "0000000000010110",
36 => "0000000000010110",
37 => "0000000000010110",
38 => "0000000000010110",
39 => "0000000000010110",
40 => "0000000000010110",
41 => "0000000000010110",
42 => "0000000000010110",
43 => "0000000000010110",
44 => "0000000000010110",
45 => "0000000000010110",
46 => "0000000000010110",
47 => "0000000000010110",
48 => "0000000000010110",
49 => "0000000000010110",
50 => "0000000000010110",
51 => "0000000000010110",
52 => "0000000000010110",
53 => "0000000000010110",
54 => "0000000000010110",
55 => "0000000000010110",
56 => "0000000000010110",
57 => "0000000000010110",
58 => "0000000000010110",
59 => "0000000000010110",
60 => "0000000000010110",
61 => "0000000000010110",
62 => "0000000000010110",
63 => "0000000000010110",
64 => "0000000000010110",
65 => "0000000000010110",
66 => "0000000000010110",
67 => "0000000000010110",
68 => "0000000000010110",
69 => "0000000000010110",
70 => "0000000000010110",
71 => "0000000000010110",
72 => "0000000000010110",
73 => "0000000000010110",
74 => "0000000000010110",
75 => "0000000000010110",
76 => "0000000000010110",
77 => "0000000000010110",
78 => "0000000000010110",
79 => "0000000000010110",
80 => "0000000000010110",
81 => "0000000000010110",
82 => "0000000000010110",
83 => "0000000000010110",
84 => "0000000000010110",
85 => "0000000000010110",
86 => "0000000000010110",
87 => "0000000000010110",
88 => "0000000000010110",
89 => "0000000000010110",
90 => "0000000000010110",
91 => "0000000000010110",
92 => "0000000000010110",
93 => "0000000000010110",
94 => "0000000000010110",
95 => "0000000000010110",
96 => "0000000000010110",
97 => "0000000000010110",
98 => "0000000000010110",
99 => "0000000000010110",
100 => "0000000000010110",
101 => "0000000000010110",
102 => "0000000000010110",
103 => "0000000000010110",
104 => "0000000000010110",
105 => "0000000000010110",
106 => "0000000000010110",
107 => "0000000000010110",
108 => "0000000000010110",
109 => "0000000000010110",
110 => "0000000000010110",
111 => "0000000000010110",
112 => "0000000000010110",
113 => "0000000000010110",
114 => "0000000000010110",
115 => "0000000000010110",
116 => "0000000000010110",
117 => "0000000000010110",
118 => "0000000000010110",
119 => "0000000000010110",
120 => "0000000000010110",
121 => "0000000000010110",
122 => "0000000000010110",
123 => "0000000000010110",
124 => "0000000000010110",
125 => "0000000000010110",
126 => "0000000000010110",
127 => "0000000000010110",
128 => "0000000000010110",
129 => "0000000000010110",
130 => "0000000000010110",
131 => "0000000000010110",
132 => "0000000000010110",
133 => "0000000000010110",
134 => "0000000000010110",
135 => "0000000000010110",
136 => "0000000000010110",
137 => "0000000000010110",
138 => "0000000000010110",
139 => "0000000000010110",
140 => "0000000000010110",
141 => "0000000000010110",
142 => "0000000000010110",
143 => "0000000000010110",
144 => "0000000000010110",
145 => "0000000000010110",
146 => "0000000000010110",
147 => "0000000000010110",
148 => "0000000000010110",
149 => "0000000000010110",
150 => "0000000000010110",
151 => "0000000000010110",
152 => "0000000000010110",
153 => "0000000000010110",
154 => "0000000000010110",
155 => "0000000000010110",
156 => "0000000000010110",
157 => "0000000000010110",
158 => "0000000000010110",
159 => "0000000000010110",
160 => "0000000000010110",
161 => "0000000000010110",
162 => "0000000000010110",
163 => "0000000000010110",
164 => "0000000000010110",
165 => "0000000000010110",
166 => "0000000000010110",
167 => "0000000000010110",
168 => "0000000000010110",
169 => "0000000000010110",
170 => "0000000000010110",
171 => "0000000000010110",
172 => "0000000000010110",
173 => "0000000000010110",
174 => "0000000000010110",
175 => "0000000000010110",
176 => "0000000000010110",
177 => "0000000000010110",
178 => "0000000000010110",
179 => "0000000000010110",
180 => "0000000000010110",
181 => "0000000000010110",
182 => "0000000000010110",
183 => "0000000000010110",
184 => "0000000000010110",
185 => "0000000000010110",
186 => "0000000000010110",
187 => "0000000000010111",
188 => "0000000000010111",
189 => "0000000000010111",
190 => "0000000000010111",
191 => "0000000000010111",
192 => "0000000000010111",
193 => "0000000000010111",
194 => "0000000000010111",
195 => "0000000000010111",
196 => "0000000000010111",
197 => "0000000000010111",
198 => "0000000000010111",
199 => "0000000000010111",
200 => "0000000000010111",
201 => "0000000000010111",
202 => "0000000000010111",
203 => "0000000000010111",
204 => "0000000000010111",
205 => "0000000000010111",
206 => "0000000000010111",
207 => "0000000000010111",
208 => "0000000000010111",
209 => "0000000000010111",
210 => "0000000000010111",
211 => "0000000000010111",
212 => "0000000000010111",
213 => "0000000000010111",
214 => "0000000000010111",
215 => "0000000000010111",
216 => "0000000000010111",
217 => "0000000000010111",
218 => "0000000000010111",
219 => "0000000000010111",
220 => "0000000000010111",
221 => "0000000000010111",
222 => "0000000000010111",
223 => "0000000000010111",
224 => "0000000000010111",
225 => "0000000000010111",
226 => "0000000000010111",
227 => "0000000000010111",
228 => "0000000000010111",
229 => "0000000000010111",
230 => "0000000000010111",
231 => "0000000000010111",
232 => "0000000000010111",
233 => "0000000000010111",
234 => "0000000000010111",
235 => "0000000000010111",
236 => "0000000000010111",
237 => "0000000000010111",
238 => "0000000000010111",
239 => "0000000000010111",
240 => "0000000000010111",
241 => "0000000000010111",
242 => "0000000000010111",
243 => "0000000000010111",
244 => "0000000000010111",
245 => "0000000000010111",
246 => "0000000000010111",
247 => "0000000000010111",
248 => "0000000000010111",
249 => "0000000000010111",
250 => "0000000000010111",
251 => "0000000000010111",
252 => "0000000000010111",
253 => "0000000000010111",
254 => "0000000000010111",
255 => "0000000000010111",
256 => "0000000000010111",
257 => "0000000000010111",
258 => "0000000000010111",
259 => "0000000000010111",
260 => "0000000000010111",
261 => "0000000000010111",
262 => "0000000000010111",
263 => "0000000000010111",
264 => "0000000000010111",
265 => "0000000000010111",
266 => "0000000000010111",
267 => "0000000000010111",
268 => "0000000000010111",
269 => "0000000000010111",
270 => "0000000000010111",
271 => "0000000000010111",
272 => "0000000000010111",
273 => "0000000000010111",
274 => "0000000000010111",
275 => "0000000000010111",
276 => "0000000000010111",
277 => "0000000000010111",
278 => "0000000000010111",
279 => "0000000000010111",
280 => "0000000000010111",
281 => "0000000000010111",
282 => "0000000000010111",
283 => "0000000000010111",
284 => "0000000000010111",
285 => "0000000000010111",
286 => "0000000000010111",
287 => "0000000000010111",
288 => "0000000000010111",
289 => "0000000000010111",
290 => "0000000000010111",
291 => "0000000000010111",
292 => "0000000000010111",
293 => "0000000000010111",
294 => "0000000000010111",
295 => "0000000000010111",
296 => "0000000000010111",
297 => "0000000000010111",
298 => "0000000000010111",
299 => "0000000000010111",
300 => "0000000000010111",
301 => "0000000000010111",
302 => "0000000000010111",
303 => "0000000000010111",
304 => "0000000000010111",
305 => "0000000000010111",
306 => "0000000000010111",
307 => "0000000000010111",
308 => "0000000000010111",
309 => "0000000000010111",
310 => "0000000000010111",
311 => "0000000000010111",
312 => "0000000000010111",
313 => "0000000000010111",
314 => "0000000000010111",
315 => "0000000000010111",
316 => "0000000000010111",
317 => "0000000000010111",
318 => "0000000000010111",
319 => "0000000000010111",
320 => "0000000000010111",
321 => "0000000000010111",
322 => "0000000000010111",
323 => "0000000000010111",
324 => "0000000000010111",
325 => "0000000000010111",
326 => "0000000000010111",
327 => "0000000000010111",
328 => "0000000000010111",
329 => "0000000000010111",
330 => "0000000000010111",
331 => "0000000000010111",
332 => "0000000000010111",
333 => "0000000000010111",
334 => "0000000000010111",
335 => "0000000000010111",
336 => "0000000000010111",
337 => "0000000000010111",
338 => "0000000000010111",
339 => "0000000000010111",
340 => "0000000000010111",
341 => "0000000000010111",
342 => "0000000000010111",
343 => "0000000000010111",
344 => "0000000000010111",
345 => "0000000000010111",
346 => "0000000000010111",
347 => "0000000000010111",
348 => "0000000000010111",
349 => "0000000000010111",
350 => "0000000000010111",
351 => "0000000000010111",
352 => "0000000000010111",
353 => "0000000000010111",
354 => "0000000000010111",
355 => "0000000000010111",
356 => "0000000000010111",
357 => "0000000000010111",
358 => "0000000000010111",
359 => "0000000000010111",
360 => "0000000000010111",
361 => "0000000000011000",
362 => "0000000000011000",
363 => "0000000000011000",
364 => "0000000000011000",
365 => "0000000000011000",
366 => "0000000000011000",
367 => "0000000000011000",
368 => "0000000000011000",
369 => "0000000000011000",
370 => "0000000000011000",
371 => "0000000000011000",
372 => "0000000000011000",
373 => "0000000000011000",
374 => "0000000000011000",
375 => "0000000000011000",
376 => "0000000000011000",
377 => "0000000000011000",
378 => "0000000000011000",
379 => "0000000000011000",
380 => "0000000000011000",
381 => "0000000000011000",
382 => "0000000000011000",
383 => "0000000000011000",
384 => "0000000000011000",
385 => "0000000000011000",
386 => "0000000000011000",
387 => "0000000000011000",
388 => "0000000000011000",
389 => "0000000000011000",
390 => "0000000000011000",
391 => "0000000000011000",
392 => "0000000000011000",
393 => "0000000000011000",
394 => "0000000000011000",
395 => "0000000000011000",
396 => "0000000000011000",
397 => "0000000000011000",
398 => "0000000000011000",
399 => "0000000000011000",
400 => "0000000000011000",
401 => "0000000000011000",
402 => "0000000000011000",
403 => "0000000000011000",
404 => "0000000000011000",
405 => "0000000000011000",
406 => "0000000000011000",
407 => "0000000000011000",
408 => "0000000000011000",
409 => "0000000000011000",
410 => "0000000000011000",
411 => "0000000000011000",
412 => "0000000000011000",
413 => "0000000000011000",
414 => "0000000000011000",
415 => "0000000000011000",
416 => "0000000000011000",
417 => "0000000000011000",
418 => "0000000000011000",
419 => "0000000000011000",
420 => "0000000000011000",
421 => "0000000000011000",
422 => "0000000000011000",
423 => "0000000000011000",
424 => "0000000000011000",
425 => "0000000000011000",
426 => "0000000000011000",
427 => "0000000000011000",
428 => "0000000000011000",
429 => "0000000000011000",
430 => "0000000000011000",
431 => "0000000000011000",
432 => "0000000000011000",
433 => "0000000000011000",
434 => "0000000000011000",
435 => "0000000000011000",
436 => "0000000000011000",
437 => "0000000000011000",
438 => "0000000000011000",
439 => "0000000000011000",
440 => "0000000000011000",
441 => "0000000000011000",
442 => "0000000000011000",
443 => "0000000000011000",
444 => "0000000000011000",
445 => "0000000000011000",
446 => "0000000000011000",
447 => "0000000000011000",
448 => "0000000000011000",
449 => "0000000000011000",
450 => "0000000000011000",
451 => "0000000000011000",
452 => "0000000000011000",
453 => "0000000000011000",
454 => "0000000000011000",
455 => "0000000000011000",
456 => "0000000000011000",
457 => "0000000000011000",
458 => "0000000000011000",
459 => "0000000000011000",
460 => "0000000000011000",
461 => "0000000000011000",
462 => "0000000000011000",
463 => "0000000000011000",
464 => "0000000000011000",
465 => "0000000000011000",
466 => "0000000000011000",
467 => "0000000000011000",
468 => "0000000000011000",
469 => "0000000000011000",
470 => "0000000000011000",
471 => "0000000000011000",
472 => "0000000000011000",
473 => "0000000000011000",
474 => "0000000000011000",
475 => "0000000000011000",
476 => "0000000000011000",
477 => "0000000000011000",
478 => "0000000000011000",
479 => "0000000000011000",
480 => "0000000000011000",
481 => "0000000000011000",
482 => "0000000000011000",
483 => "0000000000011000",
484 => "0000000000011000",
485 => "0000000000011000",
486 => "0000000000011000",
487 => "0000000000011000",
488 => "0000000000011000",
489 => "0000000000011000",
490 => "0000000000011000",
491 => "0000000000011000",
492 => "0000000000011000",
493 => "0000000000011000",
494 => "0000000000011000",
495 => "0000000000011000",
496 => "0000000000011000",
497 => "0000000000011000",
498 => "0000000000011000",
499 => "0000000000011000",
500 => "0000000000011000",
501 => "0000000000011000",
502 => "0000000000011000",
503 => "0000000000011000",
504 => "0000000000011000",
505 => "0000000000011000",
506 => "0000000000011000",
507 => "0000000000011000",
508 => "0000000000011000",
509 => "0000000000011000",
510 => "0000000000011000",
511 => "0000000000011000",
512 => "0000000000011000",
513 => "0000000000011000",
514 => "0000000000011000",
515 => "0000000000011000",
516 => "0000000000011000",
517 => "0000000000011000",
518 => "0000000000011000",
519 => "0000000000011000",
520 => "0000000000011000",
521 => "0000000000011000",
522 => "0000000000011000",
523 => "0000000000011000",
524 => "0000000000011000",
525 => "0000000000011000",
526 => "0000000000011000",
527 => "0000000000011000",
528 => "0000000000011001",
529 => "0000000000011001",
530 => "0000000000011001",
531 => "0000000000011001",
532 => "0000000000011001",
533 => "0000000000011001",
534 => "0000000000011001",
535 => "0000000000011001",
536 => "0000000000011001",
537 => "0000000000011001",
538 => "0000000000011001",
539 => "0000000000011001",
540 => "0000000000011001",
541 => "0000000000011001",
542 => "0000000000011001",
543 => "0000000000011001",
544 => "0000000000011001",
545 => "0000000000011001",
546 => "0000000000011001",
547 => "0000000000011001",
548 => "0000000000011001",
549 => "0000000000011001",
550 => "0000000000011001",
551 => "0000000000011001",
552 => "0000000000011001",
553 => "0000000000011001",
554 => "0000000000011001",
555 => "0000000000011001",
556 => "0000000000011001",
557 => "0000000000011001",
558 => "0000000000011001",
559 => "0000000000011001",
560 => "0000000000011001",
561 => "0000000000011001",
562 => "0000000000011001",
563 => "0000000000011001",
564 => "0000000000011001",
565 => "0000000000011001",
566 => "0000000000011001",
567 => "0000000000011001",
568 => "0000000000011001",
569 => "0000000000011001",
570 => "0000000000011001",
571 => "0000000000011001",
572 => "0000000000011001",
573 => "0000000000011001",
574 => "0000000000011001",
575 => "0000000000011001",
576 => "0000000000011001",
577 => "0000000000011001",
578 => "0000000000011001",
579 => "0000000000011001",
580 => "0000000000011001",
581 => "0000000000011001",
582 => "0000000000011001",
583 => "0000000000011001",
584 => "0000000000011001",
585 => "0000000000011001",
586 => "0000000000011001",
587 => "0000000000011001",
588 => "0000000000011001",
589 => "0000000000011001",
590 => "0000000000011001",
591 => "0000000000011001",
592 => "0000000000011001",
593 => "0000000000011001",
594 => "0000000000011001",
595 => "0000000000011001",
596 => "0000000000011001",
597 => "0000000000011001",
598 => "0000000000011001",
599 => "0000000000011001",
600 => "0000000000011001",
601 => "0000000000011001",
602 => "0000000000011001",
603 => "0000000000011001",
604 => "0000000000011001",
605 => "0000000000011001",
606 => "0000000000011001",
607 => "0000000000011001",
608 => "0000000000011001",
609 => "0000000000011001",
610 => "0000000000011001",
611 => "0000000000011001",
612 => "0000000000011001",
613 => "0000000000011001",
614 => "0000000000011001",
615 => "0000000000011001",
616 => "0000000000011001",
617 => "0000000000011001",
618 => "0000000000011001",
619 => "0000000000011001",
620 => "0000000000011001",
621 => "0000000000011001",
622 => "0000000000011001",
623 => "0000000000011001",
624 => "0000000000011001",
625 => "0000000000011001",
626 => "0000000000011001",
627 => "0000000000011001",
628 => "0000000000011001",
629 => "0000000000011001",
630 => "0000000000011001",
631 => "0000000000011001",
632 => "0000000000011001",
633 => "0000000000011001",
634 => "0000000000011001",
635 => "0000000000011001",
636 => "0000000000011001",
637 => "0000000000011001",
638 => "0000000000011001",
639 => "0000000000011001",
640 => "0000000000011001",
641 => "0000000000011001",
642 => "0000000000011001",
643 => "0000000000011001",
644 => "0000000000011001",
645 => "0000000000011001",
646 => "0000000000011001",
647 => "0000000000011001",
648 => "0000000000011001",
649 => "0000000000011001",
650 => "0000000000011001",
651 => "0000000000011001",
652 => "0000000000011001",
653 => "0000000000011001",
654 => "0000000000011001",
655 => "0000000000011001",
656 => "0000000000011001",
657 => "0000000000011001",
658 => "0000000000011001",
659 => "0000000000011001",
660 => "0000000000011001",
661 => "0000000000011001",
662 => "0000000000011001",
663 => "0000000000011001",
664 => "0000000000011001",
665 => "0000000000011001",
666 => "0000000000011001",
667 => "0000000000011001",
668 => "0000000000011001",
669 => "0000000000011001",
670 => "0000000000011001",
671 => "0000000000011001",
672 => "0000000000011001",
673 => "0000000000011001",
674 => "0000000000011001",
675 => "0000000000011001",
676 => "0000000000011001",
677 => "0000000000011001",
678 => "0000000000011001",
679 => "0000000000011001",
680 => "0000000000011001",
681 => "0000000000011001",
682 => "0000000000011001",
683 => "0000000000011001",
684 => "0000000000011001",
685 => "0000000000011001",
686 => "0000000000011001",
687 => "0000000000011001",
688 => "0000000000011001",
689 => "0000000000011010",
690 => "0000000000011010",
691 => "0000000000011010",
692 => "0000000000011010",
693 => "0000000000011010",
694 => "0000000000011010",
695 => "0000000000011010",
696 => "0000000000011010",
697 => "0000000000011010",
698 => "0000000000011010",
699 => "0000000000011010",
700 => "0000000000011010",
701 => "0000000000011010",
702 => "0000000000011010",
703 => "0000000000011010",
704 => "0000000000011010",
705 => "0000000000011010",
706 => "0000000000011010",
707 => "0000000000011010",
708 => "0000000000011010",
709 => "0000000000011010",
710 => "0000000000011010",
711 => "0000000000011010",
712 => "0000000000011010",
713 => "0000000000011010",
714 => "0000000000011010",
715 => "0000000000011010",
716 => "0000000000011010",
717 => "0000000000011010",
718 => "0000000000011010",
719 => "0000000000011010",
720 => "0000000000011010",
721 => "0000000000011010",
722 => "0000000000011010",
723 => "0000000000011010",
724 => "0000000000011010",
725 => "0000000000011010",
726 => "0000000000011010",
727 => "0000000000011010",
728 => "0000000000011010",
729 => "0000000000011010",
730 => "0000000000011010",
731 => "0000000000011010",
732 => "0000000000011010",
733 => "0000000000011010",
734 => "0000000000011010",
735 => "0000000000011010",
736 => "0000000000011010",
737 => "0000000000011010",
738 => "0000000000011010",
739 => "0000000000011010",
740 => "0000000000011010",
741 => "0000000000011010",
742 => "0000000000011010",
743 => "0000000000011010",
744 => "0000000000011010",
745 => "0000000000011010",
746 => "0000000000011010",
747 => "0000000000011010",
748 => "0000000000011010",
749 => "0000000000011010",
750 => "0000000000011010",
751 => "0000000000011010",
752 => "0000000000011010",
753 => "0000000000011010",
754 => "0000000000011010",
755 => "0000000000011010",
756 => "0000000000011010",
757 => "0000000000011010",
758 => "0000000000011010",
759 => "0000000000011010",
760 => "0000000000011010",
761 => "0000000000011010",
762 => "0000000000011010",
763 => "0000000000011010",
764 => "0000000000011010",
765 => "0000000000011010",
766 => "0000000000011010",
767 => "0000000000011010",
768 => "0000000000011010",
769 => "0000000000011010",
770 => "0000000000011010",
771 => "0000000000011010",
772 => "0000000000011010",
773 => "0000000000011010",
774 => "0000000000011010",
775 => "0000000000011010",
776 => "0000000000011010",
777 => "0000000000011010",
778 => "0000000000011010",
779 => "0000000000011010",
780 => "0000000000011010",
781 => "0000000000011010",
782 => "0000000000011010",
783 => "0000000000011010",
784 => "0000000000011010",
785 => "0000000000011010",
786 => "0000000000011010",
787 => "0000000000011010",
788 => "0000000000011010",
789 => "0000000000011010",
790 => "0000000000011010",
791 => "0000000000011010",
792 => "0000000000011010",
793 => "0000000000011010",
794 => "0000000000011010",
795 => "0000000000011010",
796 => "0000000000011010",
797 => "0000000000011010",
798 => "0000000000011010",
799 => "0000000000011010",
800 => "0000000000011010",
801 => "0000000000011010",
802 => "0000000000011010",
803 => "0000000000011010",
804 => "0000000000011010",
805 => "0000000000011010",
806 => "0000000000011010",
807 => "0000000000011010",
808 => "0000000000011010",
809 => "0000000000011010",
810 => "0000000000011010",
811 => "0000000000011010",
812 => "0000000000011010",
813 => "0000000000011010",
814 => "0000000000011010",
815 => "0000000000011010",
816 => "0000000000011010",
817 => "0000000000011010",
818 => "0000000000011010",
819 => "0000000000011010",
820 => "0000000000011010",
821 => "0000000000011010",
822 => "0000000000011010",
823 => "0000000000011010",
824 => "0000000000011010",
825 => "0000000000011010",
826 => "0000000000011010",
827 => "0000000000011010",
828 => "0000000000011010",
829 => "0000000000011010",
830 => "0000000000011010",
831 => "0000000000011010",
832 => "0000000000011010",
833 => "0000000000011010",
834 => "0000000000011010",
835 => "0000000000011010",
836 => "0000000000011010",
837 => "0000000000011010",
838 => "0000000000011010",
839 => "0000000000011010",
840 => "0000000000011010",
841 => "0000000000011010",
842 => "0000000000011010",
843 => "0000000000011010",
844 => "0000000000011011",
845 => "0000000000011011",
846 => "0000000000011011",
847 => "0000000000011011",
848 => "0000000000011011",
849 => "0000000000011011",
850 => "0000000000011011",
851 => "0000000000011011",
852 => "0000000000011011",
853 => "0000000000011011",
854 => "0000000000011011",
855 => "0000000000011011",
856 => "0000000000011011",
857 => "0000000000011011",
858 => "0000000000011011",
859 => "0000000000011011",
860 => "0000000000011011",
861 => "0000000000011011",
862 => "0000000000011011",
863 => "0000000000011011",
864 => "0000000000011011",
865 => "0000000000011011",
866 => "0000000000011011",
867 => "0000000000011011",
868 => "0000000000011011",
869 => "0000000000011011",
870 => "0000000000011011",
871 => "0000000000011011",
872 => "0000000000011011",
873 => "0000000000011011",
874 => "0000000000011011",
875 => "0000000000011011",
876 => "0000000000011011",
877 => "0000000000011011",
878 => "0000000000011011",
879 => "0000000000011011",
880 => "0000000000011011",
881 => "0000000000011011",
882 => "0000000000011011",
883 => "0000000000011011",
884 => "0000000000011011",
885 => "0000000000011011",
886 => "0000000000011011",
887 => "0000000000011011",
888 => "0000000000011011",
889 => "0000000000011011",
890 => "0000000000011011",
891 => "0000000000011011",
892 => "0000000000011011",
893 => "0000000000011011",
894 => "0000000000011011",
895 => "0000000000011011",
896 => "0000000000011011",
897 => "0000000000011011",
898 => "0000000000011011",
899 => "0000000000011011",
900 => "0000000000011011",
901 => "0000000000011011",
902 => "0000000000011011",
903 => "0000000000011011",
904 => "0000000000011011",
905 => "0000000000011011",
906 => "0000000000011011",
907 => "0000000000011011",
908 => "0000000000011011",
909 => "0000000000011011",
910 => "0000000000011011",
911 => "0000000000011011",
912 => "0000000000011011",
913 => "0000000000011011",
914 => "0000000000011011",
915 => "0000000000011011",
916 => "0000000000011011",
917 => "0000000000011011",
918 => "0000000000011011",
919 => "0000000000011011",
920 => "0000000000011011",
921 => "0000000000011011",
922 => "0000000000011011",
923 => "0000000000011011",
924 => "0000000000011011",
925 => "0000000000011011",
926 => "0000000000011011",
927 => "0000000000011011",
928 => "0000000000011011",
929 => "0000000000011011",
930 => "0000000000011011",
931 => "0000000000011011",
932 => "0000000000011011",
933 => "0000000000011011",
934 => "0000000000011011",
935 => "0000000000011011",
936 => "0000000000011011",
937 => "0000000000011011",
938 => "0000000000011011",
939 => "0000000000011011",
940 => "0000000000011011",
941 => "0000000000011011",
942 => "0000000000011011",
943 => "0000000000011011",
944 => "0000000000011011",
945 => "0000000000011011",
946 => "0000000000011011",
947 => "0000000000011011",
948 => "0000000000011011",
949 => "0000000000011011",
950 => "0000000000011011",
951 => "0000000000011011",
952 => "0000000000011011",
953 => "0000000000011011",
954 => "0000000000011011",
955 => "0000000000011011",
956 => "0000000000011011",
957 => "0000000000011011",
958 => "0000000000011011",
959 => "0000000000011011",
960 => "0000000000011011",
961 => "0000000000011011",
962 => "0000000000011011",
963 => "0000000000011011",
964 => "0000000000011011",
965 => "0000000000011011",
966 => "0000000000011011",
967 => "0000000000011011",
968 => "0000000000011011",
969 => "0000000000011011",
970 => "0000000000011011",
971 => "0000000000011011",
972 => "0000000000011011",
973 => "0000000000011011",
974 => "0000000000011011",
975 => "0000000000011011",
976 => "0000000000011011",
977 => "0000000000011011",
978 => "0000000000011011",
979 => "0000000000011011",
980 => "0000000000011011",
981 => "0000000000011011",
982 => "0000000000011011",
983 => "0000000000011011",
984 => "0000000000011011",
985 => "0000000000011011",
986 => "0000000000011011",
987 => "0000000000011011",
988 => "0000000000011011",
989 => "0000000000011011",
990 => "0000000000011011",
991 => "0000000000011011",
992 => "0000000000011011",
993 => "0000000000011100",
994 => "0000000000011100",
995 => "0000000000011100",
996 => "0000000000011100",
997 => "0000000000011100",
998 => "0000000000011100",
999 => "0000000000011100",
1000 => "0000000000011100",
1001 => "0000000000011100",
1002 => "0000000000011100",
1003 => "0000000000011100",
1004 => "0000000000011100",
1005 => "0000000000011100",
1006 => "0000000000011100",
1007 => "0000000000011100",
1008 => "0000000000011100",
1009 => "0000000000011100",
1010 => "0000000000011100",
1011 => "0000000000011100",
1012 => "0000000000011100",
1013 => "0000000000011100",
1014 => "0000000000011100",
1015 => "0000000000011100",
1016 => "0000000000011100",
1017 => "0000000000011100",
1018 => "0000000000011100",
1019 => "0000000000011100",
1020 => "0000000000011100",
1021 => "0000000000011100",
1022 => "0000000000011100",
1023 => "0000000000011100",
1024 => "0000000000011100",
1025 => "0000000000011100",
1026 => "0000000000011100",
1027 => "0000000000011100",
1028 => "0000000000011100",
1029 => "0000000000011100",
1030 => "0000000000011100",
1031 => "0000000000011100",
1032 => "0000000000011100",
1033 => "0000000000011100",
1034 => "0000000000011100",
1035 => "0000000000011100",
1036 => "0000000000011100",
1037 => "0000000000011100",
1038 => "0000000000011100",
1039 => "0000000000011100",
1040 => "0000000000011100",
1041 => "0000000000011100",
1042 => "0000000000011100",
1043 => "0000000000011100",
1044 => "0000000000011100",
1045 => "0000000000011100",
1046 => "0000000000011100",
1047 => "0000000000011100",
1048 => "0000000000011100",
1049 => "0000000000011100",
1050 => "0000000000011100",
1051 => "0000000000011100",
1052 => "0000000000011100",
1053 => "0000000000011100",
1054 => "0000000000011100",
1055 => "0000000000011100",
1056 => "0000000000011100",
1057 => "0000000000011100",
1058 => "0000000000011100",
1059 => "0000000000011100",
1060 => "0000000000011100",
1061 => "0000000000011100",
1062 => "0000000000011100",
1063 => "0000000000011100",
1064 => "0000000000011100",
1065 => "0000000000011100",
1066 => "0000000000011100",
1067 => "0000000000011100",
1068 => "0000000000011100",
1069 => "0000000000011100",
1070 => "0000000000011100",
1071 => "0000000000011100",
1072 => "0000000000011100",
1073 => "0000000000011100",
1074 => "0000000000011100",
1075 => "0000000000011100",
1076 => "0000000000011100",
1077 => "0000000000011100",
1078 => "0000000000011100",
1079 => "0000000000011100",
1080 => "0000000000011100",
1081 => "0000000000011100",
1082 => "0000000000011100",
1083 => "0000000000011100",
1084 => "0000000000011100",
1085 => "0000000000011100",
1086 => "0000000000011100",
1087 => "0000000000011100",
1088 => "0000000000011100",
1089 => "0000000000011100",
1090 => "0000000000011100",
1091 => "0000000000011100",
1092 => "0000000000011100",
1093 => "0000000000011100",
1094 => "0000000000011100",
1095 => "0000000000011100",
1096 => "0000000000011100",
1097 => "0000000000011100",
1098 => "0000000000011100",
1099 => "0000000000011100",
1100 => "0000000000011100",
1101 => "0000000000011100",
1102 => "0000000000011100",
1103 => "0000000000011100",
1104 => "0000000000011100",
1105 => "0000000000011100",
1106 => "0000000000011100",
1107 => "0000000000011100",
1108 => "0000000000011100",
1109 => "0000000000011100",
1110 => "0000000000011100",
1111 => "0000000000011100",
1112 => "0000000000011100",
1113 => "0000000000011100",
1114 => "0000000000011100",
1115 => "0000000000011100",
1116 => "0000000000011100",
1117 => "0000000000011100",
1118 => "0000000000011100",
1119 => "0000000000011100",
1120 => "0000000000011100",
1121 => "0000000000011100",
1122 => "0000000000011100",
1123 => "0000000000011100",
1124 => "0000000000011100",
1125 => "0000000000011100",
1126 => "0000000000011100",
1127 => "0000000000011100",
1128 => "0000000000011100",
1129 => "0000000000011100",
1130 => "0000000000011100",
1131 => "0000000000011100",
1132 => "0000000000011100",
1133 => "0000000000011100",
1134 => "0000000000011100",
1135 => "0000000000011100",
1136 => "0000000000011100",
1137 => "0000000000011101",
1138 => "0000000000011101",
1139 => "0000000000011101",
1140 => "0000000000011101",
1141 => "0000000000011101",
1142 => "0000000000011101",
1143 => "0000000000011101",
1144 => "0000000000011101",
1145 => "0000000000011101",
1146 => "0000000000011101",
1147 => "0000000000011101",
1148 => "0000000000011101",
1149 => "0000000000011101",
1150 => "0000000000011101",
1151 => "0000000000011101",
1152 => "0000000000011101",
1153 => "0000000000011101",
1154 => "0000000000011101",
1155 => "0000000000011101",
1156 => "0000000000011101",
1157 => "0000000000011101",
1158 => "0000000000011101",
1159 => "0000000000011101",
1160 => "0000000000011101",
1161 => "0000000000011101",
1162 => "0000000000011101",
1163 => "0000000000011101",
1164 => "0000000000011101",
1165 => "0000000000011101",
1166 => "0000000000011101",
1167 => "0000000000011101",
1168 => "0000000000011101",
1169 => "0000000000011101",
1170 => "0000000000011101",
1171 => "0000000000011101",
1172 => "0000000000011101",
1173 => "0000000000011101",
1174 => "0000000000011101",
1175 => "0000000000011101",
1176 => "0000000000011101",
1177 => "0000000000011101",
1178 => "0000000000011101",
1179 => "0000000000011101",
1180 => "0000000000011101",
1181 => "0000000000011101",
1182 => "0000000000011101",
1183 => "0000000000011101",
1184 => "0000000000011101",
1185 => "0000000000011101",
1186 => "0000000000011101",
1187 => "0000000000011101",
1188 => "0000000000011101",
1189 => "0000000000011101",
1190 => "0000000000011101",
1191 => "0000000000011101",
1192 => "0000000000011101",
1193 => "0000000000011101",
1194 => "0000000000011101",
1195 => "0000000000011101",
1196 => "0000000000011101",
1197 => "0000000000011101",
1198 => "0000000000011101",
1199 => "0000000000011101",
1200 => "0000000000011101",
1201 => "0000000000011101",
1202 => "0000000000011101",
1203 => "0000000000011101",
1204 => "0000000000011101",
1205 => "0000000000011101",
1206 => "0000000000011101",
1207 => "0000000000011101",
1208 => "0000000000011101",
1209 => "0000000000011101",
1210 => "0000000000011101",
1211 => "0000000000011101",
1212 => "0000000000011101",
1213 => "0000000000011101",
1214 => "0000000000011101",
1215 => "0000000000011101",
1216 => "0000000000011101",
1217 => "0000000000011101",
1218 => "0000000000011101",
1219 => "0000000000011101",
1220 => "0000000000011101",
1221 => "0000000000011101",
1222 => "0000000000011101",
1223 => "0000000000011101",
1224 => "0000000000011101",
1225 => "0000000000011101",
1226 => "0000000000011101",
1227 => "0000000000011101",
1228 => "0000000000011101",
1229 => "0000000000011101",
1230 => "0000000000011101",
1231 => "0000000000011101",
1232 => "0000000000011101",
1233 => "0000000000011101",
1234 => "0000000000011101",
1235 => "0000000000011101",
1236 => "0000000000011101",
1237 => "0000000000011101",
1238 => "0000000000011101",
1239 => "0000000000011101",
1240 => "0000000000011101",
1241 => "0000000000011101",
1242 => "0000000000011101",
1243 => "0000000000011101",
1244 => "0000000000011101",
1245 => "0000000000011101",
1246 => "0000000000011101",
1247 => "0000000000011101",
1248 => "0000000000011101",
1249 => "0000000000011101",
1250 => "0000000000011101",
1251 => "0000000000011101",
1252 => "0000000000011101",
1253 => "0000000000011101",
1254 => "0000000000011101",
1255 => "0000000000011101",
1256 => "0000000000011101",
1257 => "0000000000011101",
1258 => "0000000000011101",
1259 => "0000000000011101",
1260 => "0000000000011101",
1261 => "0000000000011101",
1262 => "0000000000011101",
1263 => "0000000000011101",
1264 => "0000000000011101",
1265 => "0000000000011101",
1266 => "0000000000011101",
1267 => "0000000000011101",
1268 => "0000000000011101",
1269 => "0000000000011101",
1270 => "0000000000011101",
1271 => "0000000000011101",
1272 => "0000000000011101",
1273 => "0000000000011101",
1274 => "0000000000011101",
1275 => "0000000000011101",
1276 => "0000000000011110",
1277 => "0000000000011110",
1278 => "0000000000011110",
1279 => "0000000000011110",
1280 => "0000000000011110",
1281 => "0000000000011110",
1282 => "0000000000011110",
1283 => "0000000000011110",
1284 => "0000000000011110",
1285 => "0000000000011110",
1286 => "0000000000011110",
1287 => "0000000000011110",
1288 => "0000000000011110",
1289 => "0000000000011110",
1290 => "0000000000011110",
1291 => "0000000000011110",
1292 => "0000000000011110",
1293 => "0000000000011110",
1294 => "0000000000011110",
1295 => "0000000000011110",
1296 => "0000000000011110",
1297 => "0000000000011110",
1298 => "0000000000011110",
1299 => "0000000000011110",
1300 => "0000000000011110",
1301 => "0000000000011110",
1302 => "0000000000011110",
1303 => "0000000000011110",
1304 => "0000000000011110",
1305 => "0000000000011110",
1306 => "0000000000011110",
1307 => "0000000000011110",
1308 => "0000000000011110",
1309 => "0000000000011110",
1310 => "0000000000011110",
1311 => "0000000000011110",
1312 => "0000000000011110",
1313 => "0000000000011110",
1314 => "0000000000011110",
1315 => "0000000000011110",
1316 => "0000000000011110",
1317 => "0000000000011110",
1318 => "0000000000011110",
1319 => "0000000000011110",
1320 => "0000000000011110",
1321 => "0000000000011110",
1322 => "0000000000011110",
1323 => "0000000000011110",
1324 => "0000000000011110",
1325 => "0000000000011110",
1326 => "0000000000011110",
1327 => "0000000000011110",
1328 => "0000000000011110",
1329 => "0000000000011110",
1330 => "0000000000011110",
1331 => "0000000000011110",
1332 => "0000000000011110",
1333 => "0000000000011110",
1334 => "0000000000011110",
1335 => "0000000000011110",
1336 => "0000000000011110",
1337 => "0000000000011110",
1338 => "0000000000011110",
1339 => "0000000000011110",
1340 => "0000000000011110",
1341 => "0000000000011110",
1342 => "0000000000011110",
1343 => "0000000000011110",
1344 => "0000000000011110",
1345 => "0000000000011110",
1346 => "0000000000011110",
1347 => "0000000000011110",
1348 => "0000000000011110",
1349 => "0000000000011110",
1350 => "0000000000011110",
1351 => "0000000000011110",
1352 => "0000000000011110",
1353 => "0000000000011110",
1354 => "0000000000011110",
1355 => "0000000000011110",
1356 => "0000000000011110",
1357 => "0000000000011110",
1358 => "0000000000011110",
1359 => "0000000000011110",
1360 => "0000000000011110",
1361 => "0000000000011110",
1362 => "0000000000011110",
1363 => "0000000000011110",
1364 => "0000000000011110",
1365 => "0000000000011110",
1366 => "0000000000011110",
1367 => "0000000000011110",
1368 => "0000000000011110",
1369 => "0000000000011110",
1370 => "0000000000011110",
1371 => "0000000000011110",
1372 => "0000000000011110",
1373 => "0000000000011110",
1374 => "0000000000011110",
1375 => "0000000000011110",
1376 => "0000000000011110",
1377 => "0000000000011110",
1378 => "0000000000011110",
1379 => "0000000000011110",
1380 => "0000000000011110",
1381 => "0000000000011110",
1382 => "0000000000011110",
1383 => "0000000000011110",
1384 => "0000000000011110",
1385 => "0000000000011110",
1386 => "0000000000011110",
1387 => "0000000000011110",
1388 => "0000000000011110",
1389 => "0000000000011110",
1390 => "0000000000011110",
1391 => "0000000000011110",
1392 => "0000000000011110",
1393 => "0000000000011110",
1394 => "0000000000011110",
1395 => "0000000000011110",
1396 => "0000000000011110",
1397 => "0000000000011110",
1398 => "0000000000011110",
1399 => "0000000000011110",
1400 => "0000000000011110",
1401 => "0000000000011110",
1402 => "0000000000011110",
1403 => "0000000000011110",
1404 => "0000000000011110",
1405 => "0000000000011110",
1406 => "0000000000011110",
1407 => "0000000000011110",
1408 => "0000000000011110",
1409 => "0000000000011110",
1410 => "0000000000011111",
1411 => "0000000000011111",
1412 => "0000000000011111",
1413 => "0000000000011111",
1414 => "0000000000011111",
1415 => "0000000000011111",
1416 => "0000000000011111",
1417 => "0000000000011111",
1418 => "0000000000011111",
1419 => "0000000000011111",
1420 => "0000000000011111",
1421 => "0000000000011111",
1422 => "0000000000011111",
1423 => "0000000000011111",
1424 => "0000000000011111",
1425 => "0000000000011111",
1426 => "0000000000011111",
1427 => "0000000000011111",
1428 => "0000000000011111",
1429 => "0000000000011111",
1430 => "0000000000011111",
1431 => "0000000000011111",
1432 => "0000000000011111",
1433 => "0000000000011111",
1434 => "0000000000011111",
1435 => "0000000000011111",
1436 => "0000000000011111",
1437 => "0000000000011111",
1438 => "0000000000011111",
1439 => "0000000000011111",
1440 => "0000000000011111",
1441 => "0000000000011111",
1442 => "0000000000011111",
1443 => "0000000000011111",
1444 => "0000000000011111",
1445 => "0000000000011111",
1446 => "0000000000011111",
1447 => "0000000000011111",
1448 => "0000000000011111",
1449 => "0000000000011111",
1450 => "0000000000011111",
1451 => "0000000000011111",
1452 => "0000000000011111",
1453 => "0000000000011111",
1454 => "0000000000011111",
1455 => "0000000000011111",
1456 => "0000000000011111",
1457 => "0000000000011111",
1458 => "0000000000011111",
1459 => "0000000000011111",
1460 => "0000000000011111",
1461 => "0000000000011111",
1462 => "0000000000011111",
1463 => "0000000000011111",
1464 => "0000000000011111",
1465 => "0000000000011111",
1466 => "0000000000011111",
1467 => "0000000000011111",
1468 => "0000000000011111",
1469 => "0000000000011111",
1470 => "0000000000011111",
1471 => "0000000000011111",
1472 => "0000000000011111",
1473 => "0000000000011111",
1474 => "0000000000011111",
1475 => "0000000000011111",
1476 => "0000000000011111",
1477 => "0000000000011111",
1478 => "0000000000011111",
1479 => "0000000000011111",
1480 => "0000000000011111",
1481 => "0000000000011111",
1482 => "0000000000011111",
1483 => "0000000000011111",
1484 => "0000000000011111",
1485 => "0000000000011111",
1486 => "0000000000011111",
1487 => "0000000000011111",
1488 => "0000000000011111",
1489 => "0000000000011111",
1490 => "0000000000011111",
1491 => "0000000000011111",
1492 => "0000000000011111",
1493 => "0000000000011111",
1494 => "0000000000011111",
1495 => "0000000000011111",
1496 => "0000000000011111",
1497 => "0000000000011111",
1498 => "0000000000011111",
1499 => "0000000000011111",
1500 => "0000000000011111",
1501 => "0000000000011111",
1502 => "0000000000011111",
1503 => "0000000000011111",
1504 => "0000000000011111",
1505 => "0000000000011111",
1506 => "0000000000011111",
1507 => "0000000000011111",
1508 => "0000000000011111",
1509 => "0000000000011111",
1510 => "0000000000011111",
1511 => "0000000000011111",
1512 => "0000000000011111",
1513 => "0000000000011111",
1514 => "0000000000011111",
1515 => "0000000000011111",
1516 => "0000000000011111",
1517 => "0000000000011111",
1518 => "0000000000011111",
1519 => "0000000000011111",
1520 => "0000000000011111",
1521 => "0000000000011111",
1522 => "0000000000011111",
1523 => "0000000000011111",
1524 => "0000000000011111",
1525 => "0000000000011111",
1526 => "0000000000011111",
1527 => "0000000000011111",
1528 => "0000000000011111",
1529 => "0000000000011111",
1530 => "0000000000011111",
1531 => "0000000000011111",
1532 => "0000000000011111",
1533 => "0000000000011111",
1534 => "0000000000011111",
1535 => "0000000000011111",
1536 => "0000000000011111",
1537 => "0000000000011111",
1538 => "0000000000011111",
1539 => "0000000000011111",
1540 => "0000000000100000",
1541 => "0000000000100000",
1542 => "0000000000100000",
1543 => "0000000000100000",
1544 => "0000000000100000",
1545 => "0000000000100000",
1546 => "0000000000100000",
1547 => "0000000000100000",
1548 => "0000000000100000",
1549 => "0000000000100000",
1550 => "0000000000100000",
1551 => "0000000000100000",
1552 => "0000000000100000",
1553 => "0000000000100000",
1554 => "0000000000100000",
1555 => "0000000000100000",
1556 => "0000000000100000",
1557 => "0000000000100000",
1558 => "0000000000100000",
1559 => "0000000000100000",
1560 => "0000000000100000",
1561 => "0000000000100000",
1562 => "0000000000100000",
1563 => "0000000000100000",
1564 => "0000000000100000",
1565 => "0000000000100000",
1566 => "0000000000100000",
1567 => "0000000000100000",
1568 => "0000000000100000",
1569 => "0000000000100000",
1570 => "0000000000100000",
1571 => "0000000000100000",
1572 => "0000000000100000",
1573 => "0000000000100000",
1574 => "0000000000100000",
1575 => "0000000000100000",
1576 => "0000000000100000",
1577 => "0000000000100000",
1578 => "0000000000100000",
1579 => "0000000000100000",
1580 => "0000000000100000",
1581 => "0000000000100000",
1582 => "0000000000100000",
1583 => "0000000000100000",
1584 => "0000000000100000",
1585 => "0000000000100000",
1586 => "0000000000100000",
1587 => "0000000000100000",
1588 => "0000000000100000",
1589 => "0000000000100000",
1590 => "0000000000100000",
1591 => "0000000000100000",
1592 => "0000000000100000",
1593 => "0000000000100000",
1594 => "0000000000100000",
1595 => "0000000000100000",
1596 => "0000000000100000",
1597 => "0000000000100000",
1598 => "0000000000100000",
1599 => "0000000000100000",
1600 => "0000000000100000",
1601 => "0000000000100000",
1602 => "0000000000100000",
1603 => "0000000000100000",
1604 => "0000000000100000",
1605 => "0000000000100000",
1606 => "0000000000100000",
1607 => "0000000000100000",
1608 => "0000000000100000",
1609 => "0000000000100000",
1610 => "0000000000100000",
1611 => "0000000000100000",
1612 => "0000000000100000",
1613 => "0000000000100000",
1614 => "0000000000100000",
1615 => "0000000000100000",
1616 => "0000000000100000",
1617 => "0000000000100000",
1618 => "0000000000100000",
1619 => "0000000000100000",
1620 => "0000000000100000",
1621 => "0000000000100000",
1622 => "0000000000100000",
1623 => "0000000000100000",
1624 => "0000000000100000",
1625 => "0000000000100000",
1626 => "0000000000100000",
1627 => "0000000000100000",
1628 => "0000000000100000",
1629 => "0000000000100000",
1630 => "0000000000100000",
1631 => "0000000000100000",
1632 => "0000000000100000",
1633 => "0000000000100000",
1634 => "0000000000100000",
1635 => "0000000000100000",
1636 => "0000000000100000",
1637 => "0000000000100000",
1638 => "0000000000100000",
1639 => "0000000000100000",
1640 => "0000000000100000",
1641 => "0000000000100000",
1642 => "0000000000100000",
1643 => "0000000000100000",
1644 => "0000000000100000",
1645 => "0000000000100000",
1646 => "0000000000100000",
1647 => "0000000000100000",
1648 => "0000000000100000",
1649 => "0000000000100000",
1650 => "0000000000100000",
1651 => "0000000000100000",
1652 => "0000000000100000",
1653 => "0000000000100000",
1654 => "0000000000100000",
1655 => "0000000000100000",
1656 => "0000000000100000",
1657 => "0000000000100000",
1658 => "0000000000100000",
1659 => "0000000000100000",
1660 => "0000000000100000",
1661 => "0000000000100000",
1662 => "0000000000100000",
1663 => "0000000000100000",
1664 => "0000000000100000",
1665 => "0000000000100000",
1666 => "0000000000100001",
1667 => "0000000000100001",
1668 => "0000000000100001",
1669 => "0000000000100001",
1670 => "0000000000100001",
1671 => "0000000000100001",
1672 => "0000000000100001",
1673 => "0000000000100001",
1674 => "0000000000100001",
1675 => "0000000000100001",
1676 => "0000000000100001",
1677 => "0000000000100001",
1678 => "0000000000100001",
1679 => "0000000000100001",
1680 => "0000000000100001",
1681 => "0000000000100001",
1682 => "0000000000100001",
1683 => "0000000000100001",
1684 => "0000000000100001",
1685 => "0000000000100001",
1686 => "0000000000100001",
1687 => "0000000000100001",
1688 => "0000000000100001",
1689 => "0000000000100001",
1690 => "0000000000100001",
1691 => "0000000000100001",
1692 => "0000000000100001",
1693 => "0000000000100001",
1694 => "0000000000100001",
1695 => "0000000000100001",
1696 => "0000000000100001",
1697 => "0000000000100001",
1698 => "0000000000100001",
1699 => "0000000000100001",
1700 => "0000000000100001",
1701 => "0000000000100001",
1702 => "0000000000100001",
1703 => "0000000000100001",
1704 => "0000000000100001",
1705 => "0000000000100001",
1706 => "0000000000100001",
1707 => "0000000000100001",
1708 => "0000000000100001",
1709 => "0000000000100001",
1710 => "0000000000100001",
1711 => "0000000000100001",
1712 => "0000000000100001",
1713 => "0000000000100001",
1714 => "0000000000100001",
1715 => "0000000000100001",
1716 => "0000000000100001",
1717 => "0000000000100001",
1718 => "0000000000100001",
1719 => "0000000000100001",
1720 => "0000000000100001",
1721 => "0000000000100001",
1722 => "0000000000100001",
1723 => "0000000000100001",
1724 => "0000000000100001",
1725 => "0000000000100001",
1726 => "0000000000100001",
1727 => "0000000000100001",
1728 => "0000000000100001",
1729 => "0000000000100001",
1730 => "0000000000100001",
1731 => "0000000000100001",
1732 => "0000000000100001",
1733 => "0000000000100001",
1734 => "0000000000100001",
1735 => "0000000000100001",
1736 => "0000000000100001",
1737 => "0000000000100001",
1738 => "0000000000100001",
1739 => "0000000000100001",
1740 => "0000000000100001",
1741 => "0000000000100001",
1742 => "0000000000100001",
1743 => "0000000000100001",
1744 => "0000000000100001",
1745 => "0000000000100001",
1746 => "0000000000100001",
1747 => "0000000000100001",
1748 => "0000000000100001",
1749 => "0000000000100001",
1750 => "0000000000100001",
1751 => "0000000000100001",
1752 => "0000000000100001",
1753 => "0000000000100001",
1754 => "0000000000100001",
1755 => "0000000000100001",
1756 => "0000000000100001",
1757 => "0000000000100001",
1758 => "0000000000100001",
1759 => "0000000000100001",
1760 => "0000000000100001",
1761 => "0000000000100001",
1762 => "0000000000100001",
1763 => "0000000000100001",
1764 => "0000000000100001",
1765 => "0000000000100001",
1766 => "0000000000100001",
1767 => "0000000000100001",
1768 => "0000000000100001",
1769 => "0000000000100001",
1770 => "0000000000100001",
1771 => "0000000000100001",
1772 => "0000000000100001",
1773 => "0000000000100001",
1774 => "0000000000100001",
1775 => "0000000000100001",
1776 => "0000000000100001",
1777 => "0000000000100001",
1778 => "0000000000100001",
1779 => "0000000000100001",
1780 => "0000000000100001",
1781 => "0000000000100001",
1782 => "0000000000100001",
1783 => "0000000000100001",
1784 => "0000000000100001",
1785 => "0000000000100001",
1786 => "0000000000100001",
1787 => "0000000000100001",
1788 => "0000000000100010",
1789 => "0000000000100010",
1790 => "0000000000100010",
1791 => "0000000000100010",
1792 => "0000000000100010",
1793 => "0000000000100010",
1794 => "0000000000100010",
1795 => "0000000000100010",
1796 => "0000000000100010",
1797 => "0000000000100010",
1798 => "0000000000100010",
1799 => "0000000000100010",
1800 => "0000000000100010",
1801 => "0000000000100010",
1802 => "0000000000100010",
1803 => "0000000000100010",
1804 => "0000000000100010",
1805 => "0000000000100010",
1806 => "0000000000100010",
1807 => "0000000000100010",
1808 => "0000000000100010",
1809 => "0000000000100010",
1810 => "0000000000100010",
1811 => "0000000000100010",
1812 => "0000000000100010",
1813 => "0000000000100010",
1814 => "0000000000100010",
1815 => "0000000000100010",
1816 => "0000000000100010",
1817 => "0000000000100010",
1818 => "0000000000100010",
1819 => "0000000000100010",
1820 => "0000000000100010",
1821 => "0000000000100010",
1822 => "0000000000100010",
1823 => "0000000000100010",
1824 => "0000000000100010",
1825 => "0000000000100010",
1826 => "0000000000100010",
1827 => "0000000000100010",
1828 => "0000000000100010",
1829 => "0000000000100010",
1830 => "0000000000100010",
1831 => "0000000000100010",
1832 => "0000000000100010",
1833 => "0000000000100010",
1834 => "0000000000100010",
1835 => "0000000000100010",
1836 => "0000000000100010",
1837 => "0000000000100010",
1838 => "0000000000100010",
1839 => "0000000000100010",
1840 => "0000000000100010",
1841 => "0000000000100010",
1842 => "0000000000100010",
1843 => "0000000000100010",
1844 => "0000000000100010",
1845 => "0000000000100010",
1846 => "0000000000100010",
1847 => "0000000000100010",
1848 => "0000000000100010",
1849 => "0000000000100010",
1850 => "0000000000100010",
1851 => "0000000000100010",
1852 => "0000000000100010",
1853 => "0000000000100010",
1854 => "0000000000100010",
1855 => "0000000000100010",
1856 => "0000000000100010",
1857 => "0000000000100010",
1858 => "0000000000100010",
1859 => "0000000000100010",
1860 => "0000000000100010",
1861 => "0000000000100010",
1862 => "0000000000100010",
1863 => "0000000000100010",
1864 => "0000000000100010",
1865 => "0000000000100010",
1866 => "0000000000100010",
1867 => "0000000000100010",
1868 => "0000000000100010",
1869 => "0000000000100010",
1870 => "0000000000100010",
1871 => "0000000000100010",
1872 => "0000000000100010",
1873 => "0000000000100010",
1874 => "0000000000100010",
1875 => "0000000000100010",
1876 => "0000000000100010",
1877 => "0000000000100010",
1878 => "0000000000100010",
1879 => "0000000000100010",
1880 => "0000000000100010",
1881 => "0000000000100010",
1882 => "0000000000100010",
1883 => "0000000000100010",
1884 => "0000000000100010",
1885 => "0000000000100010",
1886 => "0000000000100010",
1887 => "0000000000100010",
1888 => "0000000000100010",
1889 => "0000000000100010",
1890 => "0000000000100010",
1891 => "0000000000100010",
1892 => "0000000000100010",
1893 => "0000000000100010",
1894 => "0000000000100010",
1895 => "0000000000100010",
1896 => "0000000000100010",
1897 => "0000000000100010",
1898 => "0000000000100010",
1899 => "0000000000100010",
1900 => "0000000000100010",
1901 => "0000000000100010",
1902 => "0000000000100010",
1903 => "0000000000100010",
1904 => "0000000000100010",
1905 => "0000000000100010",
1906 => "0000000000100010",
1907 => "0000000000100011",
1908 => "0000000000100011",
1909 => "0000000000100011",
1910 => "0000000000100011",
1911 => "0000000000100011",
1912 => "0000000000100011",
1913 => "0000000000100011",
1914 => "0000000000100011",
1915 => "0000000000100011",
1916 => "0000000000100011",
1917 => "0000000000100011",
1918 => "0000000000100011",
1919 => "0000000000100011",
1920 => "0000000000100011",
1921 => "0000000000100011",
1922 => "0000000000100011",
1923 => "0000000000100011",
1924 => "0000000000100011",
1925 => "0000000000100011",
1926 => "0000000000100011",
1927 => "0000000000100011",
1928 => "0000000000100011",
1929 => "0000000000100011",
1930 => "0000000000100011",
1931 => "0000000000100011",
1932 => "0000000000100011",
1933 => "0000000000100011",
1934 => "0000000000100011",
1935 => "0000000000100011",
1936 => "0000000000100011",
1937 => "0000000000100011",
1938 => "0000000000100011",
1939 => "0000000000100011",
1940 => "0000000000100011",
1941 => "0000000000100011",
1942 => "0000000000100011",
1943 => "0000000000100011",
1944 => "0000000000100011",
1945 => "0000000000100011",
1946 => "0000000000100011",
1947 => "0000000000100011",
1948 => "0000000000100011",
1949 => "0000000000100011",
1950 => "0000000000100011",
1951 => "0000000000100011",
1952 => "0000000000100011",
1953 => "0000000000100011",
1954 => "0000000000100011",
1955 => "0000000000100011",
1956 => "0000000000100011",
1957 => "0000000000100011",
1958 => "0000000000100011",
1959 => "0000000000100011",
1960 => "0000000000100011",
1961 => "0000000000100011",
1962 => "0000000000100011",
1963 => "0000000000100011",
1964 => "0000000000100011",
1965 => "0000000000100011",
1966 => "0000000000100011",
1967 => "0000000000100011",
1968 => "0000000000100011",
1969 => "0000000000100011",
1970 => "0000000000100011",
1971 => "0000000000100011",
1972 => "0000000000100011",
1973 => "0000000000100011",
1974 => "0000000000100011",
1975 => "0000000000100011",
1976 => "0000000000100011",
1977 => "0000000000100011",
1978 => "0000000000100011",
1979 => "0000000000100011",
1980 => "0000000000100011",
1981 => "0000000000100011",
1982 => "0000000000100011",
1983 => "0000000000100011",
1984 => "0000000000100011",
1985 => "0000000000100011",
1986 => "0000000000100011",
1987 => "0000000000100011",
1988 => "0000000000100011",
1989 => "0000000000100011",
1990 => "0000000000100011",
1991 => "0000000000100011",
1992 => "0000000000100011",
1993 => "0000000000100011",
1994 => "0000000000100011",
1995 => "0000000000100011",
1996 => "0000000000100011",
1997 => "0000000000100011",
1998 => "0000000000100011",
1999 => "0000000000100011",
2000 => "0000000000100011",
2001 => "0000000000100011",
2002 => "0000000000100011",
2003 => "0000000000100011",
2004 => "0000000000100011",
2005 => "0000000000100011",
2006 => "0000000000100011",
2007 => "0000000000100011",
2008 => "0000000000100011",
2009 => "0000000000100011",
2010 => "0000000000100011",
2011 => "0000000000100011",
2012 => "0000000000100011",
2013 => "0000000000100011",
2014 => "0000000000100011",
2015 => "0000000000100011",
2016 => "0000000000100011",
2017 => "0000000000100011",
2018 => "0000000000100011",
2019 => "0000000000100011",
2020 => "0000000000100011",
2021 => "0000000000100011",
2022 => "0000000000100011",
2023 => "0000000000100100",
2024 => "0000000000100100",
2025 => "0000000000100100",
2026 => "0000000000100100",
2027 => "0000000000100100",
2028 => "0000000000100100",
2029 => "0000000000100100",
2030 => "0000000000100100",
2031 => "0000000000100100",
2032 => "0000000000100100",
2033 => "0000000000100100",
2034 => "0000000000100100",
2035 => "0000000000100100",
2036 => "0000000000100100",
2037 => "0000000000100100",
2038 => "0000000000100100",
2039 => "0000000000100100",
2040 => "0000000000100100",
2041 => "0000000000100100",
2042 => "0000000000100100",
2043 => "0000000000100100",
2044 => "0000000000100100",
2045 => "0000000000100100",
2046 => "0000000000100100",
2047 => "0000000000100100",
2048 => "0000000000100100",
2049 => "0000000000100100",
2050 => "0000000000100100",
2051 => "0000000000100100",
2052 => "0000000000100100",
2053 => "0000000000100100",
2054 => "0000000000100100",
2055 => "0000000000100100",
2056 => "0000000000100100",
2057 => "0000000000100100",
2058 => "0000000000100100",
2059 => "0000000000100100",
2060 => "0000000000100100",
2061 => "0000000000100100",
2062 => "0000000000100100",
2063 => "0000000000100100",
2064 => "0000000000100100",
2065 => "0000000000100100",
2066 => "0000000000100100",
2067 => "0000000000100100",
2068 => "0000000000100100",
2069 => "0000000000100100",
2070 => "0000000000100100",
2071 => "0000000000100100",
2072 => "0000000000100100",
2073 => "0000000000100100",
2074 => "0000000000100100",
2075 => "0000000000100100",
2076 => "0000000000100100",
2077 => "0000000000100100",
2078 => "0000000000100100",
2079 => "0000000000100100",
2080 => "0000000000100100",
2081 => "0000000000100100",
2082 => "0000000000100100",
2083 => "0000000000100100",
2084 => "0000000000100100",
2085 => "0000000000100100",
2086 => "0000000000100100",
2087 => "0000000000100100",
2088 => "0000000000100100",
2089 => "0000000000100100",
2090 => "0000000000100100",
2091 => "0000000000100100",
2092 => "0000000000100100",
2093 => "0000000000100100",
2094 => "0000000000100100",
2095 => "0000000000100100",
2096 => "0000000000100100",
2097 => "0000000000100100",
2098 => "0000000000100100",
2099 => "0000000000100100",
2100 => "0000000000100100",
2101 => "0000000000100100",
2102 => "0000000000100100",
2103 => "0000000000100100",
2104 => "0000000000100100",
2105 => "0000000000100100",
2106 => "0000000000100100",
2107 => "0000000000100100",
2108 => "0000000000100100",
2109 => "0000000000100100",
2110 => "0000000000100100",
2111 => "0000000000100100",
2112 => "0000000000100100",
2113 => "0000000000100100",
2114 => "0000000000100100",
2115 => "0000000000100100",
2116 => "0000000000100100",
2117 => "0000000000100100",
2118 => "0000000000100100",
2119 => "0000000000100100",
2120 => "0000000000100100",
2121 => "0000000000100100",
2122 => "0000000000100100",
2123 => "0000000000100100",
2124 => "0000000000100100",
2125 => "0000000000100100",
2126 => "0000000000100100",
2127 => "0000000000100100",
2128 => "0000000000100100",
2129 => "0000000000100100",
2130 => "0000000000100100",
2131 => "0000000000100100",
2132 => "0000000000100100",
2133 => "0000000000100100",
2134 => "0000000000100100",
2135 => "0000000000100101",
2136 => "0000000000100101",
2137 => "0000000000100101",
2138 => "0000000000100101",
2139 => "0000000000100101",
2140 => "0000000000100101",
2141 => "0000000000100101",
2142 => "0000000000100101",
2143 => "0000000000100101",
2144 => "0000000000100101",
2145 => "0000000000100101",
2146 => "0000000000100101",
2147 => "0000000000100101",
2148 => "0000000000100101",
2149 => "0000000000100101",
2150 => "0000000000100101",
2151 => "0000000000100101",
2152 => "0000000000100101",
2153 => "0000000000100101",
2154 => "0000000000100101",
2155 => "0000000000100101",
2156 => "0000000000100101",
2157 => "0000000000100101",
2158 => "0000000000100101",
2159 => "0000000000100101",
2160 => "0000000000100101",
2161 => "0000000000100101",
2162 => "0000000000100101",
2163 => "0000000000100101",
2164 => "0000000000100101",
2165 => "0000000000100101",
2166 => "0000000000100101",
2167 => "0000000000100101",
2168 => "0000000000100101",
2169 => "0000000000100101",
2170 => "0000000000100101",
2171 => "0000000000100101",
2172 => "0000000000100101",
2173 => "0000000000100101",
2174 => "0000000000100101",
2175 => "0000000000100101",
2176 => "0000000000100101",
2177 => "0000000000100101",
2178 => "0000000000100101",
2179 => "0000000000100101",
2180 => "0000000000100101",
2181 => "0000000000100101",
2182 => "0000000000100101",
2183 => "0000000000100101",
2184 => "0000000000100101",
2185 => "0000000000100101",
2186 => "0000000000100101",
2187 => "0000000000100101",
2188 => "0000000000100101",
2189 => "0000000000100101",
2190 => "0000000000100101",
2191 => "0000000000100101",
2192 => "0000000000100101",
2193 => "0000000000100101",
2194 => "0000000000100101",
2195 => "0000000000100101",
2196 => "0000000000100101",
2197 => "0000000000100101",
2198 => "0000000000100101",
2199 => "0000000000100101",
2200 => "0000000000100101",
2201 => "0000000000100101",
2202 => "0000000000100101",
2203 => "0000000000100101",
2204 => "0000000000100101",
2205 => "0000000000100101",
2206 => "0000000000100101",
2207 => "0000000000100101",
2208 => "0000000000100101",
2209 => "0000000000100101",
2210 => "0000000000100101",
2211 => "0000000000100101",
2212 => "0000000000100101",
2213 => "0000000000100101",
2214 => "0000000000100101",
2215 => "0000000000100101",
2216 => "0000000000100101",
2217 => "0000000000100101",
2218 => "0000000000100101",
2219 => "0000000000100101",
2220 => "0000000000100101",
2221 => "0000000000100101",
2222 => "0000000000100101",
2223 => "0000000000100101",
2224 => "0000000000100101",
2225 => "0000000000100101",
2226 => "0000000000100101",
2227 => "0000000000100101",
2228 => "0000000000100101",
2229 => "0000000000100101",
2230 => "0000000000100101",
2231 => "0000000000100101",
2232 => "0000000000100101",
2233 => "0000000000100101",
2234 => "0000000000100101",
2235 => "0000000000100101",
2236 => "0000000000100101",
2237 => "0000000000100101",
2238 => "0000000000100101",
2239 => "0000000000100101",
2240 => "0000000000100101",
2241 => "0000000000100101",
2242 => "0000000000100101",
2243 => "0000000000100101",
2244 => "0000000000100110",
2245 => "0000000000100110",
2246 => "0000000000100110",
2247 => "0000000000100110",
2248 => "0000000000100110",
2249 => "0000000000100110",
2250 => "0000000000100110",
2251 => "0000000000100110",
2252 => "0000000000100110",
2253 => "0000000000100110",
2254 => "0000000000100110",
2255 => "0000000000100110",
2256 => "0000000000100110",
2257 => "0000000000100110",
2258 => "0000000000100110",
2259 => "0000000000100110",
2260 => "0000000000100110",
2261 => "0000000000100110",
2262 => "0000000000100110",
2263 => "0000000000100110",
2264 => "0000000000100110",
2265 => "0000000000100110",
2266 => "0000000000100110",
2267 => "0000000000100110",
2268 => "0000000000100110",
2269 => "0000000000100110",
2270 => "0000000000100110",
2271 => "0000000000100110",
2272 => "0000000000100110",
2273 => "0000000000100110",
2274 => "0000000000100110",
2275 => "0000000000100110",
2276 => "0000000000100110",
2277 => "0000000000100110",
2278 => "0000000000100110",
2279 => "0000000000100110",
2280 => "0000000000100110",
2281 => "0000000000100110",
2282 => "0000000000100110",
2283 => "0000000000100110",
2284 => "0000000000100110",
2285 => "0000000000100110",
2286 => "0000000000100110",
2287 => "0000000000100110",
2288 => "0000000000100110",
2289 => "0000000000100110",
2290 => "0000000000100110",
2291 => "0000000000100110",
2292 => "0000000000100110",
2293 => "0000000000100110",
2294 => "0000000000100110",
2295 => "0000000000100110",
2296 => "0000000000100110",
2297 => "0000000000100110",
2298 => "0000000000100110",
2299 => "0000000000100110",
2300 => "0000000000100110",
2301 => "0000000000100110",
2302 => "0000000000100110",
2303 => "0000000000100110",
2304 => "0000000000100110",
2305 => "0000000000100110",
2306 => "0000000000100110",
2307 => "0000000000100110",
2308 => "0000000000100110",
2309 => "0000000000100110",
2310 => "0000000000100110",
2311 => "0000000000100110",
2312 => "0000000000100110",
2313 => "0000000000100110",
2314 => "0000000000100110",
2315 => "0000000000100110",
2316 => "0000000000100110",
2317 => "0000000000100110",
2318 => "0000000000100110",
2319 => "0000000000100110",
2320 => "0000000000100110",
2321 => "0000000000100110",
2322 => "0000000000100110",
2323 => "0000000000100110",
2324 => "0000000000100110",
2325 => "0000000000100110",
2326 => "0000000000100110",
2327 => "0000000000100110",
2328 => "0000000000100110",
2329 => "0000000000100110",
2330 => "0000000000100110",
2331 => "0000000000100110",
2332 => "0000000000100110",
2333 => "0000000000100110",
2334 => "0000000000100110",
2335 => "0000000000100110",
2336 => "0000000000100110",
2337 => "0000000000100110",
2338 => "0000000000100110",
2339 => "0000000000100110",
2340 => "0000000000100110",
2341 => "0000000000100110",
2342 => "0000000000100110",
2343 => "0000000000100110",
2344 => "0000000000100110",
2345 => "0000000000100110",
2346 => "0000000000100110",
2347 => "0000000000100110",
2348 => "0000000000100110",
2349 => "0000000000100110",
2350 => "0000000000100110",
2351 => "0000000000100111",
2352 => "0000000000100111",
2353 => "0000000000100111",
2354 => "0000000000100111",
2355 => "0000000000100111",
2356 => "0000000000100111",
2357 => "0000000000100111",
2358 => "0000000000100111",
2359 => "0000000000100111",
2360 => "0000000000100111",
2361 => "0000000000100111",
2362 => "0000000000100111",
2363 => "0000000000100111",
2364 => "0000000000100111",
2365 => "0000000000100111",
2366 => "0000000000100111",
2367 => "0000000000100111",
2368 => "0000000000100111",
2369 => "0000000000100111",
2370 => "0000000000100111",
2371 => "0000000000100111",
2372 => "0000000000100111",
2373 => "0000000000100111",
2374 => "0000000000100111",
2375 => "0000000000100111",
2376 => "0000000000100111",
2377 => "0000000000100111",
2378 => "0000000000100111",
2379 => "0000000000100111",
2380 => "0000000000100111",
2381 => "0000000000100111",
2382 => "0000000000100111",
2383 => "0000000000100111",
2384 => "0000000000100111",
2385 => "0000000000100111",
2386 => "0000000000100111",
2387 => "0000000000100111",
2388 => "0000000000100111",
2389 => "0000000000100111",
2390 => "0000000000100111",
2391 => "0000000000100111",
2392 => "0000000000100111",
2393 => "0000000000100111",
2394 => "0000000000100111",
2395 => "0000000000100111",
2396 => "0000000000100111",
2397 => "0000000000100111",
2398 => "0000000000100111",
2399 => "0000000000100111",
2400 => "0000000000100111",
2401 => "0000000000100111",
2402 => "0000000000100111",
2403 => "0000000000100111",
2404 => "0000000000100111",
2405 => "0000000000100111",
2406 => "0000000000100111",
2407 => "0000000000100111",
2408 => "0000000000100111",
2409 => "0000000000100111",
2410 => "0000000000100111",
2411 => "0000000000100111",
2412 => "0000000000100111",
2413 => "0000000000100111",
2414 => "0000000000100111",
2415 => "0000000000100111",
2416 => "0000000000100111",
2417 => "0000000000100111",
2418 => "0000000000100111",
2419 => "0000000000100111",
2420 => "0000000000100111",
2421 => "0000000000100111",
2422 => "0000000000100111",
2423 => "0000000000100111",
2424 => "0000000000100111",
2425 => "0000000000100111",
2426 => "0000000000100111",
2427 => "0000000000100111",
2428 => "0000000000100111",
2429 => "0000000000100111",
2430 => "0000000000100111",
2431 => "0000000000100111",
2432 => "0000000000100111",
2433 => "0000000000100111",
2434 => "0000000000100111",
2435 => "0000000000100111",
2436 => "0000000000100111",
2437 => "0000000000100111",
2438 => "0000000000100111",
2439 => "0000000000100111",
2440 => "0000000000100111",
2441 => "0000000000100111",
2442 => "0000000000100111",
2443 => "0000000000100111",
2444 => "0000000000100111",
2445 => "0000000000100111",
2446 => "0000000000100111",
2447 => "0000000000100111",
2448 => "0000000000100111",
2449 => "0000000000100111",
2450 => "0000000000100111",
2451 => "0000000000100111",
2452 => "0000000000100111",
2453 => "0000000000100111",
2454 => "0000000000100111",
2455 => "0000000000101000",
2456 => "0000000000101000",
2457 => "0000000000101000",
2458 => "0000000000101000",
2459 => "0000000000101000",
2460 => "0000000000101000",
2461 => "0000000000101000",
2462 => "0000000000101000",
2463 => "0000000000101000",
2464 => "0000000000101000",
2465 => "0000000000101000",
2466 => "0000000000101000",
2467 => "0000000000101000",
2468 => "0000000000101000",
2469 => "0000000000101000",
2470 => "0000000000101000",
2471 => "0000000000101000",
2472 => "0000000000101000",
2473 => "0000000000101000",
2474 => "0000000000101000",
2475 => "0000000000101000",
2476 => "0000000000101000",
2477 => "0000000000101000",
2478 => "0000000000101000",
2479 => "0000000000101000",
2480 => "0000000000101000",
2481 => "0000000000101000",
2482 => "0000000000101000",
2483 => "0000000000101000",
2484 => "0000000000101000",
2485 => "0000000000101000",
2486 => "0000000000101000",
2487 => "0000000000101000",
2488 => "0000000000101000",
2489 => "0000000000101000",
2490 => "0000000000101000",
2491 => "0000000000101000",
2492 => "0000000000101000",
2493 => "0000000000101000",
2494 => "0000000000101000",
2495 => "0000000000101000",
2496 => "0000000000101000",
2497 => "0000000000101000",
2498 => "0000000000101000",
2499 => "0000000000101000",
2500 => "0000000000101000",
2501 => "0000000000101000",
2502 => "0000000000101000",
2503 => "0000000000101000",
2504 => "0000000000101000",
2505 => "0000000000101000",
2506 => "0000000000101000",
2507 => "0000000000101000",
2508 => "0000000000101000",
2509 => "0000000000101000",
2510 => "0000000000101000",
2511 => "0000000000101000",
2512 => "0000000000101000",
2513 => "0000000000101000",
2514 => "0000000000101000",
2515 => "0000000000101000",
2516 => "0000000000101000",
2517 => "0000000000101000",
2518 => "0000000000101000",
2519 => "0000000000101000",
2520 => "0000000000101000",
2521 => "0000000000101000",
2522 => "0000000000101000",
2523 => "0000000000101000",
2524 => "0000000000101000",
2525 => "0000000000101000",
2526 => "0000000000101000",
2527 => "0000000000101000",
2528 => "0000000000101000",
2529 => "0000000000101000",
2530 => "0000000000101000",
2531 => "0000000000101000",
2532 => "0000000000101000",
2533 => "0000000000101000",
2534 => "0000000000101000",
2535 => "0000000000101000",
2536 => "0000000000101000",
2537 => "0000000000101000",
2538 => "0000000000101000",
2539 => "0000000000101000",
2540 => "0000000000101000",
2541 => "0000000000101000",
2542 => "0000000000101000",
2543 => "0000000000101000",
2544 => "0000000000101000",
2545 => "0000000000101000",
2546 => "0000000000101000",
2547 => "0000000000101000",
2548 => "0000000000101000",
2549 => "0000000000101000",
2550 => "0000000000101000",
2551 => "0000000000101000",
2552 => "0000000000101000",
2553 => "0000000000101000",
2554 => "0000000000101000",
2555 => "0000000000101000",
2556 => "0000000000101001",
2557 => "0000000000101001",
2558 => "0000000000101001",
2559 => "0000000000101001",
2560 => "0000000000101001",
2561 => "0000000000101001",
2562 => "0000000000101001",
2563 => "0000000000101001",
2564 => "0000000000101001",
2565 => "0000000000101001",
2566 => "0000000000101001",
2567 => "0000000000101001",
2568 => "0000000000101001",
2569 => "0000000000101001",
2570 => "0000000000101001",
2571 => "0000000000101001",
2572 => "0000000000101001",
2573 => "0000000000101001",
2574 => "0000000000101001",
2575 => "0000000000101001",
2576 => "0000000000101001",
2577 => "0000000000101001",
2578 => "0000000000101001",
2579 => "0000000000101001",
2580 => "0000000000101001",
2581 => "0000000000101001",
2582 => "0000000000101001",
2583 => "0000000000101001",
2584 => "0000000000101001",
2585 => "0000000000101001",
2586 => "0000000000101001",
2587 => "0000000000101001",
2588 => "0000000000101001",
2589 => "0000000000101001",
2590 => "0000000000101001",
2591 => "0000000000101001",
2592 => "0000000000101001",
2593 => "0000000000101001",
2594 => "0000000000101001",
2595 => "0000000000101001",
2596 => "0000000000101001",
2597 => "0000000000101001",
2598 => "0000000000101001",
2599 => "0000000000101001",
2600 => "0000000000101001",
2601 => "0000000000101001",
2602 => "0000000000101001",
2603 => "0000000000101001",
2604 => "0000000000101001",
2605 => "0000000000101001",
2606 => "0000000000101001",
2607 => "0000000000101001",
2608 => "0000000000101001",
2609 => "0000000000101001",
2610 => "0000000000101001",
2611 => "0000000000101001",
2612 => "0000000000101001",
2613 => "0000000000101001",
2614 => "0000000000101001",
2615 => "0000000000101001",
2616 => "0000000000101001",
2617 => "0000000000101001",
2618 => "0000000000101001",
2619 => "0000000000101001",
2620 => "0000000000101001",
2621 => "0000000000101001",
2622 => "0000000000101001",
2623 => "0000000000101001",
2624 => "0000000000101001",
2625 => "0000000000101001",
2626 => "0000000000101001",
2627 => "0000000000101001",
2628 => "0000000000101001",
2629 => "0000000000101001",
2630 => "0000000000101001",
2631 => "0000000000101001",
2632 => "0000000000101001",
2633 => "0000000000101001",
2634 => "0000000000101001",
2635 => "0000000000101001",
2636 => "0000000000101001",
2637 => "0000000000101001",
2638 => "0000000000101001",
2639 => "0000000000101001",
2640 => "0000000000101001",
2641 => "0000000000101001",
2642 => "0000000000101001",
2643 => "0000000000101001",
2644 => "0000000000101001",
2645 => "0000000000101001",
2646 => "0000000000101001",
2647 => "0000000000101001",
2648 => "0000000000101001",
2649 => "0000000000101001",
2650 => "0000000000101001",
2651 => "0000000000101001",
2652 => "0000000000101001",
2653 => "0000000000101001",
2654 => "0000000000101010",
2655 => "0000000000101010",
2656 => "0000000000101010",
2657 => "0000000000101010",
2658 => "0000000000101010",
2659 => "0000000000101010",
2660 => "0000000000101010",
2661 => "0000000000101010",
2662 => "0000000000101010",
2663 => "0000000000101010",
2664 => "0000000000101010",
2665 => "0000000000101010",
2666 => "0000000000101010",
2667 => "0000000000101010",
2668 => "0000000000101010",
2669 => "0000000000101010",
2670 => "0000000000101010",
2671 => "0000000000101010",
2672 => "0000000000101010",
2673 => "0000000000101010",
2674 => "0000000000101010",
2675 => "0000000000101010",
2676 => "0000000000101010",
2677 => "0000000000101010",
2678 => "0000000000101010",
2679 => "0000000000101010",
2680 => "0000000000101010",
2681 => "0000000000101010",
2682 => "0000000000101010",
2683 => "0000000000101010",
2684 => "0000000000101010",
2685 => "0000000000101010",
2686 => "0000000000101010",
2687 => "0000000000101010",
2688 => "0000000000101010",
2689 => "0000000000101010",
2690 => "0000000000101010",
2691 => "0000000000101010",
2692 => "0000000000101010",
2693 => "0000000000101010",
2694 => "0000000000101010",
2695 => "0000000000101010",
2696 => "0000000000101010",
2697 => "0000000000101010",
2698 => "0000000000101010",
2699 => "0000000000101010",
2700 => "0000000000101010",
2701 => "0000000000101010",
2702 => "0000000000101010",
2703 => "0000000000101010",
2704 => "0000000000101010",
2705 => "0000000000101010",
2706 => "0000000000101010",
2707 => "0000000000101010",
2708 => "0000000000101010",
2709 => "0000000000101010",
2710 => "0000000000101010",
2711 => "0000000000101010",
2712 => "0000000000101010",
2713 => "0000000000101010",
2714 => "0000000000101010",
2715 => "0000000000101010",
2716 => "0000000000101010",
2717 => "0000000000101010",
2718 => "0000000000101010",
2719 => "0000000000101010",
2720 => "0000000000101010",
2721 => "0000000000101010",
2722 => "0000000000101010",
2723 => "0000000000101010",
2724 => "0000000000101010",
2725 => "0000000000101010",
2726 => "0000000000101010",
2727 => "0000000000101010",
2728 => "0000000000101010",
2729 => "0000000000101010",
2730 => "0000000000101010",
2731 => "0000000000101010",
2732 => "0000000000101010",
2733 => "0000000000101010",
2734 => "0000000000101010",
2735 => "0000000000101010",
2736 => "0000000000101010",
2737 => "0000000000101010",
2738 => "0000000000101010",
2739 => "0000000000101010",
2740 => "0000000000101010",
2741 => "0000000000101010",
2742 => "0000000000101010",
2743 => "0000000000101010",
2744 => "0000000000101010",
2745 => "0000000000101010",
2746 => "0000000000101010",
2747 => "0000000000101010",
2748 => "0000000000101010",
2749 => "0000000000101010",
2750 => "0000000000101010",
2751 => "0000000000101011",
2752 => "0000000000101011",
2753 => "0000000000101011",
2754 => "0000000000101011",
2755 => "0000000000101011",
2756 => "0000000000101011",
2757 => "0000000000101011",
2758 => "0000000000101011",
2759 => "0000000000101011",
2760 => "0000000000101011",
2761 => "0000000000101011",
2762 => "0000000000101011",
2763 => "0000000000101011",
2764 => "0000000000101011",
2765 => "0000000000101011",
2766 => "0000000000101011",
2767 => "0000000000101011",
2768 => "0000000000101011",
2769 => "0000000000101011",
2770 => "0000000000101011",
2771 => "0000000000101011",
2772 => "0000000000101011",
2773 => "0000000000101011",
2774 => "0000000000101011",
2775 => "0000000000101011",
2776 => "0000000000101011",
2777 => "0000000000101011",
2778 => "0000000000101011",
2779 => "0000000000101011",
2780 => "0000000000101011",
2781 => "0000000000101011",
2782 => "0000000000101011",
2783 => "0000000000101011",
2784 => "0000000000101011",
2785 => "0000000000101011",
2786 => "0000000000101011",
2787 => "0000000000101011",
2788 => "0000000000101011",
2789 => "0000000000101011",
2790 => "0000000000101011",
2791 => "0000000000101011",
2792 => "0000000000101011",
2793 => "0000000000101011",
2794 => "0000000000101011",
2795 => "0000000000101011",
2796 => "0000000000101011",
2797 => "0000000000101011",
2798 => "0000000000101011",
2799 => "0000000000101011",
2800 => "0000000000101011",
2801 => "0000000000101011",
2802 => "0000000000101011",
2803 => "0000000000101011",
2804 => "0000000000101011",
2805 => "0000000000101011",
2806 => "0000000000101011",
2807 => "0000000000101011",
2808 => "0000000000101011",
2809 => "0000000000101011",
2810 => "0000000000101011",
2811 => "0000000000101011",
2812 => "0000000000101011",
2813 => "0000000000101011",
2814 => "0000000000101011",
2815 => "0000000000101011",
2816 => "0000000000101011",
2817 => "0000000000101011",
2818 => "0000000000101011",
2819 => "0000000000101011",
2820 => "0000000000101011",
2821 => "0000000000101011",
2822 => "0000000000101011",
2823 => "0000000000101011",
2824 => "0000000000101011",
2825 => "0000000000101011",
2826 => "0000000000101011",
2827 => "0000000000101011",
2828 => "0000000000101011",
2829 => "0000000000101011",
2830 => "0000000000101011",
2831 => "0000000000101011",
2832 => "0000000000101011",
2833 => "0000000000101011",
2834 => "0000000000101011",
2835 => "0000000000101011",
2836 => "0000000000101011",
2837 => "0000000000101011",
2838 => "0000000000101011",
2839 => "0000000000101011",
2840 => "0000000000101011",
2841 => "0000000000101011",
2842 => "0000000000101011",
2843 => "0000000000101011",
2844 => "0000000000101011",
2845 => "0000000000101100",
2846 => "0000000000101100",
2847 => "0000000000101100",
2848 => "0000000000101100",
2849 => "0000000000101100",
2850 => "0000000000101100",
2851 => "0000000000101100",
2852 => "0000000000101100",
2853 => "0000000000101100",
2854 => "0000000000101100",
2855 => "0000000000101100",
2856 => "0000000000101100",
2857 => "0000000000101100",
2858 => "0000000000101100",
2859 => "0000000000101100",
2860 => "0000000000101100",
2861 => "0000000000101100",
2862 => "0000000000101100",
2863 => "0000000000101100",
2864 => "0000000000101100",
2865 => "0000000000101100",
2866 => "0000000000101100",
2867 => "0000000000101100",
2868 => "0000000000101100",
2869 => "0000000000101100",
2870 => "0000000000101100",
2871 => "0000000000101100",
2872 => "0000000000101100",
2873 => "0000000000101100",
2874 => "0000000000101100",
2875 => "0000000000101100",
2876 => "0000000000101100",
2877 => "0000000000101100",
2878 => "0000000000101100",
2879 => "0000000000101100",
2880 => "0000000000101100",
2881 => "0000000000101100",
2882 => "0000000000101100",
2883 => "0000000000101100",
2884 => "0000000000101100",
2885 => "0000000000101100",
2886 => "0000000000101100",
2887 => "0000000000101100",
2888 => "0000000000101100",
2889 => "0000000000101100",
2890 => "0000000000101100",
2891 => "0000000000101100",
2892 => "0000000000101100",
2893 => "0000000000101100",
2894 => "0000000000101100",
2895 => "0000000000101100",
2896 => "0000000000101100",
2897 => "0000000000101100",
2898 => "0000000000101100",
2899 => "0000000000101100",
2900 => "0000000000101100",
2901 => "0000000000101100",
2902 => "0000000000101100",
2903 => "0000000000101100",
2904 => "0000000000101100",
2905 => "0000000000101100",
2906 => "0000000000101100",
2907 => "0000000000101100",
2908 => "0000000000101100",
2909 => "0000000000101100",
2910 => "0000000000101100",
2911 => "0000000000101100",
2912 => "0000000000101100",
2913 => "0000000000101100",
2914 => "0000000000101100",
2915 => "0000000000101100",
2916 => "0000000000101100",
2917 => "0000000000101100",
2918 => "0000000000101100",
2919 => "0000000000101100",
2920 => "0000000000101100",
2921 => "0000000000101100",
2922 => "0000000000101100",
2923 => "0000000000101100",
2924 => "0000000000101100",
2925 => "0000000000101100",
2926 => "0000000000101100",
2927 => "0000000000101100",
2928 => "0000000000101100",
2929 => "0000000000101100",
2930 => "0000000000101100",
2931 => "0000000000101100",
2932 => "0000000000101100",
2933 => "0000000000101100",
2934 => "0000000000101100",
2935 => "0000000000101100",
2936 => "0000000000101100",
2937 => "0000000000101101",
2938 => "0000000000101101",
2939 => "0000000000101101",
2940 => "0000000000101101",
2941 => "0000000000101101",
2942 => "0000000000101101",
2943 => "0000000000101101",
2944 => "0000000000101101",
2945 => "0000000000101101",
2946 => "0000000000101101",
2947 => "0000000000101101",
2948 => "0000000000101101",
2949 => "0000000000101101",
2950 => "0000000000101101",
2951 => "0000000000101101",
2952 => "0000000000101101",
2953 => "0000000000101101",
2954 => "0000000000101101",
2955 => "0000000000101101",
2956 => "0000000000101101",
2957 => "0000000000101101",
2958 => "0000000000101101",
2959 => "0000000000101101",
2960 => "0000000000101101",
2961 => "0000000000101101",
2962 => "0000000000101101",
2963 => "0000000000101101",
2964 => "0000000000101101",
2965 => "0000000000101101",
2966 => "0000000000101101",
2967 => "0000000000101101",
2968 => "0000000000101101",
2969 => "0000000000101101",
2970 => "0000000000101101",
2971 => "0000000000101101",
2972 => "0000000000101101",
2973 => "0000000000101101",
2974 => "0000000000101101",
2975 => "0000000000101101",
2976 => "0000000000101101",
2977 => "0000000000101101",
2978 => "0000000000101101",
2979 => "0000000000101101",
2980 => "0000000000101101",
2981 => "0000000000101101",
2982 => "0000000000101101",
2983 => "0000000000101101",
2984 => "0000000000101101",
2985 => "0000000000101101",
2986 => "0000000000101101",
2987 => "0000000000101101",
2988 => "0000000000101101",
2989 => "0000000000101101",
2990 => "0000000000101101",
2991 => "0000000000101101",
2992 => "0000000000101101",
2993 => "0000000000101101",
2994 => "0000000000101101",
2995 => "0000000000101101",
2996 => "0000000000101101",
2997 => "0000000000101101",
2998 => "0000000000101101",
2999 => "0000000000101101",
3000 => "0000000000101101",
3001 => "0000000000101101",
3002 => "0000000000101101",
3003 => "0000000000101101",
3004 => "0000000000101101",
3005 => "0000000000101101",
3006 => "0000000000101101",
3007 => "0000000000101101",
3008 => "0000000000101101",
3009 => "0000000000101101",
3010 => "0000000000101101",
3011 => "0000000000101101",
3012 => "0000000000101101",
3013 => "0000000000101101",
3014 => "0000000000101101",
3015 => "0000000000101101",
3016 => "0000000000101101",
3017 => "0000000000101101",
3018 => "0000000000101101",
3019 => "0000000000101101",
3020 => "0000000000101101",
3021 => "0000000000101101",
3022 => "0000000000101101",
3023 => "0000000000101101",
3024 => "0000000000101101",
3025 => "0000000000101101",
3026 => "0000000000101101",
3027 => "0000000000101110",
3028 => "0000000000101110",
3029 => "0000000000101110",
3030 => "0000000000101110",
3031 => "0000000000101110",
3032 => "0000000000101110",
3033 => "0000000000101110",
3034 => "0000000000101110",
3035 => "0000000000101110",
3036 => "0000000000101110",
3037 => "0000000000101110",
3038 => "0000000000101110",
3039 => "0000000000101110",
3040 => "0000000000101110",
3041 => "0000000000101110",
3042 => "0000000000101110",
3043 => "0000000000101110",
3044 => "0000000000101110",
3045 => "0000000000101110",
3046 => "0000000000101110",
3047 => "0000000000101110",
3048 => "0000000000101110",
3049 => "0000000000101110",
3050 => "0000000000101110",
3051 => "0000000000101110",
3052 => "0000000000101110",
3053 => "0000000000101110",
3054 => "0000000000101110",
3055 => "0000000000101110",
3056 => "0000000000101110",
3057 => "0000000000101110",
3058 => "0000000000101110",
3059 => "0000000000101110",
3060 => "0000000000101110",
3061 => "0000000000101110",
3062 => "0000000000101110",
3063 => "0000000000101110",
3064 => "0000000000101110",
3065 => "0000000000101110",
3066 => "0000000000101110",
3067 => "0000000000101110",
3068 => "0000000000101110",
3069 => "0000000000101110",
3070 => "0000000000101110",
3071 => "0000000000101110",
3072 => "0000000000101110",
3073 => "0000000000101110",
3074 => "0000000000101110",
3075 => "0000000000101110",
3076 => "0000000000101110",
3077 => "0000000000101110",
3078 => "0000000000101110",
3079 => "0000000000101110",
3080 => "0000000000101110",
3081 => "0000000000101110",
3082 => "0000000000101110",
3083 => "0000000000101110",
3084 => "0000000000101110",
3085 => "0000000000101110",
3086 => "0000000000101110",
3087 => "0000000000101110",
3088 => "0000000000101110",
3089 => "0000000000101110",
3090 => "0000000000101110",
3091 => "0000000000101110",
3092 => "0000000000101110",
3093 => "0000000000101110",
3094 => "0000000000101110",
3095 => "0000000000101110",
3096 => "0000000000101110",
3097 => "0000000000101110",
3098 => "0000000000101110",
3099 => "0000000000101110",
3100 => "0000000000101110",
3101 => "0000000000101110",
3102 => "0000000000101110",
3103 => "0000000000101110",
3104 => "0000000000101110",
3105 => "0000000000101110",
3106 => "0000000000101110",
3107 => "0000000000101110",
3108 => "0000000000101110",
3109 => "0000000000101110",
3110 => "0000000000101110",
3111 => "0000000000101110",
3112 => "0000000000101110",
3113 => "0000000000101110",
3114 => "0000000000101110",
3115 => "0000000000101110",
3116 => "0000000000101111",
3117 => "0000000000101111",
3118 => "0000000000101111",
3119 => "0000000000101111",
3120 => "0000000000101111",
3121 => "0000000000101111",
3122 => "0000000000101111",
3123 => "0000000000101111",
3124 => "0000000000101111",
3125 => "0000000000101111",
3126 => "0000000000101111",
3127 => "0000000000101111",
3128 => "0000000000101111",
3129 => "0000000000101111",
3130 => "0000000000101111",
3131 => "0000000000101111",
3132 => "0000000000101111",
3133 => "0000000000101111",
3134 => "0000000000101111",
3135 => "0000000000101111",
3136 => "0000000000101111",
3137 => "0000000000101111",
3138 => "0000000000101111",
3139 => "0000000000101111",
3140 => "0000000000101111",
3141 => "0000000000101111",
3142 => "0000000000101111",
3143 => "0000000000101111",
3144 => "0000000000101111",
3145 => "0000000000101111",
3146 => "0000000000101111",
3147 => "0000000000101111",
3148 => "0000000000101111",
3149 => "0000000000101111",
3150 => "0000000000101111",
3151 => "0000000000101111",
3152 => "0000000000101111",
3153 => "0000000000101111",
3154 => "0000000000101111",
3155 => "0000000000101111",
3156 => "0000000000101111",
3157 => "0000000000101111",
3158 => "0000000000101111",
3159 => "0000000000101111",
3160 => "0000000000101111",
3161 => "0000000000101111",
3162 => "0000000000101111",
3163 => "0000000000101111",
3164 => "0000000000101111",
3165 => "0000000000101111",
3166 => "0000000000101111",
3167 => "0000000000101111",
3168 => "0000000000101111",
3169 => "0000000000101111",
3170 => "0000000000101111",
3171 => "0000000000101111",
3172 => "0000000000101111",
3173 => "0000000000101111",
3174 => "0000000000101111",
3175 => "0000000000101111",
3176 => "0000000000101111",
3177 => "0000000000101111",
3178 => "0000000000101111",
3179 => "0000000000101111",
3180 => "0000000000101111",
3181 => "0000000000101111",
3182 => "0000000000101111",
3183 => "0000000000101111",
3184 => "0000000000101111",
3185 => "0000000000101111",
3186 => "0000000000101111",
3187 => "0000000000101111",
3188 => "0000000000101111",
3189 => "0000000000101111",
3190 => "0000000000101111",
3191 => "0000000000101111",
3192 => "0000000000101111",
3193 => "0000000000101111",
3194 => "0000000000101111",
3195 => "0000000000101111",
3196 => "0000000000101111",
3197 => "0000000000101111",
3198 => "0000000000101111",
3199 => "0000000000101111",
3200 => "0000000000101111",
3201 => "0000000000101111",
3202 => "0000000000110000",
3203 => "0000000000110000",
3204 => "0000000000110000",
3205 => "0000000000110000",
3206 => "0000000000110000",
3207 => "0000000000110000",
3208 => "0000000000110000",
3209 => "0000000000110000",
3210 => "0000000000110000",
3211 => "0000000000110000",
3212 => "0000000000110000",
3213 => "0000000000110000",
3214 => "0000000000110000",
3215 => "0000000000110000",
3216 => "0000000000110000",
3217 => "0000000000110000",
3218 => "0000000000110000",
3219 => "0000000000110000",
3220 => "0000000000110000",
3221 => "0000000000110000",
3222 => "0000000000110000",
3223 => "0000000000110000",
3224 => "0000000000110000",
3225 => "0000000000110000",
3226 => "0000000000110000",
3227 => "0000000000110000",
3228 => "0000000000110000",
3229 => "0000000000110000",
3230 => "0000000000110000",
3231 => "0000000000110000",
3232 => "0000000000110000",
3233 => "0000000000110000",
3234 => "0000000000110000",
3235 => "0000000000110000",
3236 => "0000000000110000",
3237 => "0000000000110000",
3238 => "0000000000110000",
3239 => "0000000000110000",
3240 => "0000000000110000",
3241 => "0000000000110000",
3242 => "0000000000110000",
3243 => "0000000000110000",
3244 => "0000000000110000",
3245 => "0000000000110000",
3246 => "0000000000110000",
3247 => "0000000000110000",
3248 => "0000000000110000",
3249 => "0000000000110000",
3250 => "0000000000110000",
3251 => "0000000000110000",
3252 => "0000000000110000",
3253 => "0000000000110000",
3254 => "0000000000110000",
3255 => "0000000000110000",
3256 => "0000000000110000",
3257 => "0000000000110000",
3258 => "0000000000110000",
3259 => "0000000000110000",
3260 => "0000000000110000",
3261 => "0000000000110000",
3262 => "0000000000110000",
3263 => "0000000000110000",
3264 => "0000000000110000",
3265 => "0000000000110000",
3266 => "0000000000110000",
3267 => "0000000000110000",
3268 => "0000000000110000",
3269 => "0000000000110000",
3270 => "0000000000110000",
3271 => "0000000000110000",
3272 => "0000000000110000",
3273 => "0000000000110000",
3274 => "0000000000110000",
3275 => "0000000000110000",
3276 => "0000000000110000",
3277 => "0000000000110000",
3278 => "0000000000110000",
3279 => "0000000000110000",
3280 => "0000000000110000",
3281 => "0000000000110000",
3282 => "0000000000110000",
3283 => "0000000000110000",
3284 => "0000000000110000",
3285 => "0000000000110000",
3286 => "0000000000110001",
3287 => "0000000000110001",
3288 => "0000000000110001",
3289 => "0000000000110001",
3290 => "0000000000110001",
3291 => "0000000000110001",
3292 => "0000000000110001",
3293 => "0000000000110001",
3294 => "0000000000110001",
3295 => "0000000000110001",
3296 => "0000000000110001",
3297 => "0000000000110001",
3298 => "0000000000110001",
3299 => "0000000000110001",
3300 => "0000000000110001",
3301 => "0000000000110001",
3302 => "0000000000110001",
3303 => "0000000000110001",
3304 => "0000000000110001",
3305 => "0000000000110001",
3306 => "0000000000110001",
3307 => "0000000000110001",
3308 => "0000000000110001",
3309 => "0000000000110001",
3310 => "0000000000110001",
3311 => "0000000000110001",
3312 => "0000000000110001",
3313 => "0000000000110001",
3314 => "0000000000110001",
3315 => "0000000000110001",
3316 => "0000000000110001",
3317 => "0000000000110001",
3318 => "0000000000110001",
3319 => "0000000000110001",
3320 => "0000000000110001",
3321 => "0000000000110001",
3322 => "0000000000110001",
3323 => "0000000000110001",
3324 => "0000000000110001",
3325 => "0000000000110001",
3326 => "0000000000110001",
3327 => "0000000000110001",
3328 => "0000000000110001",
3329 => "0000000000110001",
3330 => "0000000000110001",
3331 => "0000000000110001",
3332 => "0000000000110001",
3333 => "0000000000110001",
3334 => "0000000000110001",
3335 => "0000000000110001",
3336 => "0000000000110001",
3337 => "0000000000110001",
3338 => "0000000000110001",
3339 => "0000000000110001",
3340 => "0000000000110001",
3341 => "0000000000110001",
3342 => "0000000000110001",
3343 => "0000000000110001",
3344 => "0000000000110001",
3345 => "0000000000110001",
3346 => "0000000000110001",
3347 => "0000000000110001",
3348 => "0000000000110001",
3349 => "0000000000110001",
3350 => "0000000000110001",
3351 => "0000000000110001",
3352 => "0000000000110001",
3353 => "0000000000110001",
3354 => "0000000000110001",
3355 => "0000000000110001",
3356 => "0000000000110001",
3357 => "0000000000110001",
3358 => "0000000000110001",
3359 => "0000000000110001",
3360 => "0000000000110001",
3361 => "0000000000110001",
3362 => "0000000000110001",
3363 => "0000000000110001",
3364 => "0000000000110001",
3365 => "0000000000110001",
3366 => "0000000000110001",
3367 => "0000000000110001",
3368 => "0000000000110001",
3369 => "0000000000110010",
3370 => "0000000000110010",
3371 => "0000000000110010",
3372 => "0000000000110010",
3373 => "0000000000110010",
3374 => "0000000000110010",
3375 => "0000000000110010",
3376 => "0000000000110010",
3377 => "0000000000110010",
3378 => "0000000000110010",
3379 => "0000000000110010",
3380 => "0000000000110010",
3381 => "0000000000110010",
3382 => "0000000000110010",
3383 => "0000000000110010",
3384 => "0000000000110010",
3385 => "0000000000110010",
3386 => "0000000000110010",
3387 => "0000000000110010",
3388 => "0000000000110010",
3389 => "0000000000110010",
3390 => "0000000000110010",
3391 => "0000000000110010",
3392 => "0000000000110010",
3393 => "0000000000110010",
3394 => "0000000000110010",
3395 => "0000000000110010",
3396 => "0000000000110010",
3397 => "0000000000110010",
3398 => "0000000000110010",
3399 => "0000000000110010",
3400 => "0000000000110010",
3401 => "0000000000110010",
3402 => "0000000000110010",
3403 => "0000000000110010",
3404 => "0000000000110010",
3405 => "0000000000110010",
3406 => "0000000000110010",
3407 => "0000000000110010",
3408 => "0000000000110010",
3409 => "0000000000110010",
3410 => "0000000000110010",
3411 => "0000000000110010",
3412 => "0000000000110010",
3413 => "0000000000110010",
3414 => "0000000000110010",
3415 => "0000000000110010",
3416 => "0000000000110010",
3417 => "0000000000110010",
3418 => "0000000000110010",
3419 => "0000000000110010",
3420 => "0000000000110010",
3421 => "0000000000110010",
3422 => "0000000000110010",
3423 => "0000000000110010",
3424 => "0000000000110010",
3425 => "0000000000110010",
3426 => "0000000000110010",
3427 => "0000000000110010",
3428 => "0000000000110010",
3429 => "0000000000110010",
3430 => "0000000000110010",
3431 => "0000000000110010",
3432 => "0000000000110010",
3433 => "0000000000110010",
3434 => "0000000000110010",
3435 => "0000000000110010",
3436 => "0000000000110010",
3437 => "0000000000110010",
3438 => "0000000000110010",
3439 => "0000000000110010",
3440 => "0000000000110010",
3441 => "0000000000110010",
3442 => "0000000000110010",
3443 => "0000000000110010",
3444 => "0000000000110010",
3445 => "0000000000110010",
3446 => "0000000000110010",
3447 => "0000000000110010",
3448 => "0000000000110010",
3449 => "0000000000110010",
3450 => "0000000000110011",
3451 => "0000000000110011",
3452 => "0000000000110011",
3453 => "0000000000110011",
3454 => "0000000000110011",
3455 => "0000000000110011",
3456 => "0000000000110011",
3457 => "0000000000110011",
3458 => "0000000000110011",
3459 => "0000000000110011",
3460 => "0000000000110011",
3461 => "0000000000110011",
3462 => "0000000000110011",
3463 => "0000000000110011",
3464 => "0000000000110011",
3465 => "0000000000110011",
3466 => "0000000000110011",
3467 => "0000000000110011",
3468 => "0000000000110011",
3469 => "0000000000110011",
3470 => "0000000000110011",
3471 => "0000000000110011",
3472 => "0000000000110011",
3473 => "0000000000110011",
3474 => "0000000000110011",
3475 => "0000000000110011",
3476 => "0000000000110011",
3477 => "0000000000110011",
3478 => "0000000000110011",
3479 => "0000000000110011",
3480 => "0000000000110011",
3481 => "0000000000110011",
3482 => "0000000000110011",
3483 => "0000000000110011",
3484 => "0000000000110011",
3485 => "0000000000110011",
3486 => "0000000000110011",
3487 => "0000000000110011",
3488 => "0000000000110011",
3489 => "0000000000110011",
3490 => "0000000000110011",
3491 => "0000000000110011",
3492 => "0000000000110011",
3493 => "0000000000110011",
3494 => "0000000000110011",
3495 => "0000000000110011",
3496 => "0000000000110011",
3497 => "0000000000110011",
3498 => "0000000000110011",
3499 => "0000000000110011",
3500 => "0000000000110011",
3501 => "0000000000110011",
3502 => "0000000000110011",
3503 => "0000000000110011",
3504 => "0000000000110011",
3505 => "0000000000110011",
3506 => "0000000000110011",
3507 => "0000000000110011",
3508 => "0000000000110011",
3509 => "0000000000110011",
3510 => "0000000000110011",
3511 => "0000000000110011",
3512 => "0000000000110011",
3513 => "0000000000110011",
3514 => "0000000000110011",
3515 => "0000000000110011",
3516 => "0000000000110011",
3517 => "0000000000110011",
3518 => "0000000000110011",
3519 => "0000000000110011",
3520 => "0000000000110011",
3521 => "0000000000110011",
3522 => "0000000000110011",
3523 => "0000000000110011",
3524 => "0000000000110011",
3525 => "0000000000110011",
3526 => "0000000000110011",
3527 => "0000000000110011",
3528 => "0000000000110011",
3529 => "0000000000110011",
3530 => "0000000000110100",
3531 => "0000000000110100",
3532 => "0000000000110100",
3533 => "0000000000110100",
3534 => "0000000000110100",
3535 => "0000000000110100",
3536 => "0000000000110100",
3537 => "0000000000110100",
3538 => "0000000000110100",
3539 => "0000000000110100",
3540 => "0000000000110100",
3541 => "0000000000110100",
3542 => "0000000000110100",
3543 => "0000000000110100",
3544 => "0000000000110100",
3545 => "0000000000110100",
3546 => "0000000000110100",
3547 => "0000000000110100",
3548 => "0000000000110100",
3549 => "0000000000110100",
3550 => "0000000000110100",
3551 => "0000000000110100",
3552 => "0000000000110100",
3553 => "0000000000110100",
3554 => "0000000000110100",
3555 => "0000000000110100",
3556 => "0000000000110100",
3557 => "0000000000110100",
3558 => "0000000000110100",
3559 => "0000000000110100",
3560 => "0000000000110100",
3561 => "0000000000110100",
3562 => "0000000000110100",
3563 => "0000000000110100",
3564 => "0000000000110100",
3565 => "0000000000110100",
3566 => "0000000000110100",
3567 => "0000000000110100",
3568 => "0000000000110100",
3569 => "0000000000110100",
3570 => "0000000000110100",
3571 => "0000000000110100",
3572 => "0000000000110100",
3573 => "0000000000110100",
3574 => "0000000000110100",
3575 => "0000000000110100",
3576 => "0000000000110100",
3577 => "0000000000110100",
3578 => "0000000000110100",
3579 => "0000000000110100",
3580 => "0000000000110100",
3581 => "0000000000110100",
3582 => "0000000000110100",
3583 => "0000000000110100",
3584 => "0000000000110100",
3585 => "0000000000110100",
3586 => "0000000000110100",
3587 => "0000000000110100",
3588 => "0000000000110100",
3589 => "0000000000110100",
3590 => "0000000000110100",
3591 => "0000000000110100",
3592 => "0000000000110100",
3593 => "0000000000110100",
3594 => "0000000000110100",
3595 => "0000000000110100",
3596 => "0000000000110100",
3597 => "0000000000110100",
3598 => "0000000000110100",
3599 => "0000000000110100",
3600 => "0000000000110100",
3601 => "0000000000110100",
3602 => "0000000000110100",
3603 => "0000000000110100",
3604 => "0000000000110100",
3605 => "0000000000110100",
3606 => "0000000000110100",
3607 => "0000000000110100",
3608 => "0000000000110101",
3609 => "0000000000110101",
3610 => "0000000000110101",
3611 => "0000000000110101",
3612 => "0000000000110101",
3613 => "0000000000110101",
3614 => "0000000000110101",
3615 => "0000000000110101",
3616 => "0000000000110101",
3617 => "0000000000110101",
3618 => "0000000000110101",
3619 => "0000000000110101",
3620 => "0000000000110101",
3621 => "0000000000110101",
3622 => "0000000000110101",
3623 => "0000000000110101",
3624 => "0000000000110101",
3625 => "0000000000110101",
3626 => "0000000000110101",
3627 => "0000000000110101",
3628 => "0000000000110101",
3629 => "0000000000110101",
3630 => "0000000000110101",
3631 => "0000000000110101",
3632 => "0000000000110101",
3633 => "0000000000110101",
3634 => "0000000000110101",
3635 => "0000000000110101",
3636 => "0000000000110101",
3637 => "0000000000110101",
3638 => "0000000000110101",
3639 => "0000000000110101",
3640 => "0000000000110101",
3641 => "0000000000110101",
3642 => "0000000000110101",
3643 => "0000000000110101",
3644 => "0000000000110101",
3645 => "0000000000110101",
3646 => "0000000000110101",
3647 => "0000000000110101",
3648 => "0000000000110101",
3649 => "0000000000110101",
3650 => "0000000000110101",
3651 => "0000000000110101",
3652 => "0000000000110101",
3653 => "0000000000110101",
3654 => "0000000000110101",
3655 => "0000000000110101",
3656 => "0000000000110101",
3657 => "0000000000110101",
3658 => "0000000000110101",
3659 => "0000000000110101",
3660 => "0000000000110101",
3661 => "0000000000110101",
3662 => "0000000000110101",
3663 => "0000000000110101",
3664 => "0000000000110101",
3665 => "0000000000110101",
3666 => "0000000000110101",
3667 => "0000000000110101",
3668 => "0000000000110101",
3669 => "0000000000110101",
3670 => "0000000000110101",
3671 => "0000000000110101",
3672 => "0000000000110101",
3673 => "0000000000110101",
3674 => "0000000000110101",
3675 => "0000000000110101",
3676 => "0000000000110101",
3677 => "0000000000110101",
3678 => "0000000000110101",
3679 => "0000000000110101",
3680 => "0000000000110101",
3681 => "0000000000110101",
3682 => "0000000000110101",
3683 => "0000000000110101",
3684 => "0000000000110101",
3685 => "0000000000110110",
3686 => "0000000000110110",
3687 => "0000000000110110",
3688 => "0000000000110110",
3689 => "0000000000110110",
3690 => "0000000000110110",
3691 => "0000000000110110",
3692 => "0000000000110110",
3693 => "0000000000110110",
3694 => "0000000000110110",
3695 => "0000000000110110",
3696 => "0000000000110110",
3697 => "0000000000110110",
3698 => "0000000000110110",
3699 => "0000000000110110",
3700 => "0000000000110110",
3701 => "0000000000110110",
3702 => "0000000000110110",
3703 => "0000000000110110",
3704 => "0000000000110110",
3705 => "0000000000110110",
3706 => "0000000000110110",
3707 => "0000000000110110",
3708 => "0000000000110110",
3709 => "0000000000110110",
3710 => "0000000000110110",
3711 => "0000000000110110",
3712 => "0000000000110110",
3713 => "0000000000110110",
3714 => "0000000000110110",
3715 => "0000000000110110",
3716 => "0000000000110110",
3717 => "0000000000110110",
3718 => "0000000000110110",
3719 => "0000000000110110",
3720 => "0000000000110110",
3721 => "0000000000110110",
3722 => "0000000000110110",
3723 => "0000000000110110",
3724 => "0000000000110110",
3725 => "0000000000110110",
3726 => "0000000000110110",
3727 => "0000000000110110",
3728 => "0000000000110110",
3729 => "0000000000110110",
3730 => "0000000000110110",
3731 => "0000000000110110",
3732 => "0000000000110110",
3733 => "0000000000110110",
3734 => "0000000000110110",
3735 => "0000000000110110",
3736 => "0000000000110110",
3737 => "0000000000110110",
3738 => "0000000000110110",
3739 => "0000000000110110",
3740 => "0000000000110110",
3741 => "0000000000110110",
3742 => "0000000000110110",
3743 => "0000000000110110",
3744 => "0000000000110110",
3745 => "0000000000110110",
3746 => "0000000000110110",
3747 => "0000000000110110",
3748 => "0000000000110110",
3749 => "0000000000110110",
3750 => "0000000000110110",
3751 => "0000000000110110",
3752 => "0000000000110110",
3753 => "0000000000110110",
3754 => "0000000000110110",
3755 => "0000000000110110",
3756 => "0000000000110110",
3757 => "0000000000110110",
3758 => "0000000000110110",
3759 => "0000000000110110",
3760 => "0000000000110111",
3761 => "0000000000110111",
3762 => "0000000000110111",
3763 => "0000000000110111",
3764 => "0000000000110111",
3765 => "0000000000110111",
3766 => "0000000000110111",
3767 => "0000000000110111",
3768 => "0000000000110111",
3769 => "0000000000110111",
3770 => "0000000000110111",
3771 => "0000000000110111",
3772 => "0000000000110111",
3773 => "0000000000110111",
3774 => "0000000000110111",
3775 => "0000000000110111",
3776 => "0000000000110111",
3777 => "0000000000110111",
3778 => "0000000000110111",
3779 => "0000000000110111",
3780 => "0000000000110111",
3781 => "0000000000110111",
3782 => "0000000000110111",
3783 => "0000000000110111",
3784 => "0000000000110111",
3785 => "0000000000110111",
3786 => "0000000000110111",
3787 => "0000000000110111",
3788 => "0000000000110111",
3789 => "0000000000110111",
3790 => "0000000000110111",
3791 => "0000000000110111",
3792 => "0000000000110111",
3793 => "0000000000110111",
3794 => "0000000000110111",
3795 => "0000000000110111",
3796 => "0000000000110111",
3797 => "0000000000110111",
3798 => "0000000000110111",
3799 => "0000000000110111",
3800 => "0000000000110111",
3801 => "0000000000110111",
3802 => "0000000000110111",
3803 => "0000000000110111",
3804 => "0000000000110111",
3805 => "0000000000110111",
3806 => "0000000000110111",
3807 => "0000000000110111",
3808 => "0000000000110111",
3809 => "0000000000110111",
3810 => "0000000000110111",
3811 => "0000000000110111",
3812 => "0000000000110111",
3813 => "0000000000110111",
3814 => "0000000000110111",
3815 => "0000000000110111",
3816 => "0000000000110111",
3817 => "0000000000110111",
3818 => "0000000000110111",
3819 => "0000000000110111",
3820 => "0000000000110111",
3821 => "0000000000110111",
3822 => "0000000000110111",
3823 => "0000000000110111",
3824 => "0000000000110111",
3825 => "0000000000110111",
3826 => "0000000000110111",
3827 => "0000000000110111",
3828 => "0000000000110111",
3829 => "0000000000110111",
3830 => "0000000000110111",
3831 => "0000000000110111",
3832 => "0000000000110111",
3833 => "0000000000110111",
3834 => "0000000000111000",
3835 => "0000000000111000",
3836 => "0000000000111000",
3837 => "0000000000111000",
3838 => "0000000000111000",
3839 => "0000000000111000",
3840 => "0000000000111000",
3841 => "0000000000111000",
3842 => "0000000000111000",
3843 => "0000000000111000",
3844 => "0000000000111000",
3845 => "0000000000111000",
3846 => "0000000000111000",
3847 => "0000000000111000",
3848 => "0000000000111000",
3849 => "0000000000111000",
3850 => "0000000000111000",
3851 => "0000000000111000",
3852 => "0000000000111000",
3853 => "0000000000111000",
3854 => "0000000000111000",
3855 => "0000000000111000",
3856 => "0000000000111000",
3857 => "0000000000111000",
3858 => "0000000000111000",
3859 => "0000000000111000",
3860 => "0000000000111000",
3861 => "0000000000111000",
3862 => "0000000000111000",
3863 => "0000000000111000",
3864 => "0000000000111000",
3865 => "0000000000111000",
3866 => "0000000000111000",
3867 => "0000000000111000",
3868 => "0000000000111000",
3869 => "0000000000111000",
3870 => "0000000000111000",
3871 => "0000000000111000",
3872 => "0000000000111000",
3873 => "0000000000111000",
3874 => "0000000000111000",
3875 => "0000000000111000",
3876 => "0000000000111000",
3877 => "0000000000111000",
3878 => "0000000000111000",
3879 => "0000000000111000",
3880 => "0000000000111000",
3881 => "0000000000111000",
3882 => "0000000000111000",
3883 => "0000000000111000",
3884 => "0000000000111000",
3885 => "0000000000111000",
3886 => "0000000000111000",
3887 => "0000000000111000",
3888 => "0000000000111000",
3889 => "0000000000111000",
3890 => "0000000000111000",
3891 => "0000000000111000",
3892 => "0000000000111000",
3893 => "0000000000111000",
3894 => "0000000000111000",
3895 => "0000000000111000",
3896 => "0000000000111000",
3897 => "0000000000111000",
3898 => "0000000000111000",
3899 => "0000000000111000",
3900 => "0000000000111000",
3901 => "0000000000111000",
3902 => "0000000000111000",
3903 => "0000000000111000",
3904 => "0000000000111000",
3905 => "0000000000111000",
3906 => "0000000000111001",
3907 => "0000000000111001",
3908 => "0000000000111001",
3909 => "0000000000111001",
3910 => "0000000000111001",
3911 => "0000000000111001",
3912 => "0000000000111001",
3913 => "0000000000111001",
3914 => "0000000000111001",
3915 => "0000000000111001",
3916 => "0000000000111001",
3917 => "0000000000111001",
3918 => "0000000000111001",
3919 => "0000000000111001",
3920 => "0000000000111001",
3921 => "0000000000111001",
3922 => "0000000000111001",
3923 => "0000000000111001",
3924 => "0000000000111001",
3925 => "0000000000111001",
3926 => "0000000000111001",
3927 => "0000000000111001",
3928 => "0000000000111001",
3929 => "0000000000111001",
3930 => "0000000000111001",
3931 => "0000000000111001",
3932 => "0000000000111001",
3933 => "0000000000111001",
3934 => "0000000000111001",
3935 => "0000000000111001",
3936 => "0000000000111001",
3937 => "0000000000111001",
3938 => "0000000000111001",
3939 => "0000000000111001",
3940 => "0000000000111001",
3941 => "0000000000111001",
3942 => "0000000000111001",
3943 => "0000000000111001",
3944 => "0000000000111001",
3945 => "0000000000111001",
3946 => "0000000000111001",
3947 => "0000000000111001",
3948 => "0000000000111001",
3949 => "0000000000111001",
3950 => "0000000000111001",
3951 => "0000000000111001",
3952 => "0000000000111001",
3953 => "0000000000111001",
3954 => "0000000000111001",
3955 => "0000000000111001",
3956 => "0000000000111001",
3957 => "0000000000111001",
3958 => "0000000000111001",
3959 => "0000000000111001",
3960 => "0000000000111001",
3961 => "0000000000111001",
3962 => "0000000000111001",
3963 => "0000000000111001",
3964 => "0000000000111001",
3965 => "0000000000111001",
3966 => "0000000000111001",
3967 => "0000000000111001",
3968 => "0000000000111001",
3969 => "0000000000111001",
3970 => "0000000000111001",
3971 => "0000000000111001",
3972 => "0000000000111001",
3973 => "0000000000111001",
3974 => "0000000000111001",
3975 => "0000000000111001",
3976 => "0000000000111001",
3977 => "0000000000111001",
3978 => "0000000000111010",
3979 => "0000000000111010",
3980 => "0000000000111010",
3981 => "0000000000111010",
3982 => "0000000000111010",
3983 => "0000000000111010",
3984 => "0000000000111010",
3985 => "0000000000111010",
3986 => "0000000000111010",
3987 => "0000000000111010",
3988 => "0000000000111010",
3989 => "0000000000111010",
3990 => "0000000000111010",
3991 => "0000000000111010",
3992 => "0000000000111010",
3993 => "0000000000111010",
3994 => "0000000000111010",
3995 => "0000000000111010",
3996 => "0000000000111010",
3997 => "0000000000111010",
3998 => "0000000000111010",
3999 => "0000000000111010",
4000 => "0000000000111010",
4001 => "0000000000111010",
4002 => "0000000000111010",
4003 => "0000000000111010",
4004 => "0000000000111010",
4005 => "0000000000111010",
4006 => "0000000000111010",
4007 => "0000000000111010",
4008 => "0000000000111010",
4009 => "0000000000111010",
4010 => "0000000000111010",
4011 => "0000000000111010",
4012 => "0000000000111010",
4013 => "0000000000111010",
4014 => "0000000000111010",
4015 => "0000000000111010",
4016 => "0000000000111010",
4017 => "0000000000111010",
4018 => "0000000000111010",
4019 => "0000000000111010",
4020 => "0000000000111010",
4021 => "0000000000111010",
4022 => "0000000000111010",
4023 => "0000000000111010",
4024 => "0000000000111010",
4025 => "0000000000111010",
4026 => "0000000000111010",
4027 => "0000000000111010",
4028 => "0000000000111010",
4029 => "0000000000111010",
4030 => "0000000000111010",
4031 => "0000000000111010",
4032 => "0000000000111010",
4033 => "0000000000111010",
4034 => "0000000000111010",
4035 => "0000000000111010",
4036 => "0000000000111010",
4037 => "0000000000111010",
4038 => "0000000000111010",
4039 => "0000000000111010",
4040 => "0000000000111010",
4041 => "0000000000111010",
4042 => "0000000000111010",
4043 => "0000000000111010",
4044 => "0000000000111010",
4045 => "0000000000111010",
4046 => "0000000000111010",
4047 => "0000000000111010",
4048 => "0000000000111011",
4049 => "0000000000111011",
4050 => "0000000000111011",
4051 => "0000000000111011",
4052 => "0000000000111011",
4053 => "0000000000111011",
4054 => "0000000000111011",
4055 => "0000000000111011",
4056 => "0000000000111011",
4057 => "0000000000111011",
4058 => "0000000000111011",
4059 => "0000000000111011",
4060 => "0000000000111011",
4061 => "0000000000111011",
4062 => "0000000000111011",
4063 => "0000000000111011",
4064 => "0000000000111011",
4065 => "0000000000111011",
4066 => "0000000000111011",
4067 => "0000000000111011",
4068 => "0000000000111011",
4069 => "0000000000111011",
4070 => "0000000000111011",
4071 => "0000000000111011",
4072 => "0000000000111011",
4073 => "0000000000111011",
4074 => "0000000000111011",
4075 => "0000000000111011",
4076 => "0000000000111011",
4077 => "0000000000111011",
4078 => "0000000000111011",
4079 => "0000000000111011",
4080 => "0000000000111011",
4081 => "0000000000111011",
4082 => "0000000000111011",
4083 => "0000000000111011",
4084 => "0000000000111011",
4085 => "0000000000111011",
4086 => "0000000000111011",
4087 => "0000000000111011",
4088 => "0000000000111011",
4089 => "0000000000111011",
4090 => "0000000000111011",
4091 => "0000000000111011",
4092 => "0000000000111011",
4093 => "0000000000111011",
4094 => "0000000000111011",
4095 => "0000000000111011",
4096 => "0000000000111011",
4097 => "0000000000111011",
4098 => "0000000000111011",
4099 => "0000000000111011",
4100 => "0000000000111011",
4101 => "0000000000111011",
4102 => "0000000000111011",
4103 => "0000000000111011",
4104 => "0000000000111011",
4105 => "0000000000111011",
4106 => "0000000000111011",
4107 => "0000000000111011",
4108 => "0000000000111011",
4109 => "0000000000111011",
4110 => "0000000000111011",
4111 => "0000000000111011",
4112 => "0000000000111011",
4113 => "0000000000111011",
4114 => "0000000000111011",
4115 => "0000000000111011",
4116 => "0000000000111011",
4117 => "0000000000111100",
4118 => "0000000000111100",
4119 => "0000000000111100",
4120 => "0000000000111100",
4121 => "0000000000111100",
4122 => "0000000000111100",
4123 => "0000000000111100",
4124 => "0000000000111100",
4125 => "0000000000111100",
4126 => "0000000000111100",
4127 => "0000000000111100",
4128 => "0000000000111100",
4129 => "0000000000111100",
4130 => "0000000000111100",
4131 => "0000000000111100",
4132 => "0000000000111100",
4133 => "0000000000111100",
4134 => "0000000000111100",
4135 => "0000000000111100",
4136 => "0000000000111100",
4137 => "0000000000111100",
4138 => "0000000000111100",
4139 => "0000000000111100",
4140 => "0000000000111100",
4141 => "0000000000111100",
4142 => "0000000000111100",
4143 => "0000000000111100",
4144 => "0000000000111100",
4145 => "0000000000111100",
4146 => "0000000000111100",
4147 => "0000000000111100",
4148 => "0000000000111100",
4149 => "0000000000111100",
4150 => "0000000000111100",
4151 => "0000000000111100",
4152 => "0000000000111100",
4153 => "0000000000111100",
4154 => "0000000000111100",
4155 => "0000000000111100",
4156 => "0000000000111100",
4157 => "0000000000111100",
4158 => "0000000000111100",
4159 => "0000000000111100",
4160 => "0000000000111100",
4161 => "0000000000111100",
4162 => "0000000000111100",
4163 => "0000000000111100",
4164 => "0000000000111100",
4165 => "0000000000111100",
4166 => "0000000000111100",
4167 => "0000000000111100",
4168 => "0000000000111100",
4169 => "0000000000111100",
4170 => "0000000000111100",
4171 => "0000000000111100",
4172 => "0000000000111100",
4173 => "0000000000111100",
4174 => "0000000000111100",
4175 => "0000000000111100",
4176 => "0000000000111100",
4177 => "0000000000111100",
4178 => "0000000000111100",
4179 => "0000000000111100",
4180 => "0000000000111100",
4181 => "0000000000111100",
4182 => "0000000000111100",
4183 => "0000000000111100",
4184 => "0000000000111101",
4185 => "0000000000111101",
4186 => "0000000000111101",
4187 => "0000000000111101",
4188 => "0000000000111101",
4189 => "0000000000111101",
4190 => "0000000000111101",
4191 => "0000000000111101",
4192 => "0000000000111101",
4193 => "0000000000111101",
4194 => "0000000000111101",
4195 => "0000000000111101",
4196 => "0000000000111101",
4197 => "0000000000111101",
4198 => "0000000000111101",
4199 => "0000000000111101",
4200 => "0000000000111101",
4201 => "0000000000111101",
4202 => "0000000000111101",
4203 => "0000000000111101",
4204 => "0000000000111101",
4205 => "0000000000111101",
4206 => "0000000000111101",
4207 => "0000000000111101",
4208 => "0000000000111101",
4209 => "0000000000111101",
4210 => "0000000000111101",
4211 => "0000000000111101",
4212 => "0000000000111101",
4213 => "0000000000111101",
4214 => "0000000000111101",
4215 => "0000000000111101",
4216 => "0000000000111101",
4217 => "0000000000111101",
4218 => "0000000000111101",
4219 => "0000000000111101",
4220 => "0000000000111101",
4221 => "0000000000111101",
4222 => "0000000000111101",
4223 => "0000000000111101",
4224 => "0000000000111101",
4225 => "0000000000111101",
4226 => "0000000000111101",
4227 => "0000000000111101",
4228 => "0000000000111101",
4229 => "0000000000111101",
4230 => "0000000000111101",
4231 => "0000000000111101",
4232 => "0000000000111101",
4233 => "0000000000111101",
4234 => "0000000000111101",
4235 => "0000000000111101",
4236 => "0000000000111101",
4237 => "0000000000111101",
4238 => "0000000000111101",
4239 => "0000000000111101",
4240 => "0000000000111101",
4241 => "0000000000111101",
4242 => "0000000000111101",
4243 => "0000000000111101",
4244 => "0000000000111101",
4245 => "0000000000111101",
4246 => "0000000000111101",
4247 => "0000000000111101",
4248 => "0000000000111101",
4249 => "0000000000111101",
4250 => "0000000000111101",
4251 => "0000000000111110",
4252 => "0000000000111110",
4253 => "0000000000111110",
4254 => "0000000000111110",
4255 => "0000000000111110",
4256 => "0000000000111110",
4257 => "0000000000111110",
4258 => "0000000000111110",
4259 => "0000000000111110",
4260 => "0000000000111110",
4261 => "0000000000111110",
4262 => "0000000000111110",
4263 => "0000000000111110",
4264 => "0000000000111110",
4265 => "0000000000111110",
4266 => "0000000000111110",
4267 => "0000000000111110",
4268 => "0000000000111110",
4269 => "0000000000111110",
4270 => "0000000000111110",
4271 => "0000000000111110",
4272 => "0000000000111110",
4273 => "0000000000111110",
4274 => "0000000000111110",
4275 => "0000000000111110",
4276 => "0000000000111110",
4277 => "0000000000111110",
4278 => "0000000000111110",
4279 => "0000000000111110",
4280 => "0000000000111110",
4281 => "0000000000111110",
4282 => "0000000000111110",
4283 => "0000000000111110",
4284 => "0000000000111110",
4285 => "0000000000111110",
4286 => "0000000000111110",
4287 => "0000000000111110",
4288 => "0000000000111110",
4289 => "0000000000111110",
4290 => "0000000000111110",
4291 => "0000000000111110",
4292 => "0000000000111110",
4293 => "0000000000111110",
4294 => "0000000000111110",
4295 => "0000000000111110",
4296 => "0000000000111110",
4297 => "0000000000111110",
4298 => "0000000000111110",
4299 => "0000000000111110",
4300 => "0000000000111110",
4301 => "0000000000111110",
4302 => "0000000000111110",
4303 => "0000000000111110",
4304 => "0000000000111110",
4305 => "0000000000111110",
4306 => "0000000000111110",
4307 => "0000000000111110",
4308 => "0000000000111110",
4309 => "0000000000111110",
4310 => "0000000000111110",
4311 => "0000000000111110",
4312 => "0000000000111110",
4313 => "0000000000111110",
4314 => "0000000000111110",
4315 => "0000000000111110",
4316 => "0000000000111110",
4317 => "0000000000111111",
4318 => "0000000000111111",
4319 => "0000000000111111",
4320 => "0000000000111111",
4321 => "0000000000111111",
4322 => "0000000000111111",
4323 => "0000000000111111",
4324 => "0000000000111111",
4325 => "0000000000111111",
4326 => "0000000000111111",
4327 => "0000000000111111",
4328 => "0000000000111111",
4329 => "0000000000111111",
4330 => "0000000000111111",
4331 => "0000000000111111",
4332 => "0000000000111111",
4333 => "0000000000111111",
4334 => "0000000000111111",
4335 => "0000000000111111",
4336 => "0000000000111111",
4337 => "0000000000111111",
4338 => "0000000000111111",
4339 => "0000000000111111",
4340 => "0000000000111111",
4341 => "0000000000111111",
4342 => "0000000000111111",
4343 => "0000000000111111",
4344 => "0000000000111111",
4345 => "0000000000111111",
4346 => "0000000000111111",
4347 => "0000000000111111",
4348 => "0000000000111111",
4349 => "0000000000111111",
4350 => "0000000000111111",
4351 => "0000000000111111",
4352 => "0000000000111111",
4353 => "0000000000111111",
4354 => "0000000000111111",
4355 => "0000000000111111",
4356 => "0000000000111111",
4357 => "0000000000111111",
4358 => "0000000000111111",
4359 => "0000000000111111",
4360 => "0000000000111111",
4361 => "0000000000111111",
4362 => "0000000000111111",
4363 => "0000000000111111",
4364 => "0000000000111111",
4365 => "0000000000111111",
4366 => "0000000000111111",
4367 => "0000000000111111",
4368 => "0000000000111111",
4369 => "0000000000111111",
4370 => "0000000000111111",
4371 => "0000000000111111",
4372 => "0000000000111111",
4373 => "0000000000111111",
4374 => "0000000000111111",
4375 => "0000000000111111",
4376 => "0000000000111111",
4377 => "0000000000111111",
4378 => "0000000000111111",
4379 => "0000000000111111",
4380 => "0000000000111111",
4381 => "0000000001000000",
4382 => "0000000001000000",
4383 => "0000000001000000",
4384 => "0000000001000000",
4385 => "0000000001000000",
4386 => "0000000001000000",
4387 => "0000000001000000",
4388 => "0000000001000000",
4389 => "0000000001000000",
4390 => "0000000001000000",
4391 => "0000000001000000",
4392 => "0000000001000000",
4393 => "0000000001000000",
4394 => "0000000001000000",
4395 => "0000000001000000",
4396 => "0000000001000000",
4397 => "0000000001000000",
4398 => "0000000001000000",
4399 => "0000000001000000",
4400 => "0000000001000000",
4401 => "0000000001000000",
4402 => "0000000001000000",
4403 => "0000000001000000",
4404 => "0000000001000000",
4405 => "0000000001000000",
4406 => "0000000001000000",
4407 => "0000000001000000",
4408 => "0000000001000000",
4409 => "0000000001000000",
4410 => "0000000001000000",
4411 => "0000000001000000",
4412 => "0000000001000000",
4413 => "0000000001000000",
4414 => "0000000001000000",
4415 => "0000000001000000",
4416 => "0000000001000000",
4417 => "0000000001000000",
4418 => "0000000001000000",
4419 => "0000000001000000",
4420 => "0000000001000000",
4421 => "0000000001000000",
4422 => "0000000001000000",
4423 => "0000000001000000",
4424 => "0000000001000000",
4425 => "0000000001000000",
4426 => "0000000001000000",
4427 => "0000000001000000",
4428 => "0000000001000000",
4429 => "0000000001000000",
4430 => "0000000001000000",
4431 => "0000000001000000",
4432 => "0000000001000000",
4433 => "0000000001000000",
4434 => "0000000001000000",
4435 => "0000000001000000",
4436 => "0000000001000000",
4437 => "0000000001000000",
4438 => "0000000001000000",
4439 => "0000000001000000",
4440 => "0000000001000000",
4441 => "0000000001000000",
4442 => "0000000001000000",
4443 => "0000000001000000",
4444 => "0000000001000000",
4445 => "0000000001000001",
4446 => "0000000001000001",
4447 => "0000000001000001",
4448 => "0000000001000001",
4449 => "0000000001000001",
4450 => "0000000001000001",
4451 => "0000000001000001",
4452 => "0000000001000001",
4453 => "0000000001000001",
4454 => "0000000001000001",
4455 => "0000000001000001",
4456 => "0000000001000001",
4457 => "0000000001000001",
4458 => "0000000001000001",
4459 => "0000000001000001",
4460 => "0000000001000001",
4461 => "0000000001000001",
4462 => "0000000001000001",
4463 => "0000000001000001",
4464 => "0000000001000001",
4465 => "0000000001000001",
4466 => "0000000001000001",
4467 => "0000000001000001",
4468 => "0000000001000001",
4469 => "0000000001000001",
4470 => "0000000001000001",
4471 => "0000000001000001",
4472 => "0000000001000001",
4473 => "0000000001000001",
4474 => "0000000001000001",
4475 => "0000000001000001",
4476 => "0000000001000001",
4477 => "0000000001000001",
4478 => "0000000001000001",
4479 => "0000000001000001",
4480 => "0000000001000001",
4481 => "0000000001000001",
4482 => "0000000001000001",
4483 => "0000000001000001",
4484 => "0000000001000001",
4485 => "0000000001000001",
4486 => "0000000001000001",
4487 => "0000000001000001",
4488 => "0000000001000001",
4489 => "0000000001000001",
4490 => "0000000001000001",
4491 => "0000000001000001",
4492 => "0000000001000001",
4493 => "0000000001000001",
4494 => "0000000001000001",
4495 => "0000000001000001",
4496 => "0000000001000001",
4497 => "0000000001000001",
4498 => "0000000001000001",
4499 => "0000000001000001",
4500 => "0000000001000001",
4501 => "0000000001000001",
4502 => "0000000001000001",
4503 => "0000000001000001",
4504 => "0000000001000001",
4505 => "0000000001000001",
4506 => "0000000001000001",
4507 => "0000000001000010",
4508 => "0000000001000010",
4509 => "0000000001000010",
4510 => "0000000001000010",
4511 => "0000000001000010",
4512 => "0000000001000010",
4513 => "0000000001000010",
4514 => "0000000001000010",
4515 => "0000000001000010",
4516 => "0000000001000010",
4517 => "0000000001000010",
4518 => "0000000001000010",
4519 => "0000000001000010",
4520 => "0000000001000010",
4521 => "0000000001000010",
4522 => "0000000001000010",
4523 => "0000000001000010",
4524 => "0000000001000010",
4525 => "0000000001000010",
4526 => "0000000001000010",
4527 => "0000000001000010",
4528 => "0000000001000010",
4529 => "0000000001000010",
4530 => "0000000001000010",
4531 => "0000000001000010",
4532 => "0000000001000010",
4533 => "0000000001000010",
4534 => "0000000001000010",
4535 => "0000000001000010",
4536 => "0000000001000010",
4537 => "0000000001000010",
4538 => "0000000001000010",
4539 => "0000000001000010",
4540 => "0000000001000010",
4541 => "0000000001000010",
4542 => "0000000001000010",
4543 => "0000000001000010",
4544 => "0000000001000010",
4545 => "0000000001000010",
4546 => "0000000001000010",
4547 => "0000000001000010",
4548 => "0000000001000010",
4549 => "0000000001000010",
4550 => "0000000001000010",
4551 => "0000000001000010",
4552 => "0000000001000010",
4553 => "0000000001000010",
4554 => "0000000001000010",
4555 => "0000000001000010",
4556 => "0000000001000010",
4557 => "0000000001000010",
4558 => "0000000001000010",
4559 => "0000000001000010",
4560 => "0000000001000010",
4561 => "0000000001000010",
4562 => "0000000001000010",
4563 => "0000000001000010",
4564 => "0000000001000010",
4565 => "0000000001000010",
4566 => "0000000001000010",
4567 => "0000000001000010",
4568 => "0000000001000010",
4569 => "0000000001000011",
4570 => "0000000001000011",
4571 => "0000000001000011",
4572 => "0000000001000011",
4573 => "0000000001000011",
4574 => "0000000001000011",
4575 => "0000000001000011",
4576 => "0000000001000011",
4577 => "0000000001000011",
4578 => "0000000001000011",
4579 => "0000000001000011",
4580 => "0000000001000011",
4581 => "0000000001000011",
4582 => "0000000001000011",
4583 => "0000000001000011",
4584 => "0000000001000011",
4585 => "0000000001000011",
4586 => "0000000001000011",
4587 => "0000000001000011",
4588 => "0000000001000011",
4589 => "0000000001000011",
4590 => "0000000001000011",
4591 => "0000000001000011",
4592 => "0000000001000011",
4593 => "0000000001000011",
4594 => "0000000001000011",
4595 => "0000000001000011",
4596 => "0000000001000011",
4597 => "0000000001000011",
4598 => "0000000001000011",
4599 => "0000000001000011",
4600 => "0000000001000011",
4601 => "0000000001000011",
4602 => "0000000001000011",
4603 => "0000000001000011",
4604 => "0000000001000011",
4605 => "0000000001000011",
4606 => "0000000001000011",
4607 => "0000000001000011",
4608 => "0000000001000011",
4609 => "0000000001000011",
4610 => "0000000001000011",
4611 => "0000000001000011",
4612 => "0000000001000011",
4613 => "0000000001000011",
4614 => "0000000001000011",
4615 => "0000000001000011",
4616 => "0000000001000011",
4617 => "0000000001000011",
4618 => "0000000001000011",
4619 => "0000000001000011",
4620 => "0000000001000011",
4621 => "0000000001000011",
4622 => "0000000001000011",
4623 => "0000000001000011",
4624 => "0000000001000011",
4625 => "0000000001000011",
4626 => "0000000001000011",
4627 => "0000000001000011",
4628 => "0000000001000011",
4629 => "0000000001000011",
4630 => "0000000001000100",
4631 => "0000000001000100",
4632 => "0000000001000100",
4633 => "0000000001000100",
4634 => "0000000001000100",
4635 => "0000000001000100",
4636 => "0000000001000100",
4637 => "0000000001000100",
4638 => "0000000001000100",
4639 => "0000000001000100",
4640 => "0000000001000100",
4641 => "0000000001000100",
4642 => "0000000001000100",
4643 => "0000000001000100",
4644 => "0000000001000100",
4645 => "0000000001000100",
4646 => "0000000001000100",
4647 => "0000000001000100",
4648 => "0000000001000100",
4649 => "0000000001000100",
4650 => "0000000001000100",
4651 => "0000000001000100",
4652 => "0000000001000100",
4653 => "0000000001000100",
4654 => "0000000001000100",
4655 => "0000000001000100",
4656 => "0000000001000100",
4657 => "0000000001000100",
4658 => "0000000001000100",
4659 => "0000000001000100",
4660 => "0000000001000100",
4661 => "0000000001000100",
4662 => "0000000001000100",
4663 => "0000000001000100",
4664 => "0000000001000100",
4665 => "0000000001000100",
4666 => "0000000001000100",
4667 => "0000000001000100",
4668 => "0000000001000100",
4669 => "0000000001000100",
4670 => "0000000001000100",
4671 => "0000000001000100",
4672 => "0000000001000100",
4673 => "0000000001000100",
4674 => "0000000001000100",
4675 => "0000000001000100",
4676 => "0000000001000100",
4677 => "0000000001000100",
4678 => "0000000001000100",
4679 => "0000000001000100",
4680 => "0000000001000100",
4681 => "0000000001000100",
4682 => "0000000001000100",
4683 => "0000000001000100",
4684 => "0000000001000100",
4685 => "0000000001000100",
4686 => "0000000001000100",
4687 => "0000000001000100",
4688 => "0000000001000100",
4689 => "0000000001000100",
4690 => "0000000001000101",
4691 => "0000000001000101",
4692 => "0000000001000101",
4693 => "0000000001000101",
4694 => "0000000001000101",
4695 => "0000000001000101",
4696 => "0000000001000101",
4697 => "0000000001000101",
4698 => "0000000001000101",
4699 => "0000000001000101",
4700 => "0000000001000101",
4701 => "0000000001000101",
4702 => "0000000001000101",
4703 => "0000000001000101",
4704 => "0000000001000101",
4705 => "0000000001000101",
4706 => "0000000001000101",
4707 => "0000000001000101",
4708 => "0000000001000101",
4709 => "0000000001000101",
4710 => "0000000001000101",
4711 => "0000000001000101",
4712 => "0000000001000101",
4713 => "0000000001000101",
4714 => "0000000001000101",
4715 => "0000000001000101",
4716 => "0000000001000101",
4717 => "0000000001000101",
4718 => "0000000001000101",
4719 => "0000000001000101",
4720 => "0000000001000101",
4721 => "0000000001000101",
4722 => "0000000001000101",
4723 => "0000000001000101",
4724 => "0000000001000101",
4725 => "0000000001000101",
4726 => "0000000001000101",
4727 => "0000000001000101",
4728 => "0000000001000101",
4729 => "0000000001000101",
4730 => "0000000001000101",
4731 => "0000000001000101",
4732 => "0000000001000101",
4733 => "0000000001000101",
4734 => "0000000001000101",
4735 => "0000000001000101",
4736 => "0000000001000101",
4737 => "0000000001000101",
4738 => "0000000001000101",
4739 => "0000000001000101",
4740 => "0000000001000101",
4741 => "0000000001000101",
4742 => "0000000001000101",
4743 => "0000000001000101",
4744 => "0000000001000101",
4745 => "0000000001000101",
4746 => "0000000001000101",
4747 => "0000000001000101",
4748 => "0000000001000101",
4749 => "0000000001000110",
4750 => "0000000001000110",
4751 => "0000000001000110",
4752 => "0000000001000110",
4753 => "0000000001000110",
4754 => "0000000001000110",
4755 => "0000000001000110",
4756 => "0000000001000110",
4757 => "0000000001000110",
4758 => "0000000001000110",
4759 => "0000000001000110",
4760 => "0000000001000110",
4761 => "0000000001000110",
4762 => "0000000001000110",
4763 => "0000000001000110",
4764 => "0000000001000110",
4765 => "0000000001000110",
4766 => "0000000001000110",
4767 => "0000000001000110",
4768 => "0000000001000110",
4769 => "0000000001000110",
4770 => "0000000001000110",
4771 => "0000000001000110",
4772 => "0000000001000110",
4773 => "0000000001000110",
4774 => "0000000001000110",
4775 => "0000000001000110",
4776 => "0000000001000110",
4777 => "0000000001000110",
4778 => "0000000001000110",
4779 => "0000000001000110",
4780 => "0000000001000110",
4781 => "0000000001000110",
4782 => "0000000001000110",
4783 => "0000000001000110",
4784 => "0000000001000110",
4785 => "0000000001000110",
4786 => "0000000001000110",
4787 => "0000000001000110",
4788 => "0000000001000110",
4789 => "0000000001000110",
4790 => "0000000001000110",
4791 => "0000000001000110",
4792 => "0000000001000110",
4793 => "0000000001000110",
4794 => "0000000001000110",
4795 => "0000000001000110",
4796 => "0000000001000110",
4797 => "0000000001000110",
4798 => "0000000001000110",
4799 => "0000000001000110",
4800 => "0000000001000110",
4801 => "0000000001000110",
4802 => "0000000001000110",
4803 => "0000000001000110",
4804 => "0000000001000110",
4805 => "0000000001000110",
4806 => "0000000001000110",
4807 => "0000000001000111",
4808 => "0000000001000111",
4809 => "0000000001000111",
4810 => "0000000001000111",
4811 => "0000000001000111",
4812 => "0000000001000111",
4813 => "0000000001000111",
4814 => "0000000001000111",
4815 => "0000000001000111",
4816 => "0000000001000111",
4817 => "0000000001000111",
4818 => "0000000001000111",
4819 => "0000000001000111",
4820 => "0000000001000111",
4821 => "0000000001000111",
4822 => "0000000001000111",
4823 => "0000000001000111",
4824 => "0000000001000111",
4825 => "0000000001000111",
4826 => "0000000001000111",
4827 => "0000000001000111",
4828 => "0000000001000111",
4829 => "0000000001000111",
4830 => "0000000001000111",
4831 => "0000000001000111",
4832 => "0000000001000111",
4833 => "0000000001000111",
4834 => "0000000001000111",
4835 => "0000000001000111",
4836 => "0000000001000111",
4837 => "0000000001000111",
4838 => "0000000001000111",
4839 => "0000000001000111",
4840 => "0000000001000111",
4841 => "0000000001000111",
4842 => "0000000001000111",
4843 => "0000000001000111",
4844 => "0000000001000111",
4845 => "0000000001000111",
4846 => "0000000001000111",
4847 => "0000000001000111",
4848 => "0000000001000111",
4849 => "0000000001000111",
4850 => "0000000001000111",
4851 => "0000000001000111",
4852 => "0000000001000111",
4853 => "0000000001000111",
4854 => "0000000001000111",
4855 => "0000000001000111",
4856 => "0000000001000111",
4857 => "0000000001000111",
4858 => "0000000001000111",
4859 => "0000000001000111",
4860 => "0000000001000111",
4861 => "0000000001000111",
4862 => "0000000001000111",
4863 => "0000000001000111",
4864 => "0000000001001000",
4865 => "0000000001001000",
4866 => "0000000001001000",
4867 => "0000000001001000",
4868 => "0000000001001000",
4869 => "0000000001001000",
4870 => "0000000001001000",
4871 => "0000000001001000",
4872 => "0000000001001000",
4873 => "0000000001001000",
4874 => "0000000001001000",
4875 => "0000000001001000",
4876 => "0000000001001000",
4877 => "0000000001001000",
4878 => "0000000001001000",
4879 => "0000000001001000",
4880 => "0000000001001000",
4881 => "0000000001001000",
4882 => "0000000001001000",
4883 => "0000000001001000",
4884 => "0000000001001000",
4885 => "0000000001001000",
4886 => "0000000001001000",
4887 => "0000000001001000",
4888 => "0000000001001000",
4889 => "0000000001001000",
4890 => "0000000001001000",
4891 => "0000000001001000",
4892 => "0000000001001000",
4893 => "0000000001001000",
4894 => "0000000001001000",
4895 => "0000000001001000",
4896 => "0000000001001000",
4897 => "0000000001001000",
4898 => "0000000001001000",
4899 => "0000000001001000",
4900 => "0000000001001000",
4901 => "0000000001001000",
4902 => "0000000001001000",
4903 => "0000000001001000",
4904 => "0000000001001000",
4905 => "0000000001001000",
4906 => "0000000001001000",
4907 => "0000000001001000",
4908 => "0000000001001000",
4909 => "0000000001001000",
4910 => "0000000001001000",
4911 => "0000000001001000",
4912 => "0000000001001000",
4913 => "0000000001001000",
4914 => "0000000001001000",
4915 => "0000000001001000",
4916 => "0000000001001000",
4917 => "0000000001001000",
4918 => "0000000001001000",
4919 => "0000000001001000",
4920 => "0000000001001000",
4921 => "0000000001001001",
4922 => "0000000001001001",
4923 => "0000000001001001",
4924 => "0000000001001001",
4925 => "0000000001001001",
4926 => "0000000001001001",
4927 => "0000000001001001",
4928 => "0000000001001001",
4929 => "0000000001001001",
4930 => "0000000001001001",
4931 => "0000000001001001",
4932 => "0000000001001001",
4933 => "0000000001001001",
4934 => "0000000001001001",
4935 => "0000000001001001",
4936 => "0000000001001001",
4937 => "0000000001001001",
4938 => "0000000001001001",
4939 => "0000000001001001",
4940 => "0000000001001001",
4941 => "0000000001001001",
4942 => "0000000001001001",
4943 => "0000000001001001",
4944 => "0000000001001001",
4945 => "0000000001001001",
4946 => "0000000001001001",
4947 => "0000000001001001",
4948 => "0000000001001001",
4949 => "0000000001001001",
4950 => "0000000001001001",
4951 => "0000000001001001",
4952 => "0000000001001001",
4953 => "0000000001001001",
4954 => "0000000001001001",
4955 => "0000000001001001",
4956 => "0000000001001001",
4957 => "0000000001001001",
4958 => "0000000001001001",
4959 => "0000000001001001",
4960 => "0000000001001001",
4961 => "0000000001001001",
4962 => "0000000001001001",
4963 => "0000000001001001",
4964 => "0000000001001001",
4965 => "0000000001001001",
4966 => "0000000001001001",
4967 => "0000000001001001",
4968 => "0000000001001001",
4969 => "0000000001001001",
4970 => "0000000001001001",
4971 => "0000000001001001",
4972 => "0000000001001001",
4973 => "0000000001001001",
4974 => "0000000001001001",
4975 => "0000000001001001",
4976 => "0000000001001010",
4977 => "0000000001001010",
4978 => "0000000001001010",
4979 => "0000000001001010",
4980 => "0000000001001010",
4981 => "0000000001001010",
4982 => "0000000001001010",
4983 => "0000000001001010",
4984 => "0000000001001010",
4985 => "0000000001001010",
4986 => "0000000001001010",
4987 => "0000000001001010",
4988 => "0000000001001010",
4989 => "0000000001001010",
4990 => "0000000001001010",
4991 => "0000000001001010",
4992 => "0000000001001010",
4993 => "0000000001001010",
4994 => "0000000001001010",
4995 => "0000000001001010",
4996 => "0000000001001010",
4997 => "0000000001001010",
4998 => "0000000001001010",
4999 => "0000000001001010",
5000 => "0000000001001010",
5001 => "0000000001001010",
5002 => "0000000001001010",
5003 => "0000000001001010",
5004 => "0000000001001010",
5005 => "0000000001001010",
5006 => "0000000001001010",
5007 => "0000000001001010",
5008 => "0000000001001010",
5009 => "0000000001001010",
5010 => "0000000001001010",
5011 => "0000000001001010",
5012 => "0000000001001010",
5013 => "0000000001001010",
5014 => "0000000001001010",
5015 => "0000000001001010",
5016 => "0000000001001010",
5017 => "0000000001001010",
5018 => "0000000001001010",
5019 => "0000000001001010",
5020 => "0000000001001010",
5021 => "0000000001001010",
5022 => "0000000001001010",
5023 => "0000000001001010",
5024 => "0000000001001010",
5025 => "0000000001001010",
5026 => "0000000001001010",
5027 => "0000000001001010",
5028 => "0000000001001010",
5029 => "0000000001001010",
5030 => "0000000001001010",
5031 => "0000000001001011",
5032 => "0000000001001011",
5033 => "0000000001001011",
5034 => "0000000001001011",
5035 => "0000000001001011",
5036 => "0000000001001011",
5037 => "0000000001001011",
5038 => "0000000001001011",
5039 => "0000000001001011",
5040 => "0000000001001011",
5041 => "0000000001001011",
5042 => "0000000001001011",
5043 => "0000000001001011",
5044 => "0000000001001011",
5045 => "0000000001001011",
5046 => "0000000001001011",
5047 => "0000000001001011",
5048 => "0000000001001011",
5049 => "0000000001001011",
5050 => "0000000001001011",
5051 => "0000000001001011",
5052 => "0000000001001011",
5053 => "0000000001001011",
5054 => "0000000001001011",
5055 => "0000000001001011",
5056 => "0000000001001011",
5057 => "0000000001001011",
5058 => "0000000001001011",
5059 => "0000000001001011",
5060 => "0000000001001011",
5061 => "0000000001001011",
5062 => "0000000001001011",
5063 => "0000000001001011",
5064 => "0000000001001011",
5065 => "0000000001001011",
5066 => "0000000001001011",
5067 => "0000000001001011",
5068 => "0000000001001011",
5069 => "0000000001001011",
5070 => "0000000001001011",
5071 => "0000000001001011",
5072 => "0000000001001011",
5073 => "0000000001001011",
5074 => "0000000001001011",
5075 => "0000000001001011",
5076 => "0000000001001011",
5077 => "0000000001001011",
5078 => "0000000001001011",
5079 => "0000000001001011",
5080 => "0000000001001011",
5081 => "0000000001001011",
5082 => "0000000001001011",
5083 => "0000000001001011",
5084 => "0000000001001011",
5085 => "0000000001001011",
5086 => "0000000001001100",
5087 => "0000000001001100",
5088 => "0000000001001100",
5089 => "0000000001001100",
5090 => "0000000001001100",
5091 => "0000000001001100",
5092 => "0000000001001100",
5093 => "0000000001001100",
5094 => "0000000001001100",
5095 => "0000000001001100",
5096 => "0000000001001100",
5097 => "0000000001001100",
5098 => "0000000001001100",
5099 => "0000000001001100",
5100 => "0000000001001100",
5101 => "0000000001001100",
5102 => "0000000001001100",
5103 => "0000000001001100",
5104 => "0000000001001100",
5105 => "0000000001001100",
5106 => "0000000001001100",
5107 => "0000000001001100",
5108 => "0000000001001100",
5109 => "0000000001001100",
5110 => "0000000001001100",
5111 => "0000000001001100",
5112 => "0000000001001100",
5113 => "0000000001001100",
5114 => "0000000001001100",
5115 => "0000000001001100",
5116 => "0000000001001100",
5117 => "0000000001001100",
5118 => "0000000001001100",
5119 => "0000000001001100",
5120 => "0000000001001100",
5121 => "0000000001001100",
5122 => "0000000001001100",
5123 => "0000000001001100",
5124 => "0000000001001100",
5125 => "0000000001001100",
5126 => "0000000001001100",
5127 => "0000000001001100",
5128 => "0000000001001100",
5129 => "0000000001001100",
5130 => "0000000001001100",
5131 => "0000000001001100",
5132 => "0000000001001100",
5133 => "0000000001001100",
5134 => "0000000001001100",
5135 => "0000000001001100",
5136 => "0000000001001100",
5137 => "0000000001001100",
5138 => "0000000001001100",
5139 => "0000000001001101",
5140 => "0000000001001101",
5141 => "0000000001001101",
5142 => "0000000001001101",
5143 => "0000000001001101",
5144 => "0000000001001101",
5145 => "0000000001001101",
5146 => "0000000001001101",
5147 => "0000000001001101",
5148 => "0000000001001101",
5149 => "0000000001001101",
5150 => "0000000001001101",
5151 => "0000000001001101",
5152 => "0000000001001101",
5153 => "0000000001001101",
5154 => "0000000001001101",
5155 => "0000000001001101",
5156 => "0000000001001101",
5157 => "0000000001001101",
5158 => "0000000001001101",
5159 => "0000000001001101",
5160 => "0000000001001101",
5161 => "0000000001001101",
5162 => "0000000001001101",
5163 => "0000000001001101",
5164 => "0000000001001101",
5165 => "0000000001001101",
5166 => "0000000001001101",
5167 => "0000000001001101",
5168 => "0000000001001101",
5169 => "0000000001001101",
5170 => "0000000001001101",
5171 => "0000000001001101",
5172 => "0000000001001101",
5173 => "0000000001001101",
5174 => "0000000001001101",
5175 => "0000000001001101",
5176 => "0000000001001101",
5177 => "0000000001001101",
5178 => "0000000001001101",
5179 => "0000000001001101",
5180 => "0000000001001101",
5181 => "0000000001001101",
5182 => "0000000001001101",
5183 => "0000000001001101",
5184 => "0000000001001101",
5185 => "0000000001001101",
5186 => "0000000001001101",
5187 => "0000000001001101",
5188 => "0000000001001101",
5189 => "0000000001001101",
5190 => "0000000001001101",
5191 => "0000000001001101",
5192 => "0000000001001110",
5193 => "0000000001001110",
5194 => "0000000001001110",
5195 => "0000000001001110",
5196 => "0000000001001110",
5197 => "0000000001001110",
5198 => "0000000001001110",
5199 => "0000000001001110",
5200 => "0000000001001110",
5201 => "0000000001001110",
5202 => "0000000001001110",
5203 => "0000000001001110",
5204 => "0000000001001110",
5205 => "0000000001001110",
5206 => "0000000001001110",
5207 => "0000000001001110",
5208 => "0000000001001110",
5209 => "0000000001001110",
5210 => "0000000001001110",
5211 => "0000000001001110",
5212 => "0000000001001110",
5213 => "0000000001001110",
5214 => "0000000001001110",
5215 => "0000000001001110",
5216 => "0000000001001110",
5217 => "0000000001001110",
5218 => "0000000001001110",
5219 => "0000000001001110",
5220 => "0000000001001110",
5221 => "0000000001001110",
5222 => "0000000001001110",
5223 => "0000000001001110",
5224 => "0000000001001110",
5225 => "0000000001001110",
5226 => "0000000001001110",
5227 => "0000000001001110",
5228 => "0000000001001110",
5229 => "0000000001001110",
5230 => "0000000001001110",
5231 => "0000000001001110",
5232 => "0000000001001110",
5233 => "0000000001001110",
5234 => "0000000001001110",
5235 => "0000000001001110",
5236 => "0000000001001110",
5237 => "0000000001001110",
5238 => "0000000001001110",
5239 => "0000000001001110",
5240 => "0000000001001110",
5241 => "0000000001001110",
5242 => "0000000001001110",
5243 => "0000000001001110",
5244 => "0000000001001110",
5245 => "0000000001001111",
5246 => "0000000001001111",
5247 => "0000000001001111",
5248 => "0000000001001111",
5249 => "0000000001001111",
5250 => "0000000001001111",
5251 => "0000000001001111",
5252 => "0000000001001111",
5253 => "0000000001001111",
5254 => "0000000001001111",
5255 => "0000000001001111",
5256 => "0000000001001111",
5257 => "0000000001001111",
5258 => "0000000001001111",
5259 => "0000000001001111",
5260 => "0000000001001111",
5261 => "0000000001001111",
5262 => "0000000001001111",
5263 => "0000000001001111",
5264 => "0000000001001111",
5265 => "0000000001001111",
5266 => "0000000001001111",
5267 => "0000000001001111",
5268 => "0000000001001111",
5269 => "0000000001001111",
5270 => "0000000001001111",
5271 => "0000000001001111",
5272 => "0000000001001111",
5273 => "0000000001001111",
5274 => "0000000001001111",
5275 => "0000000001001111",
5276 => "0000000001001111",
5277 => "0000000001001111",
5278 => "0000000001001111",
5279 => "0000000001001111",
5280 => "0000000001001111",
5281 => "0000000001001111",
5282 => "0000000001001111",
5283 => "0000000001001111",
5284 => "0000000001001111",
5285 => "0000000001001111",
5286 => "0000000001001111",
5287 => "0000000001001111",
5288 => "0000000001001111",
5289 => "0000000001001111",
5290 => "0000000001001111",
5291 => "0000000001001111",
5292 => "0000000001001111",
5293 => "0000000001001111",
5294 => "0000000001001111",
5295 => "0000000001001111",
5296 => "0000000001010000",
5297 => "0000000001010000",
5298 => "0000000001010000",
5299 => "0000000001010000",
5300 => "0000000001010000",
5301 => "0000000001010000",
5302 => "0000000001010000",
5303 => "0000000001010000",
5304 => "0000000001010000",
5305 => "0000000001010000",
5306 => "0000000001010000",
5307 => "0000000001010000",
5308 => "0000000001010000",
5309 => "0000000001010000",
5310 => "0000000001010000",
5311 => "0000000001010000",
5312 => "0000000001010000",
5313 => "0000000001010000",
5314 => "0000000001010000",
5315 => "0000000001010000",
5316 => "0000000001010000",
5317 => "0000000001010000",
5318 => "0000000001010000",
5319 => "0000000001010000",
5320 => "0000000001010000",
5321 => "0000000001010000",
5322 => "0000000001010000",
5323 => "0000000001010000",
5324 => "0000000001010000",
5325 => "0000000001010000",
5326 => "0000000001010000",
5327 => "0000000001010000",
5328 => "0000000001010000",
5329 => "0000000001010000",
5330 => "0000000001010000",
5331 => "0000000001010000",
5332 => "0000000001010000",
5333 => "0000000001010000",
5334 => "0000000001010000",
5335 => "0000000001010000",
5336 => "0000000001010000",
5337 => "0000000001010000",
5338 => "0000000001010000",
5339 => "0000000001010000",
5340 => "0000000001010000",
5341 => "0000000001010000",
5342 => "0000000001010000",
5343 => "0000000001010000",
5344 => "0000000001010000",
5345 => "0000000001010000",
5346 => "0000000001010000",
5347 => "0000000001010001",
5348 => "0000000001010001",
5349 => "0000000001010001",
5350 => "0000000001010001",
5351 => "0000000001010001",
5352 => "0000000001010001",
5353 => "0000000001010001",
5354 => "0000000001010001",
5355 => "0000000001010001",
5356 => "0000000001010001",
5357 => "0000000001010001",
5358 => "0000000001010001",
5359 => "0000000001010001",
5360 => "0000000001010001",
5361 => "0000000001010001",
5362 => "0000000001010001",
5363 => "0000000001010001",
5364 => "0000000001010001",
5365 => "0000000001010001",
5366 => "0000000001010001",
5367 => "0000000001010001",
5368 => "0000000001010001",
5369 => "0000000001010001",
5370 => "0000000001010001",
5371 => "0000000001010001",
5372 => "0000000001010001",
5373 => "0000000001010001",
5374 => "0000000001010001",
5375 => "0000000001010001",
5376 => "0000000001010001",
5377 => "0000000001010001",
5378 => "0000000001010001",
5379 => "0000000001010001",
5380 => "0000000001010001",
5381 => "0000000001010001",
5382 => "0000000001010001",
5383 => "0000000001010001",
5384 => "0000000001010001",
5385 => "0000000001010001",
5386 => "0000000001010001",
5387 => "0000000001010001",
5388 => "0000000001010001",
5389 => "0000000001010001",
5390 => "0000000001010001",
5391 => "0000000001010001",
5392 => "0000000001010001",
5393 => "0000000001010001",
5394 => "0000000001010001",
5395 => "0000000001010001",
5396 => "0000000001010001",
5397 => "0000000001010010",
5398 => "0000000001010010",
5399 => "0000000001010010",
5400 => "0000000001010010",
5401 => "0000000001010010",
5402 => "0000000001010010",
5403 => "0000000001010010",
5404 => "0000000001010010",
5405 => "0000000001010010",
5406 => "0000000001010010",
5407 => "0000000001010010",
5408 => "0000000001010010",
5409 => "0000000001010010",
5410 => "0000000001010010",
5411 => "0000000001010010",
5412 => "0000000001010010",
5413 => "0000000001010010",
5414 => "0000000001010010",
5415 => "0000000001010010",
5416 => "0000000001010010",
5417 => "0000000001010010",
5418 => "0000000001010010",
5419 => "0000000001010010",
5420 => "0000000001010010",
5421 => "0000000001010010",
5422 => "0000000001010010",
5423 => "0000000001010010",
5424 => "0000000001010010",
5425 => "0000000001010010",
5426 => "0000000001010010",
5427 => "0000000001010010",
5428 => "0000000001010010",
5429 => "0000000001010010",
5430 => "0000000001010010",
5431 => "0000000001010010",
5432 => "0000000001010010",
5433 => "0000000001010010",
5434 => "0000000001010010",
5435 => "0000000001010010",
5436 => "0000000001010010",
5437 => "0000000001010010",
5438 => "0000000001010010",
5439 => "0000000001010010",
5440 => "0000000001010010",
5441 => "0000000001010010",
5442 => "0000000001010010",
5443 => "0000000001010010",
5444 => "0000000001010010",
5445 => "0000000001010010",
5446 => "0000000001010010",
5447 => "0000000001010011",
5448 => "0000000001010011",
5449 => "0000000001010011",
5450 => "0000000001010011",
5451 => "0000000001010011",
5452 => "0000000001010011",
5453 => "0000000001010011",
5454 => "0000000001010011",
5455 => "0000000001010011",
5456 => "0000000001010011",
5457 => "0000000001010011",
5458 => "0000000001010011",
5459 => "0000000001010011",
5460 => "0000000001010011",
5461 => "0000000001010011",
5462 => "0000000001010011",
5463 => "0000000001010011",
5464 => "0000000001010011",
5465 => "0000000001010011",
5466 => "0000000001010011",
5467 => "0000000001010011",
5468 => "0000000001010011",
5469 => "0000000001010011",
5470 => "0000000001010011",
5471 => "0000000001010011",
5472 => "0000000001010011",
5473 => "0000000001010011",
5474 => "0000000001010011",
5475 => "0000000001010011",
5476 => "0000000001010011",
5477 => "0000000001010011",
5478 => "0000000001010011",
5479 => "0000000001010011",
5480 => "0000000001010011",
5481 => "0000000001010011",
5482 => "0000000001010011",
5483 => "0000000001010011",
5484 => "0000000001010011",
5485 => "0000000001010011",
5486 => "0000000001010011",
5487 => "0000000001010011",
5488 => "0000000001010011",
5489 => "0000000001010011",
5490 => "0000000001010011",
5491 => "0000000001010011",
5492 => "0000000001010011",
5493 => "0000000001010011",
5494 => "0000000001010011",
5495 => "0000000001010011",
5496 => "0000000001010100",
5497 => "0000000001010100",
5498 => "0000000001010100",
5499 => "0000000001010100",
5500 => "0000000001010100",
5501 => "0000000001010100",
5502 => "0000000001010100",
5503 => "0000000001010100",
5504 => "0000000001010100",
5505 => "0000000001010100",
5506 => "0000000001010100",
5507 => "0000000001010100",
5508 => "0000000001010100",
5509 => "0000000001010100",
5510 => "0000000001010100",
5511 => "0000000001010100",
5512 => "0000000001010100",
5513 => "0000000001010100",
5514 => "0000000001010100",
5515 => "0000000001010100",
5516 => "0000000001010100",
5517 => "0000000001010100",
5518 => "0000000001010100",
5519 => "0000000001010100",
5520 => "0000000001010100",
5521 => "0000000001010100",
5522 => "0000000001010100",
5523 => "0000000001010100",
5524 => "0000000001010100",
5525 => "0000000001010100",
5526 => "0000000001010100",
5527 => "0000000001010100",
5528 => "0000000001010100",
5529 => "0000000001010100",
5530 => "0000000001010100",
5531 => "0000000001010100",
5532 => "0000000001010100",
5533 => "0000000001010100",
5534 => "0000000001010100",
5535 => "0000000001010100",
5536 => "0000000001010100",
5537 => "0000000001010100",
5538 => "0000000001010100",
5539 => "0000000001010100",
5540 => "0000000001010100",
5541 => "0000000001010100",
5542 => "0000000001010100",
5543 => "0000000001010100",
5544 => "0000000001010100",
5545 => "0000000001010101",
5546 => "0000000001010101",
5547 => "0000000001010101",
5548 => "0000000001010101",
5549 => "0000000001010101",
5550 => "0000000001010101",
5551 => "0000000001010101",
5552 => "0000000001010101",
5553 => "0000000001010101",
5554 => "0000000001010101",
5555 => "0000000001010101",
5556 => "0000000001010101",
5557 => "0000000001010101",
5558 => "0000000001010101",
5559 => "0000000001010101",
5560 => "0000000001010101",
5561 => "0000000001010101",
5562 => "0000000001010101",
5563 => "0000000001010101",
5564 => "0000000001010101",
5565 => "0000000001010101",
5566 => "0000000001010101",
5567 => "0000000001010101",
5568 => "0000000001010101",
5569 => "0000000001010101",
5570 => "0000000001010101",
5571 => "0000000001010101",
5572 => "0000000001010101",
5573 => "0000000001010101",
5574 => "0000000001010101",
5575 => "0000000001010101",
5576 => "0000000001010101",
5577 => "0000000001010101",
5578 => "0000000001010101",
5579 => "0000000001010101",
5580 => "0000000001010101",
5581 => "0000000001010101",
5582 => "0000000001010101",
5583 => "0000000001010101",
5584 => "0000000001010101",
5585 => "0000000001010101",
5586 => "0000000001010101",
5587 => "0000000001010101",
5588 => "0000000001010101",
5589 => "0000000001010101",
5590 => "0000000001010101",
5591 => "0000000001010101",
5592 => "0000000001010101",
5593 => "0000000001010110",
5594 => "0000000001010110",
5595 => "0000000001010110",
5596 => "0000000001010110",
5597 => "0000000001010110",
5598 => "0000000001010110",
5599 => "0000000001010110",
5600 => "0000000001010110",
5601 => "0000000001010110",
5602 => "0000000001010110",
5603 => "0000000001010110",
5604 => "0000000001010110",
5605 => "0000000001010110",
5606 => "0000000001010110",
5607 => "0000000001010110",
5608 => "0000000001010110",
5609 => "0000000001010110",
5610 => "0000000001010110",
5611 => "0000000001010110",
5612 => "0000000001010110",
5613 => "0000000001010110",
5614 => "0000000001010110",
5615 => "0000000001010110",
5616 => "0000000001010110",
5617 => "0000000001010110",
5618 => "0000000001010110",
5619 => "0000000001010110",
5620 => "0000000001010110",
5621 => "0000000001010110",
5622 => "0000000001010110",
5623 => "0000000001010110",
5624 => "0000000001010110",
5625 => "0000000001010110",
5626 => "0000000001010110",
5627 => "0000000001010110",
5628 => "0000000001010110",
5629 => "0000000001010110",
5630 => "0000000001010110",
5631 => "0000000001010110",
5632 => "0000000001010110",
5633 => "0000000001010110",
5634 => "0000000001010110",
5635 => "0000000001010110",
5636 => "0000000001010110",
5637 => "0000000001010110",
5638 => "0000000001010110",
5639 => "0000000001010110",
5640 => "0000000001010111",
5641 => "0000000001010111",
5642 => "0000000001010111",
5643 => "0000000001010111",
5644 => "0000000001010111",
5645 => "0000000001010111",
5646 => "0000000001010111",
5647 => "0000000001010111",
5648 => "0000000001010111",
5649 => "0000000001010111",
5650 => "0000000001010111",
5651 => "0000000001010111",
5652 => "0000000001010111",
5653 => "0000000001010111",
5654 => "0000000001010111",
5655 => "0000000001010111",
5656 => "0000000001010111",
5657 => "0000000001010111",
5658 => "0000000001010111",
5659 => "0000000001010111",
5660 => "0000000001010111",
5661 => "0000000001010111",
5662 => "0000000001010111",
5663 => "0000000001010111",
5664 => "0000000001010111",
5665 => "0000000001010111",
5666 => "0000000001010111",
5667 => "0000000001010111",
5668 => "0000000001010111",
5669 => "0000000001010111",
5670 => "0000000001010111",
5671 => "0000000001010111",
5672 => "0000000001010111",
5673 => "0000000001010111",
5674 => "0000000001010111",
5675 => "0000000001010111",
5676 => "0000000001010111",
5677 => "0000000001010111",
5678 => "0000000001010111",
5679 => "0000000001010111",
5680 => "0000000001010111",
5681 => "0000000001010111",
5682 => "0000000001010111",
5683 => "0000000001010111",
5684 => "0000000001010111",
5685 => "0000000001010111",
5686 => "0000000001010111",
5687 => "0000000001011000",
5688 => "0000000001011000",
5689 => "0000000001011000",
5690 => "0000000001011000",
5691 => "0000000001011000",
5692 => "0000000001011000",
5693 => "0000000001011000",
5694 => "0000000001011000",
5695 => "0000000001011000",
5696 => "0000000001011000",
5697 => "0000000001011000",
5698 => "0000000001011000",
5699 => "0000000001011000",
5700 => "0000000001011000",
5701 => "0000000001011000",
5702 => "0000000001011000",
5703 => "0000000001011000",
5704 => "0000000001011000",
5705 => "0000000001011000",
5706 => "0000000001011000",
5707 => "0000000001011000",
5708 => "0000000001011000",
5709 => "0000000001011000",
5710 => "0000000001011000",
5711 => "0000000001011000",
5712 => "0000000001011000",
5713 => "0000000001011000",
5714 => "0000000001011000",
5715 => "0000000001011000",
5716 => "0000000001011000",
5717 => "0000000001011000",
5718 => "0000000001011000",
5719 => "0000000001011000",
5720 => "0000000001011000",
5721 => "0000000001011000",
5722 => "0000000001011000",
5723 => "0000000001011000",
5724 => "0000000001011000",
5725 => "0000000001011000",
5726 => "0000000001011000",
5727 => "0000000001011000",
5728 => "0000000001011000",
5729 => "0000000001011000",
5730 => "0000000001011000",
5731 => "0000000001011000",
5732 => "0000000001011000",
5733 => "0000000001011001",
5734 => "0000000001011001",
5735 => "0000000001011001",
5736 => "0000000001011001",
5737 => "0000000001011001",
5738 => "0000000001011001",
5739 => "0000000001011001",
5740 => "0000000001011001",
5741 => "0000000001011001",
5742 => "0000000001011001",
5743 => "0000000001011001",
5744 => "0000000001011001",
5745 => "0000000001011001",
5746 => "0000000001011001",
5747 => "0000000001011001",
5748 => "0000000001011001",
5749 => "0000000001011001",
5750 => "0000000001011001",
5751 => "0000000001011001",
5752 => "0000000001011001",
5753 => "0000000001011001",
5754 => "0000000001011001",
5755 => "0000000001011001",
5756 => "0000000001011001",
5757 => "0000000001011001",
5758 => "0000000001011001",
5759 => "0000000001011001",
5760 => "0000000001011001",
5761 => "0000000001011001",
5762 => "0000000001011001",
5763 => "0000000001011001",
5764 => "0000000001011001",
5765 => "0000000001011001",
5766 => "0000000001011001",
5767 => "0000000001011001",
5768 => "0000000001011001",
5769 => "0000000001011001",
5770 => "0000000001011001",
5771 => "0000000001011001",
5772 => "0000000001011001",
5773 => "0000000001011001",
5774 => "0000000001011001",
5775 => "0000000001011001",
5776 => "0000000001011001",
5777 => "0000000001011001",
5778 => "0000000001011001",
5779 => "0000000001011010",
5780 => "0000000001011010",
5781 => "0000000001011010",
5782 => "0000000001011010",
5783 => "0000000001011010",
5784 => "0000000001011010",
5785 => "0000000001011010",
5786 => "0000000001011010",
5787 => "0000000001011010",
5788 => "0000000001011010",
5789 => "0000000001011010",
5790 => "0000000001011010",
5791 => "0000000001011010",
5792 => "0000000001011010",
5793 => "0000000001011010",
5794 => "0000000001011010",
5795 => "0000000001011010",
5796 => "0000000001011010",
5797 => "0000000001011010",
5798 => "0000000001011010",
5799 => "0000000001011010",
5800 => "0000000001011010",
5801 => "0000000001011010",
5802 => "0000000001011010",
5803 => "0000000001011010",
5804 => "0000000001011010",
5805 => "0000000001011010",
5806 => "0000000001011010",
5807 => "0000000001011010",
5808 => "0000000001011010",
5809 => "0000000001011010",
5810 => "0000000001011010",
5811 => "0000000001011010",
5812 => "0000000001011010",
5813 => "0000000001011010",
5814 => "0000000001011010",
5815 => "0000000001011010",
5816 => "0000000001011010",
5817 => "0000000001011010",
5818 => "0000000001011010",
5819 => "0000000001011010",
5820 => "0000000001011010",
5821 => "0000000001011010",
5822 => "0000000001011010",
5823 => "0000000001011010",
5824 => "0000000001011011",
5825 => "0000000001011011",
5826 => "0000000001011011",
5827 => "0000000001011011",
5828 => "0000000001011011",
5829 => "0000000001011011",
5830 => "0000000001011011",
5831 => "0000000001011011",
5832 => "0000000001011011",
5833 => "0000000001011011",
5834 => "0000000001011011",
5835 => "0000000001011011",
5836 => "0000000001011011",
5837 => "0000000001011011",
5838 => "0000000001011011",
5839 => "0000000001011011",
5840 => "0000000001011011",
5841 => "0000000001011011",
5842 => "0000000001011011",
5843 => "0000000001011011",
5844 => "0000000001011011",
5845 => "0000000001011011",
5846 => "0000000001011011",
5847 => "0000000001011011",
5848 => "0000000001011011",
5849 => "0000000001011011",
5850 => "0000000001011011",
5851 => "0000000001011011",
5852 => "0000000001011011",
5853 => "0000000001011011",
5854 => "0000000001011011",
5855 => "0000000001011011",
5856 => "0000000001011011",
5857 => "0000000001011011",
5858 => "0000000001011011",
5859 => "0000000001011011",
5860 => "0000000001011011",
5861 => "0000000001011011",
5862 => "0000000001011011",
5863 => "0000000001011011",
5864 => "0000000001011011",
5865 => "0000000001011011",
5866 => "0000000001011011",
5867 => "0000000001011011",
5868 => "0000000001011011",
5869 => "0000000001011100",
5870 => "0000000001011100",
5871 => "0000000001011100",
5872 => "0000000001011100",
5873 => "0000000001011100",
5874 => "0000000001011100",
5875 => "0000000001011100",
5876 => "0000000001011100",
5877 => "0000000001011100",
5878 => "0000000001011100",
5879 => "0000000001011100",
5880 => "0000000001011100",
5881 => "0000000001011100",
5882 => "0000000001011100",
5883 => "0000000001011100",
5884 => "0000000001011100",
5885 => "0000000001011100",
5886 => "0000000001011100",
5887 => "0000000001011100",
5888 => "0000000001011100",
5889 => "0000000001011100",
5890 => "0000000001011100",
5891 => "0000000001011100",
5892 => "0000000001011100",
5893 => "0000000001011100",
5894 => "0000000001011100",
5895 => "0000000001011100",
5896 => "0000000001011100",
5897 => "0000000001011100",
5898 => "0000000001011100",
5899 => "0000000001011100",
5900 => "0000000001011100",
5901 => "0000000001011100",
5902 => "0000000001011100",
5903 => "0000000001011100",
5904 => "0000000001011100",
5905 => "0000000001011100",
5906 => "0000000001011100",
5907 => "0000000001011100",
5908 => "0000000001011100",
5909 => "0000000001011100",
5910 => "0000000001011100",
5911 => "0000000001011100",
5912 => "0000000001011100",
5913 => "0000000001011100",
5914 => "0000000001011101",
5915 => "0000000001011101",
5916 => "0000000001011101",
5917 => "0000000001011101",
5918 => "0000000001011101",
5919 => "0000000001011101",
5920 => "0000000001011101",
5921 => "0000000001011101",
5922 => "0000000001011101",
5923 => "0000000001011101",
5924 => "0000000001011101",
5925 => "0000000001011101",
5926 => "0000000001011101",
5927 => "0000000001011101",
5928 => "0000000001011101",
5929 => "0000000001011101",
5930 => "0000000001011101",
5931 => "0000000001011101",
5932 => "0000000001011101",
5933 => "0000000001011101",
5934 => "0000000001011101",
5935 => "0000000001011101",
5936 => "0000000001011101",
5937 => "0000000001011101",
5938 => "0000000001011101",
5939 => "0000000001011101",
5940 => "0000000001011101",
5941 => "0000000001011101",
5942 => "0000000001011101",
5943 => "0000000001011101",
5944 => "0000000001011101",
5945 => "0000000001011101",
5946 => "0000000001011101",
5947 => "0000000001011101",
5948 => "0000000001011101",
5949 => "0000000001011101",
5950 => "0000000001011101",
5951 => "0000000001011101",
5952 => "0000000001011101",
5953 => "0000000001011101",
5954 => "0000000001011101",
5955 => "0000000001011101",
5956 => "0000000001011101",
5957 => "0000000001011101",
5958 => "0000000001011110",
5959 => "0000000001011110",
5960 => "0000000001011110",
5961 => "0000000001011110",
5962 => "0000000001011110",
5963 => "0000000001011110",
5964 => "0000000001011110",
5965 => "0000000001011110",
5966 => "0000000001011110",
5967 => "0000000001011110",
5968 => "0000000001011110",
5969 => "0000000001011110",
5970 => "0000000001011110",
5971 => "0000000001011110",
5972 => "0000000001011110",
5973 => "0000000001011110",
5974 => "0000000001011110",
5975 => "0000000001011110",
5976 => "0000000001011110",
5977 => "0000000001011110",
5978 => "0000000001011110",
5979 => "0000000001011110",
5980 => "0000000001011110",
5981 => "0000000001011110",
5982 => "0000000001011110",
5983 => "0000000001011110",
5984 => "0000000001011110",
5985 => "0000000001011110",
5986 => "0000000001011110",
5987 => "0000000001011110",
5988 => "0000000001011110",
5989 => "0000000001011110",
5990 => "0000000001011110",
5991 => "0000000001011110",
5992 => "0000000001011110",
5993 => "0000000001011110",
5994 => "0000000001011110",
5995 => "0000000001011110",
5996 => "0000000001011110",
5997 => "0000000001011110",
5998 => "0000000001011110",
5999 => "0000000001011110",
6000 => "0000000001011110",
6001 => "0000000001011111",
6002 => "0000000001011111",
6003 => "0000000001011111",
6004 => "0000000001011111",
6005 => "0000000001011111",
6006 => "0000000001011111",
6007 => "0000000001011111",
6008 => "0000000001011111",
6009 => "0000000001011111",
6010 => "0000000001011111",
6011 => "0000000001011111",
6012 => "0000000001011111",
6013 => "0000000001011111",
6014 => "0000000001011111",
6015 => "0000000001011111",
6016 => "0000000001011111",
6017 => "0000000001011111",
6018 => "0000000001011111",
6019 => "0000000001011111",
6020 => "0000000001011111",
6021 => "0000000001011111",
6022 => "0000000001011111",
6023 => "0000000001011111",
6024 => "0000000001011111",
6025 => "0000000001011111",
6026 => "0000000001011111",
6027 => "0000000001011111",
6028 => "0000000001011111",
6029 => "0000000001011111",
6030 => "0000000001011111",
6031 => "0000000001011111",
6032 => "0000000001011111",
6033 => "0000000001011111",
6034 => "0000000001011111",
6035 => "0000000001011111",
6036 => "0000000001011111",
6037 => "0000000001011111",
6038 => "0000000001011111",
6039 => "0000000001011111",
6040 => "0000000001011111",
6041 => "0000000001011111",
6042 => "0000000001011111",
6043 => "0000000001011111",
6044 => "0000000001100000",
6045 => "0000000001100000",
6046 => "0000000001100000",
6047 => "0000000001100000",
6048 => "0000000001100000",
6049 => "0000000001100000",
6050 => "0000000001100000",
6051 => "0000000001100000",
6052 => "0000000001100000",
6053 => "0000000001100000",
6054 => "0000000001100000",
6055 => "0000000001100000",
6056 => "0000000001100000",
6057 => "0000000001100000",
6058 => "0000000001100000",
6059 => "0000000001100000",
6060 => "0000000001100000",
6061 => "0000000001100000",
6062 => "0000000001100000",
6063 => "0000000001100000",
6064 => "0000000001100000",
6065 => "0000000001100000",
6066 => "0000000001100000",
6067 => "0000000001100000",
6068 => "0000000001100000",
6069 => "0000000001100000",
6070 => "0000000001100000",
6071 => "0000000001100000",
6072 => "0000000001100000",
6073 => "0000000001100000",
6074 => "0000000001100000",
6075 => "0000000001100000",
6076 => "0000000001100000",
6077 => "0000000001100000",
6078 => "0000000001100000",
6079 => "0000000001100000",
6080 => "0000000001100000",
6081 => "0000000001100000",
6082 => "0000000001100000",
6083 => "0000000001100000",
6084 => "0000000001100000",
6085 => "0000000001100000",
6086 => "0000000001100001",
6087 => "0000000001100001",
6088 => "0000000001100001",
6089 => "0000000001100001",
6090 => "0000000001100001",
6091 => "0000000001100001",
6092 => "0000000001100001",
6093 => "0000000001100001",
6094 => "0000000001100001",
6095 => "0000000001100001",
6096 => "0000000001100001",
6097 => "0000000001100001",
6098 => "0000000001100001",
6099 => "0000000001100001",
6100 => "0000000001100001",
6101 => "0000000001100001",
6102 => "0000000001100001",
6103 => "0000000001100001",
6104 => "0000000001100001",
6105 => "0000000001100001",
6106 => "0000000001100001",
6107 => "0000000001100001",
6108 => "0000000001100001",
6109 => "0000000001100001",
6110 => "0000000001100001",
6111 => "0000000001100001",
6112 => "0000000001100001",
6113 => "0000000001100001",
6114 => "0000000001100001",
6115 => "0000000001100001",
6116 => "0000000001100001",
6117 => "0000000001100001",
6118 => "0000000001100001",
6119 => "0000000001100001",
6120 => "0000000001100001",
6121 => "0000000001100001",
6122 => "0000000001100001",
6123 => "0000000001100001",
6124 => "0000000001100001",
6125 => "0000000001100001",
6126 => "0000000001100001",
6127 => "0000000001100001",
6128 => "0000000001100010",
6129 => "0000000001100010",
6130 => "0000000001100010",
6131 => "0000000001100010",
6132 => "0000000001100010",
6133 => "0000000001100010",
6134 => "0000000001100010",
6135 => "0000000001100010",
6136 => "0000000001100010",
6137 => "0000000001100010",
6138 => "0000000001100010",
6139 => "0000000001100010",
6140 => "0000000001100010",
6141 => "0000000001100010",
6142 => "0000000001100010",
6143 => "0000000001100010",
6144 => "0000000001100010",
6145 => "0000000001100010",
6146 => "0000000001100010",
6147 => "0000000001100010",
6148 => "0000000001100010",
6149 => "0000000001100010",
6150 => "0000000001100010",
6151 => "0000000001100010",
6152 => "0000000001100010",
6153 => "0000000001100010",
6154 => "0000000001100010",
6155 => "0000000001100010",
6156 => "0000000001100010",
6157 => "0000000001100010",
6158 => "0000000001100010",
6159 => "0000000001100010",
6160 => "0000000001100010",
6161 => "0000000001100010",
6162 => "0000000001100010",
6163 => "0000000001100010",
6164 => "0000000001100010",
6165 => "0000000001100010",
6166 => "0000000001100010",
6167 => "0000000001100010",
6168 => "0000000001100010",
6169 => "0000000001100010",
6170 => "0000000001100011",
6171 => "0000000001100011",
6172 => "0000000001100011",
6173 => "0000000001100011",
6174 => "0000000001100011",
6175 => "0000000001100011",
6176 => "0000000001100011",
6177 => "0000000001100011",
6178 => "0000000001100011",
6179 => "0000000001100011",
6180 => "0000000001100011",
6181 => "0000000001100011",
6182 => "0000000001100011",
6183 => "0000000001100011",
6184 => "0000000001100011",
6185 => "0000000001100011",
6186 => "0000000001100011",
6187 => "0000000001100011",
6188 => "0000000001100011",
6189 => "0000000001100011",
6190 => "0000000001100011",
6191 => "0000000001100011",
6192 => "0000000001100011",
6193 => "0000000001100011",
6194 => "0000000001100011",
6195 => "0000000001100011",
6196 => "0000000001100011",
6197 => "0000000001100011",
6198 => "0000000001100011",
6199 => "0000000001100011",
6200 => "0000000001100011",
6201 => "0000000001100011",
6202 => "0000000001100011",
6203 => "0000000001100011",
6204 => "0000000001100011",
6205 => "0000000001100011",
6206 => "0000000001100011",
6207 => "0000000001100011",
6208 => "0000000001100011",
6209 => "0000000001100011",
6210 => "0000000001100011",
6211 => "0000000001100100",
6212 => "0000000001100100",
6213 => "0000000001100100",
6214 => "0000000001100100",
6215 => "0000000001100100",
6216 => "0000000001100100",
6217 => "0000000001100100",
6218 => "0000000001100100",
6219 => "0000000001100100",
6220 => "0000000001100100",
6221 => "0000000001100100",
6222 => "0000000001100100",
6223 => "0000000001100100",
6224 => "0000000001100100",
6225 => "0000000001100100",
6226 => "0000000001100100",
6227 => "0000000001100100",
6228 => "0000000001100100",
6229 => "0000000001100100",
6230 => "0000000001100100",
6231 => "0000000001100100",
6232 => "0000000001100100",
6233 => "0000000001100100",
6234 => "0000000001100100",
6235 => "0000000001100100",
6236 => "0000000001100100",
6237 => "0000000001100100",
6238 => "0000000001100100",
6239 => "0000000001100100",
6240 => "0000000001100100",
6241 => "0000000001100100",
6242 => "0000000001100100",
6243 => "0000000001100100",
6244 => "0000000001100100",
6245 => "0000000001100100",
6246 => "0000000001100100",
6247 => "0000000001100100",
6248 => "0000000001100100",
6249 => "0000000001100100",
6250 => "0000000001100100",
6251 => "0000000001100100",
6252 => "0000000001100101",
6253 => "0000000001100101",
6254 => "0000000001100101",
6255 => "0000000001100101",
6256 => "0000000001100101",
6257 => "0000000001100101",
6258 => "0000000001100101",
6259 => "0000000001100101",
6260 => "0000000001100101",
6261 => "0000000001100101",
6262 => "0000000001100101",
6263 => "0000000001100101",
6264 => "0000000001100101",
6265 => "0000000001100101",
6266 => "0000000001100101",
6267 => "0000000001100101",
6268 => "0000000001100101",
6269 => "0000000001100101",
6270 => "0000000001100101",
6271 => "0000000001100101",
6272 => "0000000001100101",
6273 => "0000000001100101",
6274 => "0000000001100101",
6275 => "0000000001100101",
6276 => "0000000001100101",
6277 => "0000000001100101",
6278 => "0000000001100101",
6279 => "0000000001100101",
6280 => "0000000001100101",
6281 => "0000000001100101",
6282 => "0000000001100101",
6283 => "0000000001100101",
6284 => "0000000001100101",
6285 => "0000000001100101",
6286 => "0000000001100101",
6287 => "0000000001100101",
6288 => "0000000001100101",
6289 => "0000000001100101",
6290 => "0000000001100101",
6291 => "0000000001100101",
6292 => "0000000001100101",
6293 => "0000000001100110",
6294 => "0000000001100110",
6295 => "0000000001100110",
6296 => "0000000001100110",
6297 => "0000000001100110",
6298 => "0000000001100110",
6299 => "0000000001100110",
6300 => "0000000001100110",
6301 => "0000000001100110",
6302 => "0000000001100110",
6303 => "0000000001100110",
6304 => "0000000001100110",
6305 => "0000000001100110",
6306 => "0000000001100110",
6307 => "0000000001100110",
6308 => "0000000001100110",
6309 => "0000000001100110",
6310 => "0000000001100110",
6311 => "0000000001100110",
6312 => "0000000001100110",
6313 => "0000000001100110",
6314 => "0000000001100110",
6315 => "0000000001100110",
6316 => "0000000001100110",
6317 => "0000000001100110",
6318 => "0000000001100110",
6319 => "0000000001100110",
6320 => "0000000001100110",
6321 => "0000000001100110",
6322 => "0000000001100110",
6323 => "0000000001100110",
6324 => "0000000001100110",
6325 => "0000000001100110",
6326 => "0000000001100110",
6327 => "0000000001100110",
6328 => "0000000001100110",
6329 => "0000000001100110",
6330 => "0000000001100110",
6331 => "0000000001100110",
6332 => "0000000001100110",
6333 => "0000000001100111",
6334 => "0000000001100111",
6335 => "0000000001100111",
6336 => "0000000001100111",
6337 => "0000000001100111",
6338 => "0000000001100111",
6339 => "0000000001100111",
6340 => "0000000001100111",
6341 => "0000000001100111",
6342 => "0000000001100111",
6343 => "0000000001100111",
6344 => "0000000001100111",
6345 => "0000000001100111",
6346 => "0000000001100111",
6347 => "0000000001100111",
6348 => "0000000001100111",
6349 => "0000000001100111",
6350 => "0000000001100111",
6351 => "0000000001100111",
6352 => "0000000001100111",
6353 => "0000000001100111",
6354 => "0000000001100111",
6355 => "0000000001100111",
6356 => "0000000001100111",
6357 => "0000000001100111",
6358 => "0000000001100111",
6359 => "0000000001100111",
6360 => "0000000001100111",
6361 => "0000000001100111",
6362 => "0000000001100111",
6363 => "0000000001100111",
6364 => "0000000001100111",
6365 => "0000000001100111",
6366 => "0000000001100111",
6367 => "0000000001100111",
6368 => "0000000001100111",
6369 => "0000000001100111",
6370 => "0000000001100111",
6371 => "0000000001100111",
6372 => "0000000001101000",
6373 => "0000000001101000",
6374 => "0000000001101000",
6375 => "0000000001101000",
6376 => "0000000001101000",
6377 => "0000000001101000",
6378 => "0000000001101000",
6379 => "0000000001101000",
6380 => "0000000001101000",
6381 => "0000000001101000",
6382 => "0000000001101000",
6383 => "0000000001101000",
6384 => "0000000001101000",
6385 => "0000000001101000",
6386 => "0000000001101000",
6387 => "0000000001101000",
6388 => "0000000001101000",
6389 => "0000000001101000",
6390 => "0000000001101000",
6391 => "0000000001101000",
6392 => "0000000001101000",
6393 => "0000000001101000",
6394 => "0000000001101000",
6395 => "0000000001101000",
6396 => "0000000001101000",
6397 => "0000000001101000",
6398 => "0000000001101000",
6399 => "0000000001101000",
6400 => "0000000001101000",
6401 => "0000000001101000",
6402 => "0000000001101000",
6403 => "0000000001101000",
6404 => "0000000001101000",
6405 => "0000000001101000",
6406 => "0000000001101000",
6407 => "0000000001101000",
6408 => "0000000001101000",
6409 => "0000000001101000",
6410 => "0000000001101000",
6411 => "0000000001101001",
6412 => "0000000001101001",
6413 => "0000000001101001",
6414 => "0000000001101001",
6415 => "0000000001101001",
6416 => "0000000001101001",
6417 => "0000000001101001",
6418 => "0000000001101001",
6419 => "0000000001101001",
6420 => "0000000001101001",
6421 => "0000000001101001",
6422 => "0000000001101001",
6423 => "0000000001101001",
6424 => "0000000001101001",
6425 => "0000000001101001",
6426 => "0000000001101001",
6427 => "0000000001101001",
6428 => "0000000001101001",
6429 => "0000000001101001",
6430 => "0000000001101001",
6431 => "0000000001101001",
6432 => "0000000001101001",
6433 => "0000000001101001",
6434 => "0000000001101001",
6435 => "0000000001101001",
6436 => "0000000001101001",
6437 => "0000000001101001",
6438 => "0000000001101001",
6439 => "0000000001101001",
6440 => "0000000001101001",
6441 => "0000000001101001",
6442 => "0000000001101001",
6443 => "0000000001101001",
6444 => "0000000001101001",
6445 => "0000000001101001",
6446 => "0000000001101001",
6447 => "0000000001101001",
6448 => "0000000001101001",
6449 => "0000000001101001",
6450 => "0000000001101010",
6451 => "0000000001101010",
6452 => "0000000001101010",
6453 => "0000000001101010",
6454 => "0000000001101010",
6455 => "0000000001101010",
6456 => "0000000001101010",
6457 => "0000000001101010",
6458 => "0000000001101010",
6459 => "0000000001101010",
6460 => "0000000001101010",
6461 => "0000000001101010",
6462 => "0000000001101010",
6463 => "0000000001101010",
6464 => "0000000001101010",
6465 => "0000000001101010",
6466 => "0000000001101010",
6467 => "0000000001101010",
6468 => "0000000001101010",
6469 => "0000000001101010",
6470 => "0000000001101010",
6471 => "0000000001101010",
6472 => "0000000001101010",
6473 => "0000000001101010",
6474 => "0000000001101010",
6475 => "0000000001101010",
6476 => "0000000001101010",
6477 => "0000000001101010",
6478 => "0000000001101010",
6479 => "0000000001101010",
6480 => "0000000001101010",
6481 => "0000000001101010",
6482 => "0000000001101010",
6483 => "0000000001101010",
6484 => "0000000001101010",
6485 => "0000000001101010",
6486 => "0000000001101010",
6487 => "0000000001101010",
6488 => "0000000001101010",
6489 => "0000000001101011",
6490 => "0000000001101011",
6491 => "0000000001101011",
6492 => "0000000001101011",
6493 => "0000000001101011",
6494 => "0000000001101011",
6495 => "0000000001101011",
6496 => "0000000001101011",
6497 => "0000000001101011",
6498 => "0000000001101011",
6499 => "0000000001101011",
6500 => "0000000001101011",
6501 => "0000000001101011",
6502 => "0000000001101011",
6503 => "0000000001101011",
6504 => "0000000001101011",
6505 => "0000000001101011",
6506 => "0000000001101011",
6507 => "0000000001101011",
6508 => "0000000001101011",
6509 => "0000000001101011",
6510 => "0000000001101011",
6511 => "0000000001101011",
6512 => "0000000001101011",
6513 => "0000000001101011",
6514 => "0000000001101011",
6515 => "0000000001101011",
6516 => "0000000001101011",
6517 => "0000000001101011",
6518 => "0000000001101011",
6519 => "0000000001101011",
6520 => "0000000001101011",
6521 => "0000000001101011",
6522 => "0000000001101011",
6523 => "0000000001101011",
6524 => "0000000001101011",
6525 => "0000000001101011",
6526 => "0000000001101011",
6527 => "0000000001101100",
6528 => "0000000001101100",
6529 => "0000000001101100",
6530 => "0000000001101100",
6531 => "0000000001101100",
6532 => "0000000001101100",
6533 => "0000000001101100",
6534 => "0000000001101100",
6535 => "0000000001101100",
6536 => "0000000001101100",
6537 => "0000000001101100",
6538 => "0000000001101100",
6539 => "0000000001101100",
6540 => "0000000001101100",
6541 => "0000000001101100",
6542 => "0000000001101100",
6543 => "0000000001101100",
6544 => "0000000001101100",
6545 => "0000000001101100",
6546 => "0000000001101100",
6547 => "0000000001101100",
6548 => "0000000001101100",
6549 => "0000000001101100",
6550 => "0000000001101100",
6551 => "0000000001101100",
6552 => "0000000001101100",
6553 => "0000000001101100",
6554 => "0000000001101100",
6555 => "0000000001101100",
6556 => "0000000001101100",
6557 => "0000000001101100",
6558 => "0000000001101100",
6559 => "0000000001101100",
6560 => "0000000001101100",
6561 => "0000000001101100",
6562 => "0000000001101100",
6563 => "0000000001101100",
6564 => "0000000001101100",
6565 => "0000000001101101",
6566 => "0000000001101101",
6567 => "0000000001101101",
6568 => "0000000001101101",
6569 => "0000000001101101",
6570 => "0000000001101101",
6571 => "0000000001101101",
6572 => "0000000001101101",
6573 => "0000000001101101",
6574 => "0000000001101101",
6575 => "0000000001101101",
6576 => "0000000001101101",
6577 => "0000000001101101",
6578 => "0000000001101101",
6579 => "0000000001101101",
6580 => "0000000001101101",
6581 => "0000000001101101",
6582 => "0000000001101101",
6583 => "0000000001101101",
6584 => "0000000001101101",
6585 => "0000000001101101",
6586 => "0000000001101101",
6587 => "0000000001101101",
6588 => "0000000001101101",
6589 => "0000000001101101",
6590 => "0000000001101101",
6591 => "0000000001101101",
6592 => "0000000001101101",
6593 => "0000000001101101",
6594 => "0000000001101101",
6595 => "0000000001101101",
6596 => "0000000001101101",
6597 => "0000000001101101",
6598 => "0000000001101101",
6599 => "0000000001101101",
6600 => "0000000001101101",
6601 => "0000000001101101",
6602 => "0000000001101110",
6603 => "0000000001101110",
6604 => "0000000001101110",
6605 => "0000000001101110",
6606 => "0000000001101110",
6607 => "0000000001101110",
6608 => "0000000001101110",
6609 => "0000000001101110",
6610 => "0000000001101110",
6611 => "0000000001101110",
6612 => "0000000001101110",
6613 => "0000000001101110",
6614 => "0000000001101110",
6615 => "0000000001101110",
6616 => "0000000001101110",
6617 => "0000000001101110",
6618 => "0000000001101110",
6619 => "0000000001101110",
6620 => "0000000001101110",
6621 => "0000000001101110",
6622 => "0000000001101110",
6623 => "0000000001101110",
6624 => "0000000001101110",
6625 => "0000000001101110",
6626 => "0000000001101110",
6627 => "0000000001101110",
6628 => "0000000001101110",
6629 => "0000000001101110",
6630 => "0000000001101110",
6631 => "0000000001101110",
6632 => "0000000001101110",
6633 => "0000000001101110",
6634 => "0000000001101110",
6635 => "0000000001101110",
6636 => "0000000001101110",
6637 => "0000000001101110",
6638 => "0000000001101110",
6639 => "0000000001101111",
6640 => "0000000001101111",
6641 => "0000000001101111",
6642 => "0000000001101111",
6643 => "0000000001101111",
6644 => "0000000001101111",
6645 => "0000000001101111",
6646 => "0000000001101111",
6647 => "0000000001101111",
6648 => "0000000001101111",
6649 => "0000000001101111",
6650 => "0000000001101111",
6651 => "0000000001101111",
6652 => "0000000001101111",
6653 => "0000000001101111",
6654 => "0000000001101111",
6655 => "0000000001101111",
6656 => "0000000001101111",
6657 => "0000000001101111",
6658 => "0000000001101111",
6659 => "0000000001101111",
6660 => "0000000001101111",
6661 => "0000000001101111",
6662 => "0000000001101111",
6663 => "0000000001101111",
6664 => "0000000001101111",
6665 => "0000000001101111",
6666 => "0000000001101111",
6667 => "0000000001101111",
6668 => "0000000001101111",
6669 => "0000000001101111",
6670 => "0000000001101111",
6671 => "0000000001101111",
6672 => "0000000001101111",
6673 => "0000000001101111",
6674 => "0000000001101111",
6675 => "0000000001101111",
6676 => "0000000001110000",
6677 => "0000000001110000",
6678 => "0000000001110000",
6679 => "0000000001110000",
6680 => "0000000001110000",
6681 => "0000000001110000",
6682 => "0000000001110000",
6683 => "0000000001110000",
6684 => "0000000001110000",
6685 => "0000000001110000",
6686 => "0000000001110000",
6687 => "0000000001110000",
6688 => "0000000001110000",
6689 => "0000000001110000",
6690 => "0000000001110000",
6691 => "0000000001110000",
6692 => "0000000001110000",
6693 => "0000000001110000",
6694 => "0000000001110000",
6695 => "0000000001110000",
6696 => "0000000001110000",
6697 => "0000000001110000",
6698 => "0000000001110000",
6699 => "0000000001110000",
6700 => "0000000001110000",
6701 => "0000000001110000",
6702 => "0000000001110000",
6703 => "0000000001110000",
6704 => "0000000001110000",
6705 => "0000000001110000",
6706 => "0000000001110000",
6707 => "0000000001110000",
6708 => "0000000001110000",
6709 => "0000000001110000",
6710 => "0000000001110000",
6711 => "0000000001110000",
6712 => "0000000001110000",
6713 => "0000000001110001",
6714 => "0000000001110001",
6715 => "0000000001110001",
6716 => "0000000001110001",
6717 => "0000000001110001",
6718 => "0000000001110001",
6719 => "0000000001110001",
6720 => "0000000001110001",
6721 => "0000000001110001",
6722 => "0000000001110001",
6723 => "0000000001110001",
6724 => "0000000001110001",
6725 => "0000000001110001",
6726 => "0000000001110001",
6727 => "0000000001110001",
6728 => "0000000001110001",
6729 => "0000000001110001",
6730 => "0000000001110001",
6731 => "0000000001110001",
6732 => "0000000001110001",
6733 => "0000000001110001",
6734 => "0000000001110001",
6735 => "0000000001110001",
6736 => "0000000001110001",
6737 => "0000000001110001",
6738 => "0000000001110001",
6739 => "0000000001110001",
6740 => "0000000001110001",
6741 => "0000000001110001",
6742 => "0000000001110001",
6743 => "0000000001110001",
6744 => "0000000001110001",
6745 => "0000000001110001",
6746 => "0000000001110001",
6747 => "0000000001110001",
6748 => "0000000001110001",
6749 => "0000000001110010",
6750 => "0000000001110010",
6751 => "0000000001110010",
6752 => "0000000001110010",
6753 => "0000000001110010",
6754 => "0000000001110010",
6755 => "0000000001110010",
6756 => "0000000001110010",
6757 => "0000000001110010",
6758 => "0000000001110010",
6759 => "0000000001110010",
6760 => "0000000001110010",
6761 => "0000000001110010",
6762 => "0000000001110010",
6763 => "0000000001110010",
6764 => "0000000001110010",
6765 => "0000000001110010",
6766 => "0000000001110010",
6767 => "0000000001110010",
6768 => "0000000001110010",
6769 => "0000000001110010",
6770 => "0000000001110010",
6771 => "0000000001110010",
6772 => "0000000001110010",
6773 => "0000000001110010",
6774 => "0000000001110010",
6775 => "0000000001110010",
6776 => "0000000001110010",
6777 => "0000000001110010",
6778 => "0000000001110010",
6779 => "0000000001110010",
6780 => "0000000001110010",
6781 => "0000000001110010",
6782 => "0000000001110010",
6783 => "0000000001110010",
6784 => "0000000001110010",
6785 => "0000000001110011",
6786 => "0000000001110011",
6787 => "0000000001110011",
6788 => "0000000001110011",
6789 => "0000000001110011",
6790 => "0000000001110011",
6791 => "0000000001110011",
6792 => "0000000001110011",
6793 => "0000000001110011",
6794 => "0000000001110011",
6795 => "0000000001110011",
6796 => "0000000001110011",
6797 => "0000000001110011",
6798 => "0000000001110011",
6799 => "0000000001110011",
6800 => "0000000001110011",
6801 => "0000000001110011",
6802 => "0000000001110011",
6803 => "0000000001110011",
6804 => "0000000001110011",
6805 => "0000000001110011",
6806 => "0000000001110011",
6807 => "0000000001110011",
6808 => "0000000001110011",
6809 => "0000000001110011",
6810 => "0000000001110011",
6811 => "0000000001110011",
6812 => "0000000001110011",
6813 => "0000000001110011",
6814 => "0000000001110011",
6815 => "0000000001110011",
6816 => "0000000001110011",
6817 => "0000000001110011",
6818 => "0000000001110011",
6819 => "0000000001110011",
6820 => "0000000001110100",
6821 => "0000000001110100",
6822 => "0000000001110100",
6823 => "0000000001110100",
6824 => "0000000001110100",
6825 => "0000000001110100",
6826 => "0000000001110100",
6827 => "0000000001110100",
6828 => "0000000001110100",
6829 => "0000000001110100",
6830 => "0000000001110100",
6831 => "0000000001110100",
6832 => "0000000001110100",
6833 => "0000000001110100",
6834 => "0000000001110100",
6835 => "0000000001110100",
6836 => "0000000001110100",
6837 => "0000000001110100",
6838 => "0000000001110100",
6839 => "0000000001110100",
6840 => "0000000001110100",
6841 => "0000000001110100",
6842 => "0000000001110100",
6843 => "0000000001110100",
6844 => "0000000001110100",
6845 => "0000000001110100",
6846 => "0000000001110100",
6847 => "0000000001110100",
6848 => "0000000001110100",
6849 => "0000000001110100",
6850 => "0000000001110100",
6851 => "0000000001110100",
6852 => "0000000001110100",
6853 => "0000000001110100",
6854 => "0000000001110100",
6855 => "0000000001110101",
6856 => "0000000001110101",
6857 => "0000000001110101",
6858 => "0000000001110101",
6859 => "0000000001110101",
6860 => "0000000001110101",
6861 => "0000000001110101",
6862 => "0000000001110101",
6863 => "0000000001110101",
6864 => "0000000001110101",
6865 => "0000000001110101",
6866 => "0000000001110101",
6867 => "0000000001110101",
6868 => "0000000001110101",
6869 => "0000000001110101",
6870 => "0000000001110101",
6871 => "0000000001110101",
6872 => "0000000001110101",
6873 => "0000000001110101",
6874 => "0000000001110101",
6875 => "0000000001110101",
6876 => "0000000001110101",
6877 => "0000000001110101",
6878 => "0000000001110101",
6879 => "0000000001110101",
6880 => "0000000001110101",
6881 => "0000000001110101",
6882 => "0000000001110101",
6883 => "0000000001110101",
6884 => "0000000001110101",
6885 => "0000000001110101",
6886 => "0000000001110101",
6887 => "0000000001110101",
6888 => "0000000001110101",
6889 => "0000000001110101",
6890 => "0000000001110110",
6891 => "0000000001110110",
6892 => "0000000001110110",
6893 => "0000000001110110",
6894 => "0000000001110110",
6895 => "0000000001110110",
6896 => "0000000001110110",
6897 => "0000000001110110",
6898 => "0000000001110110",
6899 => "0000000001110110",
6900 => "0000000001110110",
6901 => "0000000001110110",
6902 => "0000000001110110",
6903 => "0000000001110110",
6904 => "0000000001110110",
6905 => "0000000001110110",
6906 => "0000000001110110",
6907 => "0000000001110110",
6908 => "0000000001110110",
6909 => "0000000001110110",
6910 => "0000000001110110",
6911 => "0000000001110110",
6912 => "0000000001110110",
6913 => "0000000001110110",
6914 => "0000000001110110",
6915 => "0000000001110110",
6916 => "0000000001110110",
6917 => "0000000001110110",
6918 => "0000000001110110",
6919 => "0000000001110110",
6920 => "0000000001110110",
6921 => "0000000001110110",
6922 => "0000000001110110",
6923 => "0000000001110110",
6924 => "0000000001110110",
6925 => "0000000001110111",
6926 => "0000000001110111",
6927 => "0000000001110111",
6928 => "0000000001110111",
6929 => "0000000001110111",
6930 => "0000000001110111",
6931 => "0000000001110111",
6932 => "0000000001110111",
6933 => "0000000001110111",
6934 => "0000000001110111",
6935 => "0000000001110111",
6936 => "0000000001110111",
6937 => "0000000001110111",
6938 => "0000000001110111",
6939 => "0000000001110111",
6940 => "0000000001110111",
6941 => "0000000001110111",
6942 => "0000000001110111",
6943 => "0000000001110111",
6944 => "0000000001110111",
6945 => "0000000001110111",
6946 => "0000000001110111",
6947 => "0000000001110111",
6948 => "0000000001110111",
6949 => "0000000001110111",
6950 => "0000000001110111",
6951 => "0000000001110111",
6952 => "0000000001110111",
6953 => "0000000001110111",
6954 => "0000000001110111",
6955 => "0000000001110111",
6956 => "0000000001110111",
6957 => "0000000001110111",
6958 => "0000000001110111",
6959 => "0000000001111000",
6960 => "0000000001111000",
6961 => "0000000001111000",
6962 => "0000000001111000",
6963 => "0000000001111000",
6964 => "0000000001111000",
6965 => "0000000001111000",
6966 => "0000000001111000",
6967 => "0000000001111000",
6968 => "0000000001111000",
6969 => "0000000001111000",
6970 => "0000000001111000",
6971 => "0000000001111000",
6972 => "0000000001111000",
6973 => "0000000001111000",
6974 => "0000000001111000",
6975 => "0000000001111000",
6976 => "0000000001111000",
6977 => "0000000001111000",
6978 => "0000000001111000",
6979 => "0000000001111000",
6980 => "0000000001111000",
6981 => "0000000001111000",
6982 => "0000000001111000",
6983 => "0000000001111000",
6984 => "0000000001111000",
6985 => "0000000001111000",
6986 => "0000000001111000",
6987 => "0000000001111000",
6988 => "0000000001111000",
6989 => "0000000001111000",
6990 => "0000000001111000",
6991 => "0000000001111000",
6992 => "0000000001111000",
6993 => "0000000001111001",
6994 => "0000000001111001",
6995 => "0000000001111001",
6996 => "0000000001111001",
6997 => "0000000001111001",
6998 => "0000000001111001",
6999 => "0000000001111001",
7000 => "0000000001111001",
7001 => "0000000001111001",
7002 => "0000000001111001",
7003 => "0000000001111001",
7004 => "0000000001111001",
7005 => "0000000001111001",
7006 => "0000000001111001",
7007 => "0000000001111001",
7008 => "0000000001111001",
7009 => "0000000001111001",
7010 => "0000000001111001",
7011 => "0000000001111001",
7012 => "0000000001111001",
7013 => "0000000001111001",
7014 => "0000000001111001",
7015 => "0000000001111001",
7016 => "0000000001111001",
7017 => "0000000001111001",
7018 => "0000000001111001",
7019 => "0000000001111001",
7020 => "0000000001111001",
7021 => "0000000001111001",
7022 => "0000000001111001",
7023 => "0000000001111001",
7024 => "0000000001111001",
7025 => "0000000001111001",
7026 => "0000000001111001",
7027 => "0000000001111010",
7028 => "0000000001111010",
7029 => "0000000001111010",
7030 => "0000000001111010",
7031 => "0000000001111010",
7032 => "0000000001111010",
7033 => "0000000001111010",
7034 => "0000000001111010",
7035 => "0000000001111010",
7036 => "0000000001111010",
7037 => "0000000001111010",
7038 => "0000000001111010",
7039 => "0000000001111010",
7040 => "0000000001111010",
7041 => "0000000001111010",
7042 => "0000000001111010",
7043 => "0000000001111010",
7044 => "0000000001111010",
7045 => "0000000001111010",
7046 => "0000000001111010",
7047 => "0000000001111010",
7048 => "0000000001111010",
7049 => "0000000001111010",
7050 => "0000000001111010",
7051 => "0000000001111010",
7052 => "0000000001111010",
7053 => "0000000001111010",
7054 => "0000000001111010",
7055 => "0000000001111010",
7056 => "0000000001111010",
7057 => "0000000001111010",
7058 => "0000000001111010",
7059 => "0000000001111010",
7060 => "0000000001111010",
7061 => "0000000001111011",
7062 => "0000000001111011",
7063 => "0000000001111011",
7064 => "0000000001111011",
7065 => "0000000001111011",
7066 => "0000000001111011",
7067 => "0000000001111011",
7068 => "0000000001111011",
7069 => "0000000001111011",
7070 => "0000000001111011",
7071 => "0000000001111011",
7072 => "0000000001111011",
7073 => "0000000001111011",
7074 => "0000000001111011",
7075 => "0000000001111011",
7076 => "0000000001111011",
7077 => "0000000001111011",
7078 => "0000000001111011",
7079 => "0000000001111011",
7080 => "0000000001111011",
7081 => "0000000001111011",
7082 => "0000000001111011",
7083 => "0000000001111011",
7084 => "0000000001111011",
7085 => "0000000001111011",
7086 => "0000000001111011",
7087 => "0000000001111011",
7088 => "0000000001111011",
7089 => "0000000001111011",
7090 => "0000000001111011",
7091 => "0000000001111011",
7092 => "0000000001111011",
7093 => "0000000001111011",
7094 => "0000000001111100",
7095 => "0000000001111100",
7096 => "0000000001111100",
7097 => "0000000001111100",
7098 => "0000000001111100",
7099 => "0000000001111100",
7100 => "0000000001111100",
7101 => "0000000001111100",
7102 => "0000000001111100",
7103 => "0000000001111100",
7104 => "0000000001111100",
7105 => "0000000001111100",
7106 => "0000000001111100",
7107 => "0000000001111100",
7108 => "0000000001111100",
7109 => "0000000001111100",
7110 => "0000000001111100",
7111 => "0000000001111100",
7112 => "0000000001111100",
7113 => "0000000001111100",
7114 => "0000000001111100",
7115 => "0000000001111100",
7116 => "0000000001111100",
7117 => "0000000001111100",
7118 => "0000000001111100",
7119 => "0000000001111100",
7120 => "0000000001111100",
7121 => "0000000001111100",
7122 => "0000000001111100",
7123 => "0000000001111100",
7124 => "0000000001111100",
7125 => "0000000001111100",
7126 => "0000000001111100",
7127 => "0000000001111101",
7128 => "0000000001111101",
7129 => "0000000001111101",
7130 => "0000000001111101",
7131 => "0000000001111101",
7132 => "0000000001111101",
7133 => "0000000001111101",
7134 => "0000000001111101",
7135 => "0000000001111101",
7136 => "0000000001111101",
7137 => "0000000001111101",
7138 => "0000000001111101",
7139 => "0000000001111101",
7140 => "0000000001111101",
7141 => "0000000001111101",
7142 => "0000000001111101",
7143 => "0000000001111101",
7144 => "0000000001111101",
7145 => "0000000001111101",
7146 => "0000000001111101",
7147 => "0000000001111101",
7148 => "0000000001111101",
7149 => "0000000001111101",
7150 => "0000000001111101",
7151 => "0000000001111101",
7152 => "0000000001111101",
7153 => "0000000001111101",
7154 => "0000000001111101",
7155 => "0000000001111101",
7156 => "0000000001111101",
7157 => "0000000001111101",
7158 => "0000000001111101",
7159 => "0000000001111101",
7160 => "0000000001111110",
7161 => "0000000001111110",
7162 => "0000000001111110",
7163 => "0000000001111110",
7164 => "0000000001111110",
7165 => "0000000001111110",
7166 => "0000000001111110",
7167 => "0000000001111110",
7168 => "0000000001111110",
7169 => "0000000001111110",
7170 => "0000000001111110",
7171 => "0000000001111110",
7172 => "0000000001111110",
7173 => "0000000001111110",
7174 => "0000000001111110",
7175 => "0000000001111110",
7176 => "0000000001111110",
7177 => "0000000001111110",
7178 => "0000000001111110",
7179 => "0000000001111110",
7180 => "0000000001111110",
7181 => "0000000001111110",
7182 => "0000000001111110",
7183 => "0000000001111110",
7184 => "0000000001111110",
7185 => "0000000001111110",
7186 => "0000000001111110",
7187 => "0000000001111110",
7188 => "0000000001111110",
7189 => "0000000001111110",
7190 => "0000000001111110",
7191 => "0000000001111110",
7192 => "0000000001111111",
7193 => "0000000001111111",
7194 => "0000000001111111",
7195 => "0000000001111111",
7196 => "0000000001111111",
7197 => "0000000001111111",
7198 => "0000000001111111",
7199 => "0000000001111111",
7200 => "0000000001111111",
7201 => "0000000001111111",
7202 => "0000000001111111",
7203 => "0000000001111111",
7204 => "0000000001111111",
7205 => "0000000001111111",
7206 => "0000000001111111",
7207 => "0000000001111111",
7208 => "0000000001111111",
7209 => "0000000001111111",
7210 => "0000000001111111",
7211 => "0000000001111111",
7212 => "0000000001111111",
7213 => "0000000001111111",
7214 => "0000000001111111",
7215 => "0000000001111111",
7216 => "0000000001111111",
7217 => "0000000001111111",
7218 => "0000000001111111",
7219 => "0000000001111111",
7220 => "0000000001111111",
7221 => "0000000001111111",
7222 => "0000000001111111",
7223 => "0000000001111111",
7224 => "0000000010000000",
7225 => "0000000010000000",
7226 => "0000000010000000",
7227 => "0000000010000000",
7228 => "0000000010000000",
7229 => "0000000010000000",
7230 => "0000000010000000",
7231 => "0000000010000000",
7232 => "0000000010000000",
7233 => "0000000010000000",
7234 => "0000000010000000",
7235 => "0000000010000000",
7236 => "0000000010000000",
7237 => "0000000010000000",
7238 => "0000000010000000",
7239 => "0000000010000000",
7240 => "0000000010000000",
7241 => "0000000010000000",
7242 => "0000000010000000",
7243 => "0000000010000000",
7244 => "0000000010000000",
7245 => "0000000010000000",
7246 => "0000000010000000",
7247 => "0000000010000000",
7248 => "0000000010000000",
7249 => "0000000010000000",
7250 => "0000000010000000",
7251 => "0000000010000000",
7252 => "0000000010000000",
7253 => "0000000010000000",
7254 => "0000000010000000",
7255 => "0000000010000000",
7256 => "0000000010000001",
7257 => "0000000010000001",
7258 => "0000000010000001",
7259 => "0000000010000001",
7260 => "0000000010000001",
7261 => "0000000010000001",
7262 => "0000000010000001",
7263 => "0000000010000001",
7264 => "0000000010000001",
7265 => "0000000010000001",
7266 => "0000000010000001",
7267 => "0000000010000001",
7268 => "0000000010000001",
7269 => "0000000010000001",
7270 => "0000000010000001",
7271 => "0000000010000001",
7272 => "0000000010000001",
7273 => "0000000010000001",
7274 => "0000000010000001",
7275 => "0000000010000001",
7276 => "0000000010000001",
7277 => "0000000010000001",
7278 => "0000000010000001",
7279 => "0000000010000001",
7280 => "0000000010000001",
7281 => "0000000010000001",
7282 => "0000000010000001",
7283 => "0000000010000001",
7284 => "0000000010000001",
7285 => "0000000010000001",
7286 => "0000000010000001",
7287 => "0000000010000001",
7288 => "0000000010000010",
7289 => "0000000010000010",
7290 => "0000000010000010",
7291 => "0000000010000010",
7292 => "0000000010000010",
7293 => "0000000010000010",
7294 => "0000000010000010",
7295 => "0000000010000010",
7296 => "0000000010000010",
7297 => "0000000010000010",
7298 => "0000000010000010",
7299 => "0000000010000010",
7300 => "0000000010000010",
7301 => "0000000010000010",
7302 => "0000000010000010",
7303 => "0000000010000010",
7304 => "0000000010000010",
7305 => "0000000010000010",
7306 => "0000000010000010",
7307 => "0000000010000010",
7308 => "0000000010000010",
7309 => "0000000010000010",
7310 => "0000000010000010",
7311 => "0000000010000010",
7312 => "0000000010000010",
7313 => "0000000010000010",
7314 => "0000000010000010",
7315 => "0000000010000010",
7316 => "0000000010000010",
7317 => "0000000010000010",
7318 => "0000000010000010",
7319 => "0000000010000011",
7320 => "0000000010000011",
7321 => "0000000010000011",
7322 => "0000000010000011",
7323 => "0000000010000011",
7324 => "0000000010000011",
7325 => "0000000010000011",
7326 => "0000000010000011",
7327 => "0000000010000011",
7328 => "0000000010000011",
7329 => "0000000010000011",
7330 => "0000000010000011",
7331 => "0000000010000011",
7332 => "0000000010000011",
7333 => "0000000010000011",
7334 => "0000000010000011",
7335 => "0000000010000011",
7336 => "0000000010000011",
7337 => "0000000010000011",
7338 => "0000000010000011",
7339 => "0000000010000011",
7340 => "0000000010000011",
7341 => "0000000010000011",
7342 => "0000000010000011",
7343 => "0000000010000011",
7344 => "0000000010000011",
7345 => "0000000010000011",
7346 => "0000000010000011",
7347 => "0000000010000011",
7348 => "0000000010000011",
7349 => "0000000010000011",
7350 => "0000000010000011",
7351 => "0000000010000100",
7352 => "0000000010000100",
7353 => "0000000010000100",
7354 => "0000000010000100",
7355 => "0000000010000100",
7356 => "0000000010000100",
7357 => "0000000010000100",
7358 => "0000000010000100",
7359 => "0000000010000100",
7360 => "0000000010000100",
7361 => "0000000010000100",
7362 => "0000000010000100",
7363 => "0000000010000100",
7364 => "0000000010000100",
7365 => "0000000010000100",
7366 => "0000000010000100",
7367 => "0000000010000100",
7368 => "0000000010000100",
7369 => "0000000010000100",
7370 => "0000000010000100",
7371 => "0000000010000100",
7372 => "0000000010000100",
7373 => "0000000010000100",
7374 => "0000000010000100",
7375 => "0000000010000100",
7376 => "0000000010000100",
7377 => "0000000010000100",
7378 => "0000000010000100",
7379 => "0000000010000100",
7380 => "0000000010000100",
7381 => "0000000010000101",
7382 => "0000000010000101",
7383 => "0000000010000101",
7384 => "0000000010000101",
7385 => "0000000010000101",
7386 => "0000000010000101",
7387 => "0000000010000101",
7388 => "0000000010000101",
7389 => "0000000010000101",
7390 => "0000000010000101",
7391 => "0000000010000101",
7392 => "0000000010000101",
7393 => "0000000010000101",
7394 => "0000000010000101",
7395 => "0000000010000101",
7396 => "0000000010000101",
7397 => "0000000010000101",
7398 => "0000000010000101",
7399 => "0000000010000101",
7400 => "0000000010000101",
7401 => "0000000010000101",
7402 => "0000000010000101",
7403 => "0000000010000101",
7404 => "0000000010000101",
7405 => "0000000010000101",
7406 => "0000000010000101",
7407 => "0000000010000101",
7408 => "0000000010000101",
7409 => "0000000010000101",
7410 => "0000000010000101",
7411 => "0000000010000101",
7412 => "0000000010000110",
7413 => "0000000010000110",
7414 => "0000000010000110",
7415 => "0000000010000110",
7416 => "0000000010000110",
7417 => "0000000010000110",
7418 => "0000000010000110",
7419 => "0000000010000110",
7420 => "0000000010000110",
7421 => "0000000010000110",
7422 => "0000000010000110",
7423 => "0000000010000110",
7424 => "0000000010000110",
7425 => "0000000010000110",
7426 => "0000000010000110",
7427 => "0000000010000110",
7428 => "0000000010000110",
7429 => "0000000010000110",
7430 => "0000000010000110",
7431 => "0000000010000110",
7432 => "0000000010000110",
7433 => "0000000010000110",
7434 => "0000000010000110",
7435 => "0000000010000110",
7436 => "0000000010000110",
7437 => "0000000010000110",
7438 => "0000000010000110",
7439 => "0000000010000110",
7440 => "0000000010000110",
7441 => "0000000010000110",
7442 => "0000000010000110",
7443 => "0000000010000111",
7444 => "0000000010000111",
7445 => "0000000010000111",
7446 => "0000000010000111",
7447 => "0000000010000111",
7448 => "0000000010000111",
7449 => "0000000010000111",
7450 => "0000000010000111",
7451 => "0000000010000111",
7452 => "0000000010000111",
7453 => "0000000010000111",
7454 => "0000000010000111",
7455 => "0000000010000111",
7456 => "0000000010000111",
7457 => "0000000010000111",
7458 => "0000000010000111",
7459 => "0000000010000111",
7460 => "0000000010000111",
7461 => "0000000010000111",
7462 => "0000000010000111",
7463 => "0000000010000111",
7464 => "0000000010000111",
7465 => "0000000010000111",
7466 => "0000000010000111",
7467 => "0000000010000111",
7468 => "0000000010000111",
7469 => "0000000010000111",
7470 => "0000000010000111",
7471 => "0000000010000111",
7472 => "0000000010000111",
7473 => "0000000010001000",
7474 => "0000000010001000",
7475 => "0000000010001000",
7476 => "0000000010001000",
7477 => "0000000010001000",
7478 => "0000000010001000",
7479 => "0000000010001000",
7480 => "0000000010001000",
7481 => "0000000010001000",
7482 => "0000000010001000",
7483 => "0000000010001000",
7484 => "0000000010001000",
7485 => "0000000010001000",
7486 => "0000000010001000",
7487 => "0000000010001000",
7488 => "0000000010001000",
7489 => "0000000010001000",
7490 => "0000000010001000",
7491 => "0000000010001000",
7492 => "0000000010001000",
7493 => "0000000010001000",
7494 => "0000000010001000",
7495 => "0000000010001000",
7496 => "0000000010001000",
7497 => "0000000010001000",
7498 => "0000000010001000",
7499 => "0000000010001000",
7500 => "0000000010001000",
7501 => "0000000010001000",
7502 => "0000000010001000",
7503 => "0000000010001001",
7504 => "0000000010001001",
7505 => "0000000010001001",
7506 => "0000000010001001",
7507 => "0000000010001001",
7508 => "0000000010001001",
7509 => "0000000010001001",
7510 => "0000000010001001",
7511 => "0000000010001001",
7512 => "0000000010001001",
7513 => "0000000010001001",
7514 => "0000000010001001",
7515 => "0000000010001001",
7516 => "0000000010001001",
7517 => "0000000010001001",
7518 => "0000000010001001",
7519 => "0000000010001001",
7520 => "0000000010001001",
7521 => "0000000010001001",
7522 => "0000000010001001",
7523 => "0000000010001001",
7524 => "0000000010001001",
7525 => "0000000010001001",
7526 => "0000000010001001",
7527 => "0000000010001001",
7528 => "0000000010001001",
7529 => "0000000010001001",
7530 => "0000000010001001",
7531 => "0000000010001001",
7532 => "0000000010001001",
7533 => "0000000010001010",
7534 => "0000000010001010",
7535 => "0000000010001010",
7536 => "0000000010001010",
7537 => "0000000010001010",
7538 => "0000000010001010",
7539 => "0000000010001010",
7540 => "0000000010001010",
7541 => "0000000010001010",
7542 => "0000000010001010",
7543 => "0000000010001010",
7544 => "0000000010001010",
7545 => "0000000010001010",
7546 => "0000000010001010",
7547 => "0000000010001010",
7548 => "0000000010001010",
7549 => "0000000010001010",
7550 => "0000000010001010",
7551 => "0000000010001010",
7552 => "0000000010001010",
7553 => "0000000010001010",
7554 => "0000000010001010",
7555 => "0000000010001010",
7556 => "0000000010001010",
7557 => "0000000010001010",
7558 => "0000000010001010",
7559 => "0000000010001010",
7560 => "0000000010001010",
7561 => "0000000010001010",
7562 => "0000000010001010",
7563 => "0000000010001011",
7564 => "0000000010001011",
7565 => "0000000010001011",
7566 => "0000000010001011",
7567 => "0000000010001011",
7568 => "0000000010001011",
7569 => "0000000010001011",
7570 => "0000000010001011",
7571 => "0000000010001011",
7572 => "0000000010001011",
7573 => "0000000010001011",
7574 => "0000000010001011",
7575 => "0000000010001011",
7576 => "0000000010001011",
7577 => "0000000010001011",
7578 => "0000000010001011",
7579 => "0000000010001011",
7580 => "0000000010001011",
7581 => "0000000010001011",
7582 => "0000000010001011",
7583 => "0000000010001011",
7584 => "0000000010001011",
7585 => "0000000010001011",
7586 => "0000000010001011",
7587 => "0000000010001011",
7588 => "0000000010001011",
7589 => "0000000010001011",
7590 => "0000000010001011",
7591 => "0000000010001011",
7592 => "0000000010001100",
7593 => "0000000010001100",
7594 => "0000000010001100",
7595 => "0000000010001100",
7596 => "0000000010001100",
7597 => "0000000010001100",
7598 => "0000000010001100",
7599 => "0000000010001100",
7600 => "0000000010001100",
7601 => "0000000010001100",
7602 => "0000000010001100",
7603 => "0000000010001100",
7604 => "0000000010001100",
7605 => "0000000010001100",
7606 => "0000000010001100",
7607 => "0000000010001100",
7608 => "0000000010001100",
7609 => "0000000010001100",
7610 => "0000000010001100",
7611 => "0000000010001100",
7612 => "0000000010001100",
7613 => "0000000010001100",
7614 => "0000000010001100",
7615 => "0000000010001100",
7616 => "0000000010001100",
7617 => "0000000010001100",
7618 => "0000000010001100",
7619 => "0000000010001100",
7620 => "0000000010001100",
7621 => "0000000010001101",
7622 => "0000000010001101",
7623 => "0000000010001101",
7624 => "0000000010001101",
7625 => "0000000010001101",
7626 => "0000000010001101",
7627 => "0000000010001101",
7628 => "0000000010001101",
7629 => "0000000010001101",
7630 => "0000000010001101",
7631 => "0000000010001101",
7632 => "0000000010001101",
7633 => "0000000010001101",
7634 => "0000000010001101",
7635 => "0000000010001101",
7636 => "0000000010001101",
7637 => "0000000010001101",
7638 => "0000000010001101",
7639 => "0000000010001101",
7640 => "0000000010001101",
7641 => "0000000010001101",
7642 => "0000000010001101",
7643 => "0000000010001101",
7644 => "0000000010001101",
7645 => "0000000010001101",
7646 => "0000000010001101",
7647 => "0000000010001101",
7648 => "0000000010001101",
7649 => "0000000010001101",
7650 => "0000000010001110",
7651 => "0000000010001110",
7652 => "0000000010001110",
7653 => "0000000010001110",
7654 => "0000000010001110",
7655 => "0000000010001110",
7656 => "0000000010001110",
7657 => "0000000010001110",
7658 => "0000000010001110",
7659 => "0000000010001110",
7660 => "0000000010001110",
7661 => "0000000010001110",
7662 => "0000000010001110",
7663 => "0000000010001110",
7664 => "0000000010001110",
7665 => "0000000010001110",
7666 => "0000000010001110",
7667 => "0000000010001110",
7668 => "0000000010001110",
7669 => "0000000010001110",
7670 => "0000000010001110",
7671 => "0000000010001110",
7672 => "0000000010001110",
7673 => "0000000010001110",
7674 => "0000000010001110",
7675 => "0000000010001110",
7676 => "0000000010001110",
7677 => "0000000010001110",
7678 => "0000000010001110",
7679 => "0000000010001111",
7680 => "0000000010001111",
7681 => "0000000010001111",
7682 => "0000000010001111",
7683 => "0000000010001111",
7684 => "0000000010001111",
7685 => "0000000010001111",
7686 => "0000000010001111",
7687 => "0000000010001111",
7688 => "0000000010001111",
7689 => "0000000010001111",
7690 => "0000000010001111",
7691 => "0000000010001111",
7692 => "0000000010001111",
7693 => "0000000010001111",
7694 => "0000000010001111",
7695 => "0000000010001111",
7696 => "0000000010001111",
7697 => "0000000010001111",
7698 => "0000000010001111",
7699 => "0000000010001111",
7700 => "0000000010001111",
7701 => "0000000010001111",
7702 => "0000000010001111",
7703 => "0000000010001111",
7704 => "0000000010001111",
7705 => "0000000010001111",
7706 => "0000000010001111",
7707 => "0000000010001111",
7708 => "0000000010010000",
7709 => "0000000010010000",
7710 => "0000000010010000",
7711 => "0000000010010000",
7712 => "0000000010010000",
7713 => "0000000010010000",
7714 => "0000000010010000",
7715 => "0000000010010000",
7716 => "0000000010010000",
7717 => "0000000010010000",
7718 => "0000000010010000",
7719 => "0000000010010000",
7720 => "0000000010010000",
7721 => "0000000010010000",
7722 => "0000000010010000",
7723 => "0000000010010000",
7724 => "0000000010010000",
7725 => "0000000010010000",
7726 => "0000000010010000",
7727 => "0000000010010000",
7728 => "0000000010010000",
7729 => "0000000010010000",
7730 => "0000000010010000",
7731 => "0000000010010000",
7732 => "0000000010010000",
7733 => "0000000010010000",
7734 => "0000000010010000",
7735 => "0000000010010000",
7736 => "0000000010010001",
7737 => "0000000010010001",
7738 => "0000000010010001",
7739 => "0000000010010001",
7740 => "0000000010010001",
7741 => "0000000010010001",
7742 => "0000000010010001",
7743 => "0000000010010001",
7744 => "0000000010010001",
7745 => "0000000010010001",
7746 => "0000000010010001",
7747 => "0000000010010001",
7748 => "0000000010010001",
7749 => "0000000010010001",
7750 => "0000000010010001",
7751 => "0000000010010001",
7752 => "0000000010010001",
7753 => "0000000010010001",
7754 => "0000000010010001",
7755 => "0000000010010001",
7756 => "0000000010010001",
7757 => "0000000010010001",
7758 => "0000000010010001",
7759 => "0000000010010001",
7760 => "0000000010010001",
7761 => "0000000010010001",
7762 => "0000000010010001",
7763 => "0000000010010001",
7764 => "0000000010010010",
7765 => "0000000010010010",
7766 => "0000000010010010",
7767 => "0000000010010010",
7768 => "0000000010010010",
7769 => "0000000010010010",
7770 => "0000000010010010",
7771 => "0000000010010010",
7772 => "0000000010010010",
7773 => "0000000010010010",
7774 => "0000000010010010",
7775 => "0000000010010010",
7776 => "0000000010010010",
7777 => "0000000010010010",
7778 => "0000000010010010",
7779 => "0000000010010010",
7780 => "0000000010010010",
7781 => "0000000010010010",
7782 => "0000000010010010",
7783 => "0000000010010010",
7784 => "0000000010010010",
7785 => "0000000010010010",
7786 => "0000000010010010",
7787 => "0000000010010010",
7788 => "0000000010010010",
7789 => "0000000010010010",
7790 => "0000000010010010",
7791 => "0000000010010010",
7792 => "0000000010010011",
7793 => "0000000010010011",
7794 => "0000000010010011",
7795 => "0000000010010011",
7796 => "0000000010010011",
7797 => "0000000010010011",
7798 => "0000000010010011",
7799 => "0000000010010011",
7800 => "0000000010010011",
7801 => "0000000010010011",
7802 => "0000000010010011",
7803 => "0000000010010011",
7804 => "0000000010010011",
7805 => "0000000010010011",
7806 => "0000000010010011",
7807 => "0000000010010011",
7808 => "0000000010010011",
7809 => "0000000010010011",
7810 => "0000000010010011",
7811 => "0000000010010011",
7812 => "0000000010010011",
7813 => "0000000010010011",
7814 => "0000000010010011",
7815 => "0000000010010011",
7816 => "0000000010010011",
7817 => "0000000010010011",
7818 => "0000000010010011",
7819 => "0000000010010011",
7820 => "0000000010010100",
7821 => "0000000010010100",
7822 => "0000000010010100",
7823 => "0000000010010100",
7824 => "0000000010010100",
7825 => "0000000010010100",
7826 => "0000000010010100",
7827 => "0000000010010100",
7828 => "0000000010010100",
7829 => "0000000010010100",
7830 => "0000000010010100",
7831 => "0000000010010100",
7832 => "0000000010010100",
7833 => "0000000010010100",
7834 => "0000000010010100",
7835 => "0000000010010100",
7836 => "0000000010010100",
7837 => "0000000010010100",
7838 => "0000000010010100",
7839 => "0000000010010100",
7840 => "0000000010010100",
7841 => "0000000010010100",
7842 => "0000000010010100",
7843 => "0000000010010100",
7844 => "0000000010010100",
7845 => "0000000010010100",
7846 => "0000000010010100",
7847 => "0000000010010100",
7848 => "0000000010010101",
7849 => "0000000010010101",
7850 => "0000000010010101",
7851 => "0000000010010101",
7852 => "0000000010010101",
7853 => "0000000010010101",
7854 => "0000000010010101",
7855 => "0000000010010101",
7856 => "0000000010010101",
7857 => "0000000010010101",
7858 => "0000000010010101",
7859 => "0000000010010101",
7860 => "0000000010010101",
7861 => "0000000010010101",
7862 => "0000000010010101",
7863 => "0000000010010101",
7864 => "0000000010010101",
7865 => "0000000010010101",
7866 => "0000000010010101",
7867 => "0000000010010101",
7868 => "0000000010010101",
7869 => "0000000010010101",
7870 => "0000000010010101",
7871 => "0000000010010101",
7872 => "0000000010010101",
7873 => "0000000010010101",
7874 => "0000000010010101",
7875 => "0000000010010110",
7876 => "0000000010010110",
7877 => "0000000010010110",
7878 => "0000000010010110",
7879 => "0000000010010110",
7880 => "0000000010010110",
7881 => "0000000010010110",
7882 => "0000000010010110",
7883 => "0000000010010110",
7884 => "0000000010010110",
7885 => "0000000010010110",
7886 => "0000000010010110",
7887 => "0000000010010110",
7888 => "0000000010010110",
7889 => "0000000010010110",
7890 => "0000000010010110",
7891 => "0000000010010110",
7892 => "0000000010010110",
7893 => "0000000010010110",
7894 => "0000000010010110",
7895 => "0000000010010110",
7896 => "0000000010010110",
7897 => "0000000010010110",
7898 => "0000000010010110",
7899 => "0000000010010110",
7900 => "0000000010010110",
7901 => "0000000010010110",
7902 => "0000000010010110",
7903 => "0000000010010111",
7904 => "0000000010010111",
7905 => "0000000010010111",
7906 => "0000000010010111",
7907 => "0000000010010111",
7908 => "0000000010010111",
7909 => "0000000010010111",
7910 => "0000000010010111",
7911 => "0000000010010111",
7912 => "0000000010010111",
7913 => "0000000010010111",
7914 => "0000000010010111",
7915 => "0000000010010111",
7916 => "0000000010010111",
7917 => "0000000010010111",
7918 => "0000000010010111",
7919 => "0000000010010111",
7920 => "0000000010010111",
7921 => "0000000010010111",
7922 => "0000000010010111",
7923 => "0000000010010111",
7924 => "0000000010010111",
7925 => "0000000010010111",
7926 => "0000000010010111",
7927 => "0000000010010111",
7928 => "0000000010010111",
7929 => "0000000010010111",
7930 => "0000000010011000",
7931 => "0000000010011000",
7932 => "0000000010011000",
7933 => "0000000010011000",
7934 => "0000000010011000",
7935 => "0000000010011000",
7936 => "0000000010011000",
7937 => "0000000010011000",
7938 => "0000000010011000",
7939 => "0000000010011000",
7940 => "0000000010011000",
7941 => "0000000010011000",
7942 => "0000000010011000",
7943 => "0000000010011000",
7944 => "0000000010011000",
7945 => "0000000010011000",
7946 => "0000000010011000",
7947 => "0000000010011000",
7948 => "0000000010011000",
7949 => "0000000010011000",
7950 => "0000000010011000",
7951 => "0000000010011000",
7952 => "0000000010011000",
7953 => "0000000010011000",
7954 => "0000000010011000",
7955 => "0000000010011000",
7956 => "0000000010011000",
7957 => "0000000010011001",
7958 => "0000000010011001",
7959 => "0000000010011001",
7960 => "0000000010011001",
7961 => "0000000010011001",
7962 => "0000000010011001",
7963 => "0000000010011001",
7964 => "0000000010011001",
7965 => "0000000010011001",
7966 => "0000000010011001",
7967 => "0000000010011001",
7968 => "0000000010011001",
7969 => "0000000010011001",
7970 => "0000000010011001",
7971 => "0000000010011001",
7972 => "0000000010011001",
7973 => "0000000010011001",
7974 => "0000000010011001",
7975 => "0000000010011001",
7976 => "0000000010011001",
7977 => "0000000010011001",
7978 => "0000000010011001",
7979 => "0000000010011001",
7980 => "0000000010011001",
7981 => "0000000010011001",
7982 => "0000000010011001",
7983 => "0000000010011010",
7984 => "0000000010011010",
7985 => "0000000010011010",
7986 => "0000000010011010",
7987 => "0000000010011010",
7988 => "0000000010011010",
7989 => "0000000010011010",
7990 => "0000000010011010",
7991 => "0000000010011010",
7992 => "0000000010011010",
7993 => "0000000010011010",
7994 => "0000000010011010",
7995 => "0000000010011010",
7996 => "0000000010011010",
7997 => "0000000010011010",
7998 => "0000000010011010",
7999 => "0000000010011010",
8000 => "0000000010011010",
8001 => "0000000010011010",
8002 => "0000000010011010",
8003 => "0000000010011010",
8004 => "0000000010011010",
8005 => "0000000010011010",
8006 => "0000000010011010",
8007 => "0000000010011010",
8008 => "0000000010011010",
8009 => "0000000010011010",
8010 => "0000000010011011",
8011 => "0000000010011011",
8012 => "0000000010011011",
8013 => "0000000010011011",
8014 => "0000000010011011",
8015 => "0000000010011011",
8016 => "0000000010011011",
8017 => "0000000010011011",
8018 => "0000000010011011",
8019 => "0000000010011011",
8020 => "0000000010011011",
8021 => "0000000010011011",
8022 => "0000000010011011",
8023 => "0000000010011011",
8024 => "0000000010011011",
8025 => "0000000010011011",
8026 => "0000000010011011",
8027 => "0000000010011011",
8028 => "0000000010011011",
8029 => "0000000010011011",
8030 => "0000000010011011",
8031 => "0000000010011011",
8032 => "0000000010011011",
8033 => "0000000010011011",
8034 => "0000000010011011",
8035 => "0000000010011011",
8036 => "0000000010011100",
8037 => "0000000010011100",
8038 => "0000000010011100",
8039 => "0000000010011100",
8040 => "0000000010011100",
8041 => "0000000010011100",
8042 => "0000000010011100",
8043 => "0000000010011100",
8044 => "0000000010011100",
8045 => "0000000010011100",
8046 => "0000000010011100",
8047 => "0000000010011100",
8048 => "0000000010011100",
8049 => "0000000010011100",
8050 => "0000000010011100",
8051 => "0000000010011100",
8052 => "0000000010011100",
8053 => "0000000010011100",
8054 => "0000000010011100",
8055 => "0000000010011100",
8056 => "0000000010011100",
8057 => "0000000010011100",
8058 => "0000000010011100",
8059 => "0000000010011100",
8060 => "0000000010011100",
8061 => "0000000010011100",
8062 => "0000000010011101",
8063 => "0000000010011101",
8064 => "0000000010011101",
8065 => "0000000010011101",
8066 => "0000000010011101",
8067 => "0000000010011101",
8068 => "0000000010011101",
8069 => "0000000010011101",
8070 => "0000000010011101",
8071 => "0000000010011101",
8072 => "0000000010011101",
8073 => "0000000010011101",
8074 => "0000000010011101",
8075 => "0000000010011101",
8076 => "0000000010011101",
8077 => "0000000010011101",
8078 => "0000000010011101",
8079 => "0000000010011101",
8080 => "0000000010011101",
8081 => "0000000010011101",
8082 => "0000000010011101",
8083 => "0000000010011101",
8084 => "0000000010011101",
8085 => "0000000010011101",
8086 => "0000000010011101",
8087 => "0000000010011101",
8088 => "0000000010011101",
8089 => "0000000010011110",
8090 => "0000000010011110",
8091 => "0000000010011110",
8092 => "0000000010011110",
8093 => "0000000010011110",
8094 => "0000000010011110",
8095 => "0000000010011110",
8096 => "0000000010011110",
8097 => "0000000010011110",
8098 => "0000000010011110",
8099 => "0000000010011110",
8100 => "0000000010011110",
8101 => "0000000010011110",
8102 => "0000000010011110",
8103 => "0000000010011110",
8104 => "0000000010011110",
8105 => "0000000010011110",
8106 => "0000000010011110",
8107 => "0000000010011110",
8108 => "0000000010011110",
8109 => "0000000010011110",
8110 => "0000000010011110",
8111 => "0000000010011110",
8112 => "0000000010011110",
8113 => "0000000010011110",
8114 => "0000000010011111",
8115 => "0000000010011111",
8116 => "0000000010011111",
8117 => "0000000010011111",
8118 => "0000000010011111",
8119 => "0000000010011111",
8120 => "0000000010011111",
8121 => "0000000010011111",
8122 => "0000000010011111",
8123 => "0000000010011111",
8124 => "0000000010011111",
8125 => "0000000010011111",
8126 => "0000000010011111",
8127 => "0000000010011111",
8128 => "0000000010011111",
8129 => "0000000010011111",
8130 => "0000000010011111",
8131 => "0000000010011111",
8132 => "0000000010011111",
8133 => "0000000010011111",
8134 => "0000000010011111",
8135 => "0000000010011111",
8136 => "0000000010011111",
8137 => "0000000010011111",
8138 => "0000000010011111",
8139 => "0000000010011111",
8140 => "0000000010100000",
8141 => "0000000010100000",
8142 => "0000000010100000",
8143 => "0000000010100000",
8144 => "0000000010100000",
8145 => "0000000010100000",
8146 => "0000000010100000",
8147 => "0000000010100000",
8148 => "0000000010100000",
8149 => "0000000010100000",
8150 => "0000000010100000",
8151 => "0000000010100000",
8152 => "0000000010100000",
8153 => "0000000010100000",
8154 => "0000000010100000",
8155 => "0000000010100000",
8156 => "0000000010100000",
8157 => "0000000010100000",
8158 => "0000000010100000",
8159 => "0000000010100000",
8160 => "0000000010100000",
8161 => "0000000010100000",
8162 => "0000000010100000",
8163 => "0000000010100000",
8164 => "0000000010100000",
8165 => "0000000010100000",
8166 => "0000000010100001",
8167 => "0000000010100001",
8168 => "0000000010100001",
8169 => "0000000010100001",
8170 => "0000000010100001",
8171 => "0000000010100001",
8172 => "0000000010100001",
8173 => "0000000010100001",
8174 => "0000000010100001",
8175 => "0000000010100001",
8176 => "0000000010100001",
8177 => "0000000010100001",
8178 => "0000000010100001",
8179 => "0000000010100001",
8180 => "0000000010100001",
8181 => "0000000010100001",
8182 => "0000000010100001",
8183 => "0000000010100001",
8184 => "0000000010100001",
8185 => "0000000010100001",
8186 => "0000000010100001",
8187 => "0000000010100001",
8188 => "0000000010100001",
8189 => "0000000010100001",
8190 => "0000000010100001",
8191 => "0000000010100010",
8192 => "0000000010100010",
8193 => "0000000010100010",
8194 => "0000000010100010",
8195 => "0000000010100010",
8196 => "0000000010100010",
8197 => "0000000010100010",
8198 => "0000000010100010",
8199 => "0000000010100010",
8200 => "0000000010100010",
8201 => "0000000010100010",
8202 => "0000000010100010",
8203 => "0000000010100010",
8204 => "0000000010100010",
8205 => "0000000010100010",
8206 => "0000000010100010",
8207 => "0000000010100010",
8208 => "0000000010100010",
8209 => "0000000010100010",
8210 => "0000000010100010",
8211 => "0000000010100010",
8212 => "0000000010100010",
8213 => "0000000010100010",
8214 => "0000000010100010",
8215 => "0000000010100010",
8216 => "0000000010100011",
8217 => "0000000010100011",
8218 => "0000000010100011",
8219 => "0000000010100011",
8220 => "0000000010100011",
8221 => "0000000010100011",
8222 => "0000000010100011",
8223 => "0000000010100011",
8224 => "0000000010100011",
8225 => "0000000010100011",
8226 => "0000000010100011",
8227 => "0000000010100011",
8228 => "0000000010100011",
8229 => "0000000010100011",
8230 => "0000000010100011",
8231 => "0000000010100011",
8232 => "0000000010100011",
8233 => "0000000010100011",
8234 => "0000000010100011",
8235 => "0000000010100011",
8236 => "0000000010100011",
8237 => "0000000010100011",
8238 => "0000000010100011",
8239 => "0000000010100011",
8240 => "0000000010100011",
8241 => "0000000010100011",
8242 => "0000000010100100",
8243 => "0000000010100100",
8244 => "0000000010100100",
8245 => "0000000010100100",
8246 => "0000000010100100",
8247 => "0000000010100100",
8248 => "0000000010100100",
8249 => "0000000010100100",
8250 => "0000000010100100",
8251 => "0000000010100100",
8252 => "0000000010100100",
8253 => "0000000010100100",
8254 => "0000000010100100",
8255 => "0000000010100100",
8256 => "0000000010100100",
8257 => "0000000010100100",
8258 => "0000000010100100",
8259 => "0000000010100100",
8260 => "0000000010100100",
8261 => "0000000010100100",
8262 => "0000000010100100",
8263 => "0000000010100100",
8264 => "0000000010100100",
8265 => "0000000010100100",
8266 => "0000000010100100",
8267 => "0000000010100101",
8268 => "0000000010100101",
8269 => "0000000010100101",
8270 => "0000000010100101",
8271 => "0000000010100101",
8272 => "0000000010100101",
8273 => "0000000010100101",
8274 => "0000000010100101",
8275 => "0000000010100101",
8276 => "0000000010100101",
8277 => "0000000010100101",
8278 => "0000000010100101",
8279 => "0000000010100101",
8280 => "0000000010100101",
8281 => "0000000010100101",
8282 => "0000000010100101",
8283 => "0000000010100101",
8284 => "0000000010100101",
8285 => "0000000010100101",
8286 => "0000000010100101",
8287 => "0000000010100101",
8288 => "0000000010100101",
8289 => "0000000010100101",
8290 => "0000000010100101",
8291 => "0000000010100110",
8292 => "0000000010100110",
8293 => "0000000010100110",
8294 => "0000000010100110",
8295 => "0000000010100110",
8296 => "0000000010100110",
8297 => "0000000010100110",
8298 => "0000000010100110",
8299 => "0000000010100110",
8300 => "0000000010100110",
8301 => "0000000010100110",
8302 => "0000000010100110",
8303 => "0000000010100110",
8304 => "0000000010100110",
8305 => "0000000010100110",
8306 => "0000000010100110",
8307 => "0000000010100110",
8308 => "0000000010100110",
8309 => "0000000010100110",
8310 => "0000000010100110",
8311 => "0000000010100110",
8312 => "0000000010100110",
8313 => "0000000010100110",
8314 => "0000000010100110",
8315 => "0000000010100110",
8316 => "0000000010100111",
8317 => "0000000010100111",
8318 => "0000000010100111",
8319 => "0000000010100111",
8320 => "0000000010100111",
8321 => "0000000010100111",
8322 => "0000000010100111",
8323 => "0000000010100111",
8324 => "0000000010100111",
8325 => "0000000010100111",
8326 => "0000000010100111",
8327 => "0000000010100111",
8328 => "0000000010100111",
8329 => "0000000010100111",
8330 => "0000000010100111",
8331 => "0000000010100111",
8332 => "0000000010100111",
8333 => "0000000010100111",
8334 => "0000000010100111",
8335 => "0000000010100111",
8336 => "0000000010100111",
8337 => "0000000010100111",
8338 => "0000000010100111",
8339 => "0000000010100111",
8340 => "0000000010100111",
8341 => "0000000010101000",
8342 => "0000000010101000",
8343 => "0000000010101000",
8344 => "0000000010101000",
8345 => "0000000010101000",
8346 => "0000000010101000",
8347 => "0000000010101000",
8348 => "0000000010101000",
8349 => "0000000010101000",
8350 => "0000000010101000",
8351 => "0000000010101000",
8352 => "0000000010101000",
8353 => "0000000010101000",
8354 => "0000000010101000",
8355 => "0000000010101000",
8356 => "0000000010101000",
8357 => "0000000010101000",
8358 => "0000000010101000",
8359 => "0000000010101000",
8360 => "0000000010101000",
8361 => "0000000010101000",
8362 => "0000000010101000",
8363 => "0000000010101000",
8364 => "0000000010101000",
8365 => "0000000010101001",
8366 => "0000000010101001",
8367 => "0000000010101001",
8368 => "0000000010101001",
8369 => "0000000010101001",
8370 => "0000000010101001",
8371 => "0000000010101001",
8372 => "0000000010101001",
8373 => "0000000010101001",
8374 => "0000000010101001",
8375 => "0000000010101001",
8376 => "0000000010101001",
8377 => "0000000010101001",
8378 => "0000000010101001",
8379 => "0000000010101001",
8380 => "0000000010101001",
8381 => "0000000010101001",
8382 => "0000000010101001",
8383 => "0000000010101001",
8384 => "0000000010101001",
8385 => "0000000010101001",
8386 => "0000000010101001",
8387 => "0000000010101001",
8388 => "0000000010101001",
8389 => "0000000010101010",
8390 => "0000000010101010",
8391 => "0000000010101010",
8392 => "0000000010101010",
8393 => "0000000010101010",
8394 => "0000000010101010",
8395 => "0000000010101010",
8396 => "0000000010101010",
8397 => "0000000010101010",
8398 => "0000000010101010",
8399 => "0000000010101010",
8400 => "0000000010101010",
8401 => "0000000010101010",
8402 => "0000000010101010",
8403 => "0000000010101010",
8404 => "0000000010101010",
8405 => "0000000010101010",
8406 => "0000000010101010",
8407 => "0000000010101010",
8408 => "0000000010101010",
8409 => "0000000010101010",
8410 => "0000000010101010",
8411 => "0000000010101010",
8412 => "0000000010101010",
8413 => "0000000010101011",
8414 => "0000000010101011",
8415 => "0000000010101011",
8416 => "0000000010101011",
8417 => "0000000010101011",
8418 => "0000000010101011",
8419 => "0000000010101011",
8420 => "0000000010101011",
8421 => "0000000010101011",
8422 => "0000000010101011",
8423 => "0000000010101011",
8424 => "0000000010101011",
8425 => "0000000010101011",
8426 => "0000000010101011",
8427 => "0000000010101011",
8428 => "0000000010101011",
8429 => "0000000010101011",
8430 => "0000000010101011",
8431 => "0000000010101011",
8432 => "0000000010101011",
8433 => "0000000010101011",
8434 => "0000000010101011",
8435 => "0000000010101011",
8436 => "0000000010101011",
8437 => "0000000010101100",
8438 => "0000000010101100",
8439 => "0000000010101100",
8440 => "0000000010101100",
8441 => "0000000010101100",
8442 => "0000000010101100",
8443 => "0000000010101100",
8444 => "0000000010101100",
8445 => "0000000010101100",
8446 => "0000000010101100",
8447 => "0000000010101100",
8448 => "0000000010101100",
8449 => "0000000010101100",
8450 => "0000000010101100",
8451 => "0000000010101100",
8452 => "0000000010101100",
8453 => "0000000010101100",
8454 => "0000000010101100",
8455 => "0000000010101100",
8456 => "0000000010101100",
8457 => "0000000010101100",
8458 => "0000000010101100",
8459 => "0000000010101100",
8460 => "0000000010101100",
8461 => "0000000010101101",
8462 => "0000000010101101",
8463 => "0000000010101101",
8464 => "0000000010101101",
8465 => "0000000010101101",
8466 => "0000000010101101",
8467 => "0000000010101101",
8468 => "0000000010101101",
8469 => "0000000010101101",
8470 => "0000000010101101",
8471 => "0000000010101101",
8472 => "0000000010101101",
8473 => "0000000010101101",
8474 => "0000000010101101",
8475 => "0000000010101101",
8476 => "0000000010101101",
8477 => "0000000010101101",
8478 => "0000000010101101",
8479 => "0000000010101101",
8480 => "0000000010101101",
8481 => "0000000010101101",
8482 => "0000000010101101",
8483 => "0000000010101101",
8484 => "0000000010101101",
8485 => "0000000010101110",
8486 => "0000000010101110",
8487 => "0000000010101110",
8488 => "0000000010101110",
8489 => "0000000010101110",
8490 => "0000000010101110",
8491 => "0000000010101110",
8492 => "0000000010101110",
8493 => "0000000010101110",
8494 => "0000000010101110",
8495 => "0000000010101110",
8496 => "0000000010101110",
8497 => "0000000010101110",
8498 => "0000000010101110",
8499 => "0000000010101110",
8500 => "0000000010101110",
8501 => "0000000010101110",
8502 => "0000000010101110",
8503 => "0000000010101110",
8504 => "0000000010101110",
8505 => "0000000010101110",
8506 => "0000000010101110",
8507 => "0000000010101110",
8508 => "0000000010101111",
8509 => "0000000010101111",
8510 => "0000000010101111",
8511 => "0000000010101111",
8512 => "0000000010101111",
8513 => "0000000010101111",
8514 => "0000000010101111",
8515 => "0000000010101111",
8516 => "0000000010101111",
8517 => "0000000010101111",
8518 => "0000000010101111",
8519 => "0000000010101111",
8520 => "0000000010101111",
8521 => "0000000010101111",
8522 => "0000000010101111",
8523 => "0000000010101111",
8524 => "0000000010101111",
8525 => "0000000010101111",
8526 => "0000000010101111",
8527 => "0000000010101111",
8528 => "0000000010101111",
8529 => "0000000010101111",
8530 => "0000000010101111",
8531 => "0000000010101111",
8532 => "0000000010110000",
8533 => "0000000010110000",
8534 => "0000000010110000",
8535 => "0000000010110000",
8536 => "0000000010110000",
8537 => "0000000010110000",
8538 => "0000000010110000",
8539 => "0000000010110000",
8540 => "0000000010110000",
8541 => "0000000010110000",
8542 => "0000000010110000",
8543 => "0000000010110000",
8544 => "0000000010110000",
8545 => "0000000010110000",
8546 => "0000000010110000",
8547 => "0000000010110000",
8548 => "0000000010110000",
8549 => "0000000010110000",
8550 => "0000000010110000",
8551 => "0000000010110000",
8552 => "0000000010110000",
8553 => "0000000010110000",
8554 => "0000000010110000",
8555 => "0000000010110001",
8556 => "0000000010110001",
8557 => "0000000010110001",
8558 => "0000000010110001",
8559 => "0000000010110001",
8560 => "0000000010110001",
8561 => "0000000010110001",
8562 => "0000000010110001",
8563 => "0000000010110001",
8564 => "0000000010110001",
8565 => "0000000010110001",
8566 => "0000000010110001",
8567 => "0000000010110001",
8568 => "0000000010110001",
8569 => "0000000010110001",
8570 => "0000000010110001",
8571 => "0000000010110001",
8572 => "0000000010110001",
8573 => "0000000010110001",
8574 => "0000000010110001",
8575 => "0000000010110001",
8576 => "0000000010110001",
8577 => "0000000010110001",
8578 => "0000000010110010",
8579 => "0000000010110010",
8580 => "0000000010110010",
8581 => "0000000010110010",
8582 => "0000000010110010",
8583 => "0000000010110010",
8584 => "0000000010110010",
8585 => "0000000010110010",
8586 => "0000000010110010",
8587 => "0000000010110010",
8588 => "0000000010110010",
8589 => "0000000010110010",
8590 => "0000000010110010",
8591 => "0000000010110010",
8592 => "0000000010110010",
8593 => "0000000010110010",
8594 => "0000000010110010",
8595 => "0000000010110010",
8596 => "0000000010110010",
8597 => "0000000010110010",
8598 => "0000000010110010",
8599 => "0000000010110010",
8600 => "0000000010110010",
8601 => "0000000010110011",
8602 => "0000000010110011",
8603 => "0000000010110011",
8604 => "0000000010110011",
8605 => "0000000010110011",
8606 => "0000000010110011",
8607 => "0000000010110011",
8608 => "0000000010110011",
8609 => "0000000010110011",
8610 => "0000000010110011",
8611 => "0000000010110011",
8612 => "0000000010110011",
8613 => "0000000010110011",
8614 => "0000000010110011",
8615 => "0000000010110011",
8616 => "0000000010110011",
8617 => "0000000010110011",
8618 => "0000000010110011",
8619 => "0000000010110011",
8620 => "0000000010110011",
8621 => "0000000010110011",
8622 => "0000000010110011",
8623 => "0000000010110011",
8624 => "0000000010110100",
8625 => "0000000010110100",
8626 => "0000000010110100",
8627 => "0000000010110100",
8628 => "0000000010110100",
8629 => "0000000010110100",
8630 => "0000000010110100",
8631 => "0000000010110100",
8632 => "0000000010110100",
8633 => "0000000010110100",
8634 => "0000000010110100",
8635 => "0000000010110100",
8636 => "0000000010110100",
8637 => "0000000010110100",
8638 => "0000000010110100",
8639 => "0000000010110100",
8640 => "0000000010110100",
8641 => "0000000010110100",
8642 => "0000000010110100",
8643 => "0000000010110100",
8644 => "0000000010110100",
8645 => "0000000010110100",
8646 => "0000000010110100",
8647 => "0000000010110101",
8648 => "0000000010110101",
8649 => "0000000010110101",
8650 => "0000000010110101",
8651 => "0000000010110101",
8652 => "0000000010110101",
8653 => "0000000010110101",
8654 => "0000000010110101",
8655 => "0000000010110101",
8656 => "0000000010110101",
8657 => "0000000010110101",
8658 => "0000000010110101",
8659 => "0000000010110101",
8660 => "0000000010110101",
8661 => "0000000010110101",
8662 => "0000000010110101",
8663 => "0000000010110101",
8664 => "0000000010110101",
8665 => "0000000010110101",
8666 => "0000000010110101",
8667 => "0000000010110101",
8668 => "0000000010110101",
8669 => "0000000010110110",
8670 => "0000000010110110",
8671 => "0000000010110110",
8672 => "0000000010110110",
8673 => "0000000010110110",
8674 => "0000000010110110",
8675 => "0000000010110110",
8676 => "0000000010110110",
8677 => "0000000010110110",
8678 => "0000000010110110",
8679 => "0000000010110110",
8680 => "0000000010110110",
8681 => "0000000010110110",
8682 => "0000000010110110",
8683 => "0000000010110110",
8684 => "0000000010110110",
8685 => "0000000010110110",
8686 => "0000000010110110",
8687 => "0000000010110110",
8688 => "0000000010110110",
8689 => "0000000010110110",
8690 => "0000000010110110",
8691 => "0000000010110110",
8692 => "0000000010110111",
8693 => "0000000010110111",
8694 => "0000000010110111",
8695 => "0000000010110111",
8696 => "0000000010110111",
8697 => "0000000010110111",
8698 => "0000000010110111",
8699 => "0000000010110111",
8700 => "0000000010110111",
8701 => "0000000010110111",
8702 => "0000000010110111",
8703 => "0000000010110111",
8704 => "0000000010110111",
8705 => "0000000010110111",
8706 => "0000000010110111",
8707 => "0000000010110111",
8708 => "0000000010110111",
8709 => "0000000010110111",
8710 => "0000000010110111",
8711 => "0000000010110111",
8712 => "0000000010110111",
8713 => "0000000010110111",
8714 => "0000000010111000",
8715 => "0000000010111000",
8716 => "0000000010111000",
8717 => "0000000010111000",
8718 => "0000000010111000",
8719 => "0000000010111000",
8720 => "0000000010111000",
8721 => "0000000010111000",
8722 => "0000000010111000",
8723 => "0000000010111000",
8724 => "0000000010111000",
8725 => "0000000010111000",
8726 => "0000000010111000",
8727 => "0000000010111000",
8728 => "0000000010111000",
8729 => "0000000010111000",
8730 => "0000000010111000",
8731 => "0000000010111000",
8732 => "0000000010111000",
8733 => "0000000010111000",
8734 => "0000000010111000",
8735 => "0000000010111000",
8736 => "0000000010111001",
8737 => "0000000010111001",
8738 => "0000000010111001",
8739 => "0000000010111001",
8740 => "0000000010111001",
8741 => "0000000010111001",
8742 => "0000000010111001",
8743 => "0000000010111001",
8744 => "0000000010111001",
8745 => "0000000010111001",
8746 => "0000000010111001",
8747 => "0000000010111001",
8748 => "0000000010111001",
8749 => "0000000010111001",
8750 => "0000000010111001",
8751 => "0000000010111001",
8752 => "0000000010111001",
8753 => "0000000010111001",
8754 => "0000000010111001",
8755 => "0000000010111001",
8756 => "0000000010111001",
8757 => "0000000010111001",
8758 => "0000000010111001",
8759 => "0000000010111010",
8760 => "0000000010111010",
8761 => "0000000010111010",
8762 => "0000000010111010",
8763 => "0000000010111010",
8764 => "0000000010111010",
8765 => "0000000010111010",
8766 => "0000000010111010",
8767 => "0000000010111010",
8768 => "0000000010111010",
8769 => "0000000010111010",
8770 => "0000000010111010",
8771 => "0000000010111010",
8772 => "0000000010111010",
8773 => "0000000010111010",
8774 => "0000000010111010",
8775 => "0000000010111010",
8776 => "0000000010111010",
8777 => "0000000010111010",
8778 => "0000000010111010",
8779 => "0000000010111010",
8780 => "0000000010111010",
8781 => "0000000010111011",
8782 => "0000000010111011",
8783 => "0000000010111011",
8784 => "0000000010111011",
8785 => "0000000010111011",
8786 => "0000000010111011",
8787 => "0000000010111011",
8788 => "0000000010111011",
8789 => "0000000010111011",
8790 => "0000000010111011",
8791 => "0000000010111011",
8792 => "0000000010111011",
8793 => "0000000010111011",
8794 => "0000000010111011",
8795 => "0000000010111011",
8796 => "0000000010111011",
8797 => "0000000010111011",
8798 => "0000000010111011",
8799 => "0000000010111011",
8800 => "0000000010111011",
8801 => "0000000010111011",
8802 => "0000000010111011",
8803 => "0000000010111100",
8804 => "0000000010111100",
8805 => "0000000010111100",
8806 => "0000000010111100",
8807 => "0000000010111100",
8808 => "0000000010111100",
8809 => "0000000010111100",
8810 => "0000000010111100",
8811 => "0000000010111100",
8812 => "0000000010111100",
8813 => "0000000010111100",
8814 => "0000000010111100",
8815 => "0000000010111100",
8816 => "0000000010111100",
8817 => "0000000010111100",
8818 => "0000000010111100",
8819 => "0000000010111100",
8820 => "0000000010111100",
8821 => "0000000010111100",
8822 => "0000000010111100",
8823 => "0000000010111100",
8824 => "0000000010111101",
8825 => "0000000010111101",
8826 => "0000000010111101",
8827 => "0000000010111101",
8828 => "0000000010111101",
8829 => "0000000010111101",
8830 => "0000000010111101",
8831 => "0000000010111101",
8832 => "0000000010111101",
8833 => "0000000010111101",
8834 => "0000000010111101",
8835 => "0000000010111101",
8836 => "0000000010111101",
8837 => "0000000010111101",
8838 => "0000000010111101",
8839 => "0000000010111101",
8840 => "0000000010111101",
8841 => "0000000010111101",
8842 => "0000000010111101",
8843 => "0000000010111101",
8844 => "0000000010111101",
8845 => "0000000010111101",
8846 => "0000000010111110",
8847 => "0000000010111110",
8848 => "0000000010111110",
8849 => "0000000010111110",
8850 => "0000000010111110",
8851 => "0000000010111110",
8852 => "0000000010111110",
8853 => "0000000010111110",
8854 => "0000000010111110",
8855 => "0000000010111110",
8856 => "0000000010111110",
8857 => "0000000010111110",
8858 => "0000000010111110",
8859 => "0000000010111110",
8860 => "0000000010111110",
8861 => "0000000010111110",
8862 => "0000000010111110",
8863 => "0000000010111110",
8864 => "0000000010111110",
8865 => "0000000010111110",
8866 => "0000000010111110",
8867 => "0000000010111110",
8868 => "0000000010111111",
8869 => "0000000010111111",
8870 => "0000000010111111",
8871 => "0000000010111111",
8872 => "0000000010111111",
8873 => "0000000010111111",
8874 => "0000000010111111",
8875 => "0000000010111111",
8876 => "0000000010111111",
8877 => "0000000010111111",
8878 => "0000000010111111",
8879 => "0000000010111111",
8880 => "0000000010111111",
8881 => "0000000010111111",
8882 => "0000000010111111",
8883 => "0000000010111111",
8884 => "0000000010111111",
8885 => "0000000010111111",
8886 => "0000000010111111",
8887 => "0000000010111111",
8888 => "0000000010111111",
8889 => "0000000011000000",
8890 => "0000000011000000",
8891 => "0000000011000000",
8892 => "0000000011000000",
8893 => "0000000011000000",
8894 => "0000000011000000",
8895 => "0000000011000000",
8896 => "0000000011000000",
8897 => "0000000011000000",
8898 => "0000000011000000",
8899 => "0000000011000000",
8900 => "0000000011000000",
8901 => "0000000011000000",
8902 => "0000000011000000",
8903 => "0000000011000000",
8904 => "0000000011000000",
8905 => "0000000011000000",
8906 => "0000000011000000",
8907 => "0000000011000000",
8908 => "0000000011000000",
8909 => "0000000011000000",
8910 => "0000000011000001",
8911 => "0000000011000001",
8912 => "0000000011000001",
8913 => "0000000011000001",
8914 => "0000000011000001",
8915 => "0000000011000001",
8916 => "0000000011000001",
8917 => "0000000011000001",
8918 => "0000000011000001",
8919 => "0000000011000001",
8920 => "0000000011000001",
8921 => "0000000011000001",
8922 => "0000000011000001",
8923 => "0000000011000001",
8924 => "0000000011000001",
8925 => "0000000011000001",
8926 => "0000000011000001",
8927 => "0000000011000001",
8928 => "0000000011000001",
8929 => "0000000011000001",
8930 => "0000000011000001",
8931 => "0000000011000001",
8932 => "0000000011000010",
8933 => "0000000011000010",
8934 => "0000000011000010",
8935 => "0000000011000010",
8936 => "0000000011000010",
8937 => "0000000011000010",
8938 => "0000000011000010",
8939 => "0000000011000010",
8940 => "0000000011000010",
8941 => "0000000011000010",
8942 => "0000000011000010",
8943 => "0000000011000010",
8944 => "0000000011000010",
8945 => "0000000011000010",
8946 => "0000000011000010",
8947 => "0000000011000010",
8948 => "0000000011000010",
8949 => "0000000011000010",
8950 => "0000000011000010",
8951 => "0000000011000010",
8952 => "0000000011000010",
8953 => "0000000011000011",
8954 => "0000000011000011",
8955 => "0000000011000011",
8956 => "0000000011000011",
8957 => "0000000011000011",
8958 => "0000000011000011",
8959 => "0000000011000011",
8960 => "0000000011000011",
8961 => "0000000011000011",
8962 => "0000000011000011",
8963 => "0000000011000011",
8964 => "0000000011000011",
8965 => "0000000011000011",
8966 => "0000000011000011",
8967 => "0000000011000011",
8968 => "0000000011000011",
8969 => "0000000011000011",
8970 => "0000000011000011",
8971 => "0000000011000011",
8972 => "0000000011000011",
8973 => "0000000011000011",
8974 => "0000000011000100",
8975 => "0000000011000100",
8976 => "0000000011000100",
8977 => "0000000011000100",
8978 => "0000000011000100",
8979 => "0000000011000100",
8980 => "0000000011000100",
8981 => "0000000011000100",
8982 => "0000000011000100",
8983 => "0000000011000100",
8984 => "0000000011000100",
8985 => "0000000011000100",
8986 => "0000000011000100",
8987 => "0000000011000100",
8988 => "0000000011000100",
8989 => "0000000011000100",
8990 => "0000000011000100",
8991 => "0000000011000100",
8992 => "0000000011000100",
8993 => "0000000011000100",
8994 => "0000000011000100",
8995 => "0000000011000101",
8996 => "0000000011000101",
8997 => "0000000011000101",
8998 => "0000000011000101",
8999 => "0000000011000101",
9000 => "0000000011000101",
9001 => "0000000011000101",
9002 => "0000000011000101",
9003 => "0000000011000101",
9004 => "0000000011000101",
9005 => "0000000011000101",
9006 => "0000000011000101",
9007 => "0000000011000101",
9008 => "0000000011000101",
9009 => "0000000011000101",
9010 => "0000000011000101",
9011 => "0000000011000101",
9012 => "0000000011000101",
9013 => "0000000011000101",
9014 => "0000000011000101",
9015 => "0000000011000110",
9016 => "0000000011000110",
9017 => "0000000011000110",
9018 => "0000000011000110",
9019 => "0000000011000110",
9020 => "0000000011000110",
9021 => "0000000011000110",
9022 => "0000000011000110",
9023 => "0000000011000110",
9024 => "0000000011000110",
9025 => "0000000011000110",
9026 => "0000000011000110",
9027 => "0000000011000110",
9028 => "0000000011000110",
9029 => "0000000011000110",
9030 => "0000000011000110",
9031 => "0000000011000110",
9032 => "0000000011000110",
9033 => "0000000011000110",
9034 => "0000000011000110",
9035 => "0000000011000110",
9036 => "0000000011000111",
9037 => "0000000011000111",
9038 => "0000000011000111",
9039 => "0000000011000111",
9040 => "0000000011000111",
9041 => "0000000011000111",
9042 => "0000000011000111",
9043 => "0000000011000111",
9044 => "0000000011000111",
9045 => "0000000011000111",
9046 => "0000000011000111",
9047 => "0000000011000111",
9048 => "0000000011000111",
9049 => "0000000011000111",
9050 => "0000000011000111",
9051 => "0000000011000111",
9052 => "0000000011000111",
9053 => "0000000011000111",
9054 => "0000000011000111",
9055 => "0000000011000111",
9056 => "0000000011000111",
9057 => "0000000011001000",
9058 => "0000000011001000",
9059 => "0000000011001000",
9060 => "0000000011001000",
9061 => "0000000011001000",
9062 => "0000000011001000",
9063 => "0000000011001000",
9064 => "0000000011001000",
9065 => "0000000011001000",
9066 => "0000000011001000",
9067 => "0000000011001000",
9068 => "0000000011001000",
9069 => "0000000011001000",
9070 => "0000000011001000",
9071 => "0000000011001000",
9072 => "0000000011001000",
9073 => "0000000011001000",
9074 => "0000000011001000",
9075 => "0000000011001000",
9076 => "0000000011001000",
9077 => "0000000011001001",
9078 => "0000000011001001",
9079 => "0000000011001001",
9080 => "0000000011001001",
9081 => "0000000011001001",
9082 => "0000000011001001",
9083 => "0000000011001001",
9084 => "0000000011001001",
9085 => "0000000011001001",
9086 => "0000000011001001",
9087 => "0000000011001001",
9088 => "0000000011001001",
9089 => "0000000011001001",
9090 => "0000000011001001",
9091 => "0000000011001001",
9092 => "0000000011001001",
9093 => "0000000011001001",
9094 => "0000000011001001",
9095 => "0000000011001001",
9096 => "0000000011001001",
9097 => "0000000011001001",
9098 => "0000000011001010",
9099 => "0000000011001010",
9100 => "0000000011001010",
9101 => "0000000011001010",
9102 => "0000000011001010",
9103 => "0000000011001010",
9104 => "0000000011001010",
9105 => "0000000011001010",
9106 => "0000000011001010",
9107 => "0000000011001010",
9108 => "0000000011001010",
9109 => "0000000011001010",
9110 => "0000000011001010",
9111 => "0000000011001010",
9112 => "0000000011001010",
9113 => "0000000011001010",
9114 => "0000000011001010",
9115 => "0000000011001010",
9116 => "0000000011001010",
9117 => "0000000011001010",
9118 => "0000000011001011",
9119 => "0000000011001011",
9120 => "0000000011001011",
9121 => "0000000011001011",
9122 => "0000000011001011",
9123 => "0000000011001011",
9124 => "0000000011001011",
9125 => "0000000011001011",
9126 => "0000000011001011",
9127 => "0000000011001011",
9128 => "0000000011001011",
9129 => "0000000011001011",
9130 => "0000000011001011",
9131 => "0000000011001011",
9132 => "0000000011001011",
9133 => "0000000011001011",
9134 => "0000000011001011",
9135 => "0000000011001011",
9136 => "0000000011001011",
9137 => "0000000011001011",
9138 => "0000000011001100",
9139 => "0000000011001100",
9140 => "0000000011001100",
9141 => "0000000011001100",
9142 => "0000000011001100",
9143 => "0000000011001100",
9144 => "0000000011001100",
9145 => "0000000011001100",
9146 => "0000000011001100",
9147 => "0000000011001100",
9148 => "0000000011001100",
9149 => "0000000011001100",
9150 => "0000000011001100",
9151 => "0000000011001100",
9152 => "0000000011001100",
9153 => "0000000011001100",
9154 => "0000000011001100",
9155 => "0000000011001100",
9156 => "0000000011001100",
9157 => "0000000011001100",
9158 => "0000000011001101",
9159 => "0000000011001101",
9160 => "0000000011001101",
9161 => "0000000011001101",
9162 => "0000000011001101",
9163 => "0000000011001101",
9164 => "0000000011001101",
9165 => "0000000011001101",
9166 => "0000000011001101",
9167 => "0000000011001101",
9168 => "0000000011001101",
9169 => "0000000011001101",
9170 => "0000000011001101",
9171 => "0000000011001101",
9172 => "0000000011001101",
9173 => "0000000011001101",
9174 => "0000000011001101",
9175 => "0000000011001101",
9176 => "0000000011001101",
9177 => "0000000011001101",
9178 => "0000000011001110",
9179 => "0000000011001110",
9180 => "0000000011001110",
9181 => "0000000011001110",
9182 => "0000000011001110",
9183 => "0000000011001110",
9184 => "0000000011001110",
9185 => "0000000011001110",
9186 => "0000000011001110",
9187 => "0000000011001110",
9188 => "0000000011001110",
9189 => "0000000011001110",
9190 => "0000000011001110",
9191 => "0000000011001110",
9192 => "0000000011001110",
9193 => "0000000011001110",
9194 => "0000000011001110",
9195 => "0000000011001110",
9196 => "0000000011001110",
9197 => "0000000011001110",
9198 => "0000000011001111",
9199 => "0000000011001111",
9200 => "0000000011001111",
9201 => "0000000011001111",
9202 => "0000000011001111",
9203 => "0000000011001111",
9204 => "0000000011001111",
9205 => "0000000011001111",
9206 => "0000000011001111",
9207 => "0000000011001111",
9208 => "0000000011001111",
9209 => "0000000011001111",
9210 => "0000000011001111",
9211 => "0000000011001111",
9212 => "0000000011001111",
9213 => "0000000011001111",
9214 => "0000000011001111",
9215 => "0000000011001111",
9216 => "0000000011001111",
9217 => "0000000011001111",
9218 => "0000000011010000",
9219 => "0000000011010000",
9220 => "0000000011010000",
9221 => "0000000011010000",
9222 => "0000000011010000",
9223 => "0000000011010000",
9224 => "0000000011010000",
9225 => "0000000011010000",
9226 => "0000000011010000",
9227 => "0000000011010000",
9228 => "0000000011010000",
9229 => "0000000011010000",
9230 => "0000000011010000",
9231 => "0000000011010000",
9232 => "0000000011010000",
9233 => "0000000011010000",
9234 => "0000000011010000",
9235 => "0000000011010000",
9236 => "0000000011010000",
9237 => "0000000011010000",
9238 => "0000000011010001",
9239 => "0000000011010001",
9240 => "0000000011010001",
9241 => "0000000011010001",
9242 => "0000000011010001",
9243 => "0000000011010001",
9244 => "0000000011010001",
9245 => "0000000011010001",
9246 => "0000000011010001",
9247 => "0000000011010001",
9248 => "0000000011010001",
9249 => "0000000011010001",
9250 => "0000000011010001",
9251 => "0000000011010001",
9252 => "0000000011010001",
9253 => "0000000011010001",
9254 => "0000000011010001",
9255 => "0000000011010001",
9256 => "0000000011010001",
9257 => "0000000011010010",
9258 => "0000000011010010",
9259 => "0000000011010010",
9260 => "0000000011010010",
9261 => "0000000011010010",
9262 => "0000000011010010",
9263 => "0000000011010010",
9264 => "0000000011010010",
9265 => "0000000011010010",
9266 => "0000000011010010",
9267 => "0000000011010010",
9268 => "0000000011010010",
9269 => "0000000011010010",
9270 => "0000000011010010",
9271 => "0000000011010010",
9272 => "0000000011010010",
9273 => "0000000011010010",
9274 => "0000000011010010",
9275 => "0000000011010010",
9276 => "0000000011010010",
9277 => "0000000011010011",
9278 => "0000000011010011",
9279 => "0000000011010011",
9280 => "0000000011010011",
9281 => "0000000011010011",
9282 => "0000000011010011",
9283 => "0000000011010011",
9284 => "0000000011010011",
9285 => "0000000011010011",
9286 => "0000000011010011",
9287 => "0000000011010011",
9288 => "0000000011010011",
9289 => "0000000011010011",
9290 => "0000000011010011",
9291 => "0000000011010011",
9292 => "0000000011010011",
9293 => "0000000011010011",
9294 => "0000000011010011",
9295 => "0000000011010011",
9296 => "0000000011010100",
9297 => "0000000011010100",
9298 => "0000000011010100",
9299 => "0000000011010100",
9300 => "0000000011010100",
9301 => "0000000011010100",
9302 => "0000000011010100",
9303 => "0000000011010100",
9304 => "0000000011010100",
9305 => "0000000011010100",
9306 => "0000000011010100",
9307 => "0000000011010100",
9308 => "0000000011010100",
9309 => "0000000011010100",
9310 => "0000000011010100",
9311 => "0000000011010100",
9312 => "0000000011010100",
9313 => "0000000011010100",
9314 => "0000000011010100",
9315 => "0000000011010101",
9316 => "0000000011010101",
9317 => "0000000011010101",
9318 => "0000000011010101",
9319 => "0000000011010101",
9320 => "0000000011010101",
9321 => "0000000011010101",
9322 => "0000000011010101",
9323 => "0000000011010101",
9324 => "0000000011010101",
9325 => "0000000011010101",
9326 => "0000000011010101",
9327 => "0000000011010101",
9328 => "0000000011010101",
9329 => "0000000011010101",
9330 => "0000000011010101",
9331 => "0000000011010101",
9332 => "0000000011010101",
9333 => "0000000011010101",
9334 => "0000000011010101",
9335 => "0000000011010110",
9336 => "0000000011010110",
9337 => "0000000011010110",
9338 => "0000000011010110",
9339 => "0000000011010110",
9340 => "0000000011010110",
9341 => "0000000011010110",
9342 => "0000000011010110",
9343 => "0000000011010110",
9344 => "0000000011010110",
9345 => "0000000011010110",
9346 => "0000000011010110",
9347 => "0000000011010110",
9348 => "0000000011010110",
9349 => "0000000011010110",
9350 => "0000000011010110",
9351 => "0000000011010110",
9352 => "0000000011010110",
9353 => "0000000011010110",
9354 => "0000000011010111",
9355 => "0000000011010111",
9356 => "0000000011010111",
9357 => "0000000011010111",
9358 => "0000000011010111",
9359 => "0000000011010111",
9360 => "0000000011010111",
9361 => "0000000011010111",
9362 => "0000000011010111",
9363 => "0000000011010111",
9364 => "0000000011010111",
9365 => "0000000011010111",
9366 => "0000000011010111",
9367 => "0000000011010111",
9368 => "0000000011010111",
9369 => "0000000011010111",
9370 => "0000000011010111",
9371 => "0000000011010111",
9372 => "0000000011010111",
9373 => "0000000011011000",
9374 => "0000000011011000",
9375 => "0000000011011000",
9376 => "0000000011011000",
9377 => "0000000011011000",
9378 => "0000000011011000",
9379 => "0000000011011000",
9380 => "0000000011011000",
9381 => "0000000011011000",
9382 => "0000000011011000",
9383 => "0000000011011000",
9384 => "0000000011011000",
9385 => "0000000011011000",
9386 => "0000000011011000",
9387 => "0000000011011000",
9388 => "0000000011011000",
9389 => "0000000011011000",
9390 => "0000000011011000",
9391 => "0000000011011000",
9392 => "0000000011011001",
9393 => "0000000011011001",
9394 => "0000000011011001",
9395 => "0000000011011001",
9396 => "0000000011011001",
9397 => "0000000011011001",
9398 => "0000000011011001",
9399 => "0000000011011001",
9400 => "0000000011011001",
9401 => "0000000011011001",
9402 => "0000000011011001",
9403 => "0000000011011001",
9404 => "0000000011011001",
9405 => "0000000011011001",
9406 => "0000000011011001",
9407 => "0000000011011001",
9408 => "0000000011011001",
9409 => "0000000011011001",
9410 => "0000000011011001",
9411 => "0000000011011010",
9412 => "0000000011011010",
9413 => "0000000011011010",
9414 => "0000000011011010",
9415 => "0000000011011010",
9416 => "0000000011011010",
9417 => "0000000011011010",
9418 => "0000000011011010",
9419 => "0000000011011010",
9420 => "0000000011011010",
9421 => "0000000011011010",
9422 => "0000000011011010",
9423 => "0000000011011010",
9424 => "0000000011011010",
9425 => "0000000011011010",
9426 => "0000000011011010",
9427 => "0000000011011010",
9428 => "0000000011011010",
9429 => "0000000011011010",
9430 => "0000000011011011",
9431 => "0000000011011011",
9432 => "0000000011011011",
9433 => "0000000011011011",
9434 => "0000000011011011",
9435 => "0000000011011011",
9436 => "0000000011011011",
9437 => "0000000011011011",
9438 => "0000000011011011",
9439 => "0000000011011011",
9440 => "0000000011011011",
9441 => "0000000011011011",
9442 => "0000000011011011",
9443 => "0000000011011011",
9444 => "0000000011011011",
9445 => "0000000011011011",
9446 => "0000000011011011",
9447 => "0000000011011011",
9448 => "0000000011011100",
9449 => "0000000011011100",
9450 => "0000000011011100",
9451 => "0000000011011100",
9452 => "0000000011011100",
9453 => "0000000011011100",
9454 => "0000000011011100",
9455 => "0000000011011100",
9456 => "0000000011011100",
9457 => "0000000011011100",
9458 => "0000000011011100",
9459 => "0000000011011100",
9460 => "0000000011011100",
9461 => "0000000011011100",
9462 => "0000000011011100",
9463 => "0000000011011100",
9464 => "0000000011011100",
9465 => "0000000011011100",
9466 => "0000000011011100",
9467 => "0000000011011101",
9468 => "0000000011011101",
9469 => "0000000011011101",
9470 => "0000000011011101",
9471 => "0000000011011101",
9472 => "0000000011011101",
9473 => "0000000011011101",
9474 => "0000000011011101",
9475 => "0000000011011101",
9476 => "0000000011011101",
9477 => "0000000011011101",
9478 => "0000000011011101",
9479 => "0000000011011101",
9480 => "0000000011011101",
9481 => "0000000011011101",
9482 => "0000000011011101",
9483 => "0000000011011101",
9484 => "0000000011011101",
9485 => "0000000011011101",
9486 => "0000000011011110",
9487 => "0000000011011110",
9488 => "0000000011011110",
9489 => "0000000011011110",
9490 => "0000000011011110",
9491 => "0000000011011110",
9492 => "0000000011011110",
9493 => "0000000011011110",
9494 => "0000000011011110",
9495 => "0000000011011110",
9496 => "0000000011011110",
9497 => "0000000011011110",
9498 => "0000000011011110",
9499 => "0000000011011110",
9500 => "0000000011011110",
9501 => "0000000011011110",
9502 => "0000000011011110",
9503 => "0000000011011110",
9504 => "0000000011011111",
9505 => "0000000011011111",
9506 => "0000000011011111",
9507 => "0000000011011111",
9508 => "0000000011011111",
9509 => "0000000011011111",
9510 => "0000000011011111",
9511 => "0000000011011111",
9512 => "0000000011011111",
9513 => "0000000011011111",
9514 => "0000000011011111",
9515 => "0000000011011111",
9516 => "0000000011011111",
9517 => "0000000011011111",
9518 => "0000000011011111",
9519 => "0000000011011111",
9520 => "0000000011011111",
9521 => "0000000011011111",
9522 => "0000000011100000",
9523 => "0000000011100000",
9524 => "0000000011100000",
9525 => "0000000011100000",
9526 => "0000000011100000",
9527 => "0000000011100000",
9528 => "0000000011100000",
9529 => "0000000011100000",
9530 => "0000000011100000",
9531 => "0000000011100000",
9532 => "0000000011100000",
9533 => "0000000011100000",
9534 => "0000000011100000",
9535 => "0000000011100000",
9536 => "0000000011100000",
9537 => "0000000011100000",
9538 => "0000000011100000",
9539 => "0000000011100000",
9540 => "0000000011100000",
9541 => "0000000011100001",
9542 => "0000000011100001",
9543 => "0000000011100001",
9544 => "0000000011100001",
9545 => "0000000011100001",
9546 => "0000000011100001",
9547 => "0000000011100001",
9548 => "0000000011100001",
9549 => "0000000011100001",
9550 => "0000000011100001",
9551 => "0000000011100001",
9552 => "0000000011100001",
9553 => "0000000011100001",
9554 => "0000000011100001",
9555 => "0000000011100001",
9556 => "0000000011100001",
9557 => "0000000011100001",
9558 => "0000000011100001",
9559 => "0000000011100010",
9560 => "0000000011100010",
9561 => "0000000011100010",
9562 => "0000000011100010",
9563 => "0000000011100010",
9564 => "0000000011100010",
9565 => "0000000011100010",
9566 => "0000000011100010",
9567 => "0000000011100010",
9568 => "0000000011100010",
9569 => "0000000011100010",
9570 => "0000000011100010",
9571 => "0000000011100010",
9572 => "0000000011100010",
9573 => "0000000011100010",
9574 => "0000000011100010",
9575 => "0000000011100010",
9576 => "0000000011100010",
9577 => "0000000011100011",
9578 => "0000000011100011",
9579 => "0000000011100011",
9580 => "0000000011100011",
9581 => "0000000011100011",
9582 => "0000000011100011",
9583 => "0000000011100011",
9584 => "0000000011100011",
9585 => "0000000011100011",
9586 => "0000000011100011",
9587 => "0000000011100011",
9588 => "0000000011100011",
9589 => "0000000011100011",
9590 => "0000000011100011",
9591 => "0000000011100011",
9592 => "0000000011100011",
9593 => "0000000011100011",
9594 => "0000000011100011",
9595 => "0000000011100100",
9596 => "0000000011100100",
9597 => "0000000011100100",
9598 => "0000000011100100",
9599 => "0000000011100100",
9600 => "0000000011100100",
9601 => "0000000011100100",
9602 => "0000000011100100",
9603 => "0000000011100100",
9604 => "0000000011100100",
9605 => "0000000011100100",
9606 => "0000000011100100",
9607 => "0000000011100100",
9608 => "0000000011100100",
9609 => "0000000011100100",
9610 => "0000000011100100",
9611 => "0000000011100100",
9612 => "0000000011100100",
9613 => "0000000011100101",
9614 => "0000000011100101",
9615 => "0000000011100101",
9616 => "0000000011100101",
9617 => "0000000011100101",
9618 => "0000000011100101",
9619 => "0000000011100101",
9620 => "0000000011100101",
9621 => "0000000011100101",
9622 => "0000000011100101",
9623 => "0000000011100101",
9624 => "0000000011100101",
9625 => "0000000011100101",
9626 => "0000000011100101",
9627 => "0000000011100101",
9628 => "0000000011100101",
9629 => "0000000011100101",
9630 => "0000000011100101",
9631 => "0000000011100110",
9632 => "0000000011100110",
9633 => "0000000011100110",
9634 => "0000000011100110",
9635 => "0000000011100110",
9636 => "0000000011100110",
9637 => "0000000011100110",
9638 => "0000000011100110",
9639 => "0000000011100110",
9640 => "0000000011100110",
9641 => "0000000011100110",
9642 => "0000000011100110",
9643 => "0000000011100110",
9644 => "0000000011100110",
9645 => "0000000011100110",
9646 => "0000000011100110",
9647 => "0000000011100110",
9648 => "0000000011100110",
9649 => "0000000011100111",
9650 => "0000000011100111",
9651 => "0000000011100111",
9652 => "0000000011100111",
9653 => "0000000011100111",
9654 => "0000000011100111",
9655 => "0000000011100111",
9656 => "0000000011100111",
9657 => "0000000011100111",
9658 => "0000000011100111",
9659 => "0000000011100111",
9660 => "0000000011100111",
9661 => "0000000011100111",
9662 => "0000000011100111",
9663 => "0000000011100111",
9664 => "0000000011100111",
9665 => "0000000011100111",
9666 => "0000000011100111",
9667 => "0000000011101000",
9668 => "0000000011101000",
9669 => "0000000011101000",
9670 => "0000000011101000",
9671 => "0000000011101000",
9672 => "0000000011101000",
9673 => "0000000011101000",
9674 => "0000000011101000",
9675 => "0000000011101000",
9676 => "0000000011101000",
9677 => "0000000011101000",
9678 => "0000000011101000",
9679 => "0000000011101000",
9680 => "0000000011101000",
9681 => "0000000011101000",
9682 => "0000000011101000",
9683 => "0000000011101000",
9684 => "0000000011101001",
9685 => "0000000011101001",
9686 => "0000000011101001",
9687 => "0000000011101001",
9688 => "0000000011101001",
9689 => "0000000011101001",
9690 => "0000000011101001",
9691 => "0000000011101001",
9692 => "0000000011101001",
9693 => "0000000011101001",
9694 => "0000000011101001",
9695 => "0000000011101001",
9696 => "0000000011101001",
9697 => "0000000011101001",
9698 => "0000000011101001",
9699 => "0000000011101001",
9700 => "0000000011101001",
9701 => "0000000011101001",
9702 => "0000000011101010",
9703 => "0000000011101010",
9704 => "0000000011101010",
9705 => "0000000011101010",
9706 => "0000000011101010",
9707 => "0000000011101010",
9708 => "0000000011101010",
9709 => "0000000011101010",
9710 => "0000000011101010",
9711 => "0000000011101010",
9712 => "0000000011101010",
9713 => "0000000011101010",
9714 => "0000000011101010",
9715 => "0000000011101010",
9716 => "0000000011101010",
9717 => "0000000011101010",
9718 => "0000000011101010",
9719 => "0000000011101011",
9720 => "0000000011101011",
9721 => "0000000011101011",
9722 => "0000000011101011",
9723 => "0000000011101011",
9724 => "0000000011101011",
9725 => "0000000011101011",
9726 => "0000000011101011",
9727 => "0000000011101011",
9728 => "0000000011101011",
9729 => "0000000011101011",
9730 => "0000000011101011",
9731 => "0000000011101011",
9732 => "0000000011101011",
9733 => "0000000011101011",
9734 => "0000000011101011",
9735 => "0000000011101011",
9736 => "0000000011101011",
9737 => "0000000011101100",
9738 => "0000000011101100",
9739 => "0000000011101100",
9740 => "0000000011101100",
9741 => "0000000011101100",
9742 => "0000000011101100",
9743 => "0000000011101100",
9744 => "0000000011101100",
9745 => "0000000011101100",
9746 => "0000000011101100",
9747 => "0000000011101100",
9748 => "0000000011101100",
9749 => "0000000011101100",
9750 => "0000000011101100",
9751 => "0000000011101100",
9752 => "0000000011101100",
9753 => "0000000011101100",
9754 => "0000000011101101",
9755 => "0000000011101101",
9756 => "0000000011101101",
9757 => "0000000011101101",
9758 => "0000000011101101",
9759 => "0000000011101101",
9760 => "0000000011101101",
9761 => "0000000011101101",
9762 => "0000000011101101",
9763 => "0000000011101101",
9764 => "0000000011101101",
9765 => "0000000011101101",
9766 => "0000000011101101",
9767 => "0000000011101101",
9768 => "0000000011101101",
9769 => "0000000011101101",
9770 => "0000000011101101",
9771 => "0000000011101101",
9772 => "0000000011101110",
9773 => "0000000011101110",
9774 => "0000000011101110",
9775 => "0000000011101110",
9776 => "0000000011101110",
9777 => "0000000011101110",
9778 => "0000000011101110",
9779 => "0000000011101110",
9780 => "0000000011101110",
9781 => "0000000011101110",
9782 => "0000000011101110",
9783 => "0000000011101110",
9784 => "0000000011101110",
9785 => "0000000011101110",
9786 => "0000000011101110",
9787 => "0000000011101110",
9788 => "0000000011101110",
9789 => "0000000011101111",
9790 => "0000000011101111",
9791 => "0000000011101111",
9792 => "0000000011101111",
9793 => "0000000011101111",
9794 => "0000000011101111",
9795 => "0000000011101111",
9796 => "0000000011101111",
9797 => "0000000011101111",
9798 => "0000000011101111",
9799 => "0000000011101111",
9800 => "0000000011101111",
9801 => "0000000011101111",
9802 => "0000000011101111",
9803 => "0000000011101111",
9804 => "0000000011101111",
9805 => "0000000011101111",
9806 => "0000000011110000",
9807 => "0000000011110000",
9808 => "0000000011110000",
9809 => "0000000011110000",
9810 => "0000000011110000",
9811 => "0000000011110000",
9812 => "0000000011110000",
9813 => "0000000011110000",
9814 => "0000000011110000",
9815 => "0000000011110000",
9816 => "0000000011110000",
9817 => "0000000011110000",
9818 => "0000000011110000",
9819 => "0000000011110000",
9820 => "0000000011110000",
9821 => "0000000011110000",
9822 => "0000000011110000",
9823 => "0000000011110001",
9824 => "0000000011110001",
9825 => "0000000011110001",
9826 => "0000000011110001",
9827 => "0000000011110001",
9828 => "0000000011110001",
9829 => "0000000011110001",
9830 => "0000000011110001",
9831 => "0000000011110001",
9832 => "0000000011110001",
9833 => "0000000011110001",
9834 => "0000000011110001",
9835 => "0000000011110001",
9836 => "0000000011110001",
9837 => "0000000011110001",
9838 => "0000000011110001",
9839 => "0000000011110001",
9840 => "0000000011110010",
9841 => "0000000011110010",
9842 => "0000000011110010",
9843 => "0000000011110010",
9844 => "0000000011110010",
9845 => "0000000011110010",
9846 => "0000000011110010",
9847 => "0000000011110010",
9848 => "0000000011110010",
9849 => "0000000011110010",
9850 => "0000000011110010",
9851 => "0000000011110010",
9852 => "0000000011110010",
9853 => "0000000011110010",
9854 => "0000000011110010",
9855 => "0000000011110010",
9856 => "0000000011110010",
9857 => "0000000011110011",
9858 => "0000000011110011",
9859 => "0000000011110011",
9860 => "0000000011110011",
9861 => "0000000011110011",
9862 => "0000000011110011",
9863 => "0000000011110011",
9864 => "0000000011110011",
9865 => "0000000011110011",
9866 => "0000000011110011",
9867 => "0000000011110011",
9868 => "0000000011110011",
9869 => "0000000011110011",
9870 => "0000000011110011",
9871 => "0000000011110011",
9872 => "0000000011110011",
9873 => "0000000011110011",
9874 => "0000000011110100",
9875 => "0000000011110100",
9876 => "0000000011110100",
9877 => "0000000011110100",
9878 => "0000000011110100",
9879 => "0000000011110100",
9880 => "0000000011110100",
9881 => "0000000011110100",
9882 => "0000000011110100",
9883 => "0000000011110100",
9884 => "0000000011110100",
9885 => "0000000011110100",
9886 => "0000000011110100",
9887 => "0000000011110100",
9888 => "0000000011110100",
9889 => "0000000011110100",
9890 => "0000000011110100",
9891 => "0000000011110101",
9892 => "0000000011110101",
9893 => "0000000011110101",
9894 => "0000000011110101",
9895 => "0000000011110101",
9896 => "0000000011110101",
9897 => "0000000011110101",
9898 => "0000000011110101",
9899 => "0000000011110101",
9900 => "0000000011110101",
9901 => "0000000011110101",
9902 => "0000000011110101",
9903 => "0000000011110101",
9904 => "0000000011110101",
9905 => "0000000011110101",
9906 => "0000000011110101",
9907 => "0000000011110110",
9908 => "0000000011110110",
9909 => "0000000011110110",
9910 => "0000000011110110",
9911 => "0000000011110110",
9912 => "0000000011110110",
9913 => "0000000011110110",
9914 => "0000000011110110",
9915 => "0000000011110110",
9916 => "0000000011110110",
9917 => "0000000011110110",
9918 => "0000000011110110",
9919 => "0000000011110110",
9920 => "0000000011110110",
9921 => "0000000011110110",
9922 => "0000000011110110",
9923 => "0000000011110110",
9924 => "0000000011110111",
9925 => "0000000011110111",
9926 => "0000000011110111",
9927 => "0000000011110111",
9928 => "0000000011110111",
9929 => "0000000011110111",
9930 => "0000000011110111",
9931 => "0000000011110111",
9932 => "0000000011110111",
9933 => "0000000011110111",
9934 => "0000000011110111",
9935 => "0000000011110111",
9936 => "0000000011110111",
9937 => "0000000011110111",
9938 => "0000000011110111",
9939 => "0000000011110111",
9940 => "0000000011110111",
9941 => "0000000011111000",
9942 => "0000000011111000",
9943 => "0000000011111000",
9944 => "0000000011111000",
9945 => "0000000011111000",
9946 => "0000000011111000",
9947 => "0000000011111000",
9948 => "0000000011111000",
9949 => "0000000011111000",
9950 => "0000000011111000",
9951 => "0000000011111000",
9952 => "0000000011111000",
9953 => "0000000011111000",
9954 => "0000000011111000",
9955 => "0000000011111000",
9956 => "0000000011111000",
9957 => "0000000011111001",
9958 => "0000000011111001",
9959 => "0000000011111001",
9960 => "0000000011111001",
9961 => "0000000011111001",
9962 => "0000000011111001",
9963 => "0000000011111001",
9964 => "0000000011111001",
9965 => "0000000011111001",
9966 => "0000000011111001",
9967 => "0000000011111001",
9968 => "0000000011111001",
9969 => "0000000011111001",
9970 => "0000000011111001",
9971 => "0000000011111001",
9972 => "0000000011111001",
9973 => "0000000011111001",
9974 => "0000000011111010",
9975 => "0000000011111010",
9976 => "0000000011111010",
9977 => "0000000011111010",
9978 => "0000000011111010",
9979 => "0000000011111010",
9980 => "0000000011111010",
9981 => "0000000011111010",
9982 => "0000000011111010",
9983 => "0000000011111010",
9984 => "0000000011111010",
9985 => "0000000011111010",
9986 => "0000000011111010",
9987 => "0000000011111010",
9988 => "0000000011111010",
9989 => "0000000011111010",
9990 => "0000000011111011",
9991 => "0000000011111011",
9992 => "0000000011111011",
9993 => "0000000011111011",
9994 => "0000000011111011",
9995 => "0000000011111011",
9996 => "0000000011111011",
9997 => "0000000011111011",
9998 => "0000000011111011",
9999 => "0000000011111011",
10000 => "0000000011111011",
10001 => "0000000011111011",
10002 => "0000000011111011",
10003 => "0000000011111011",
10004 => "0000000011111011",
10005 => "0000000011111011",
10006 => "0000000011111011",
10007 => "0000000011111100",
10008 => "0000000011111100",
10009 => "0000000011111100",
10010 => "0000000011111100",
10011 => "0000000011111100",
10012 => "0000000011111100",
10013 => "0000000011111100",
10014 => "0000000011111100",
10015 => "0000000011111100",
10016 => "0000000011111100",
10017 => "0000000011111100",
10018 => "0000000011111100",
10019 => "0000000011111100",
10020 => "0000000011111100",
10021 => "0000000011111100",
10022 => "0000000011111100",
10023 => "0000000011111101",
10024 => "0000000011111101",
10025 => "0000000011111101",
10026 => "0000000011111101",
10027 => "0000000011111101",
10028 => "0000000011111101",
10029 => "0000000011111101",
10030 => "0000000011111101",
10031 => "0000000011111101",
10032 => "0000000011111101",
10033 => "0000000011111101",
10034 => "0000000011111101",
10035 => "0000000011111101",
10036 => "0000000011111101",
10037 => "0000000011111101",
10038 => "0000000011111101",
10039 => "0000000011111110",
10040 => "0000000011111110",
10041 => "0000000011111110",
10042 => "0000000011111110",
10043 => "0000000011111110",
10044 => "0000000011111110",
10045 => "0000000011111110",
10046 => "0000000011111110",
10047 => "0000000011111110",
10048 => "0000000011111110",
10049 => "0000000011111110",
10050 => "0000000011111110",
10051 => "0000000011111110",
10052 => "0000000011111110",
10053 => "0000000011111110",
10054 => "0000000011111110",
10055 => "0000000011111111",
10056 => "0000000011111111",
10057 => "0000000011111111",
10058 => "0000000011111111",
10059 => "0000000011111111",
10060 => "0000000011111111",
10061 => "0000000011111111",
10062 => "0000000011111111",
10063 => "0000000011111111",
10064 => "0000000011111111",
10065 => "0000000011111111",
10066 => "0000000011111111",
10067 => "0000000011111111",
10068 => "0000000011111111",
10069 => "0000000011111111",
10070 => "0000000011111111",
10071 => "0000000100000000",
10072 => "0000000100000000",
10073 => "0000000100000000",
10074 => "0000000100000000",
10075 => "0000000100000000",
10076 => "0000000100000000",
10077 => "0000000100000000",
10078 => "0000000100000000",
10079 => "0000000100000000",
10080 => "0000000100000000",
10081 => "0000000100000000",
10082 => "0000000100000000",
10083 => "0000000100000000",
10084 => "0000000100000000",
10085 => "0000000100000000",
10086 => "0000000100000000",
10087 => "0000000100000001",
10088 => "0000000100000001",
10089 => "0000000100000001",
10090 => "0000000100000001",
10091 => "0000000100000001",
10092 => "0000000100000001",
10093 => "0000000100000001",
10094 => "0000000100000001",
10095 => "0000000100000001",
10096 => "0000000100000001",
10097 => "0000000100000001",
10098 => "0000000100000001",
10099 => "0000000100000001",
10100 => "0000000100000001",
10101 => "0000000100000001",
10102 => "0000000100000001",
10103 => "0000000100000010",
10104 => "0000000100000010",
10105 => "0000000100000010",
10106 => "0000000100000010",
10107 => "0000000100000010",
10108 => "0000000100000010",
10109 => "0000000100000010",
10110 => "0000000100000010",
10111 => "0000000100000010",
10112 => "0000000100000010",
10113 => "0000000100000010",
10114 => "0000000100000010",
10115 => "0000000100000010",
10116 => "0000000100000010",
10117 => "0000000100000010",
10118 => "0000000100000010",
10119 => "0000000100000011",
10120 => "0000000100000011",
10121 => "0000000100000011",
10122 => "0000000100000011",
10123 => "0000000100000011",
10124 => "0000000100000011",
10125 => "0000000100000011",
10126 => "0000000100000011",
10127 => "0000000100000011",
10128 => "0000000100000011",
10129 => "0000000100000011",
10130 => "0000000100000011",
10131 => "0000000100000011",
10132 => "0000000100000011",
10133 => "0000000100000011",
10134 => "0000000100000011",
10135 => "0000000100000100",
10136 => "0000000100000100",
10137 => "0000000100000100",
10138 => "0000000100000100",
10139 => "0000000100000100",
10140 => "0000000100000100",
10141 => "0000000100000100",
10142 => "0000000100000100",
10143 => "0000000100000100",
10144 => "0000000100000100",
10145 => "0000000100000100",
10146 => "0000000100000100",
10147 => "0000000100000100",
10148 => "0000000100000100",
10149 => "0000000100000100",
10150 => "0000000100000100",
10151 => "0000000100000101",
10152 => "0000000100000101",
10153 => "0000000100000101",
10154 => "0000000100000101",
10155 => "0000000100000101",
10156 => "0000000100000101",
10157 => "0000000100000101",
10158 => "0000000100000101",
10159 => "0000000100000101",
10160 => "0000000100000101",
10161 => "0000000100000101",
10162 => "0000000100000101",
10163 => "0000000100000101",
10164 => "0000000100000101",
10165 => "0000000100000101",
10166 => "0000000100000101",
10167 => "0000000100000110",
10168 => "0000000100000110",
10169 => "0000000100000110",
10170 => "0000000100000110",
10171 => "0000000100000110",
10172 => "0000000100000110",
10173 => "0000000100000110",
10174 => "0000000100000110",
10175 => "0000000100000110",
10176 => "0000000100000110",
10177 => "0000000100000110",
10178 => "0000000100000110",
10179 => "0000000100000110",
10180 => "0000000100000110",
10181 => "0000000100000110",
10182 => "0000000100000111",
10183 => "0000000100000111",
10184 => "0000000100000111",
10185 => "0000000100000111",
10186 => "0000000100000111",
10187 => "0000000100000111",
10188 => "0000000100000111",
10189 => "0000000100000111",
10190 => "0000000100000111",
10191 => "0000000100000111",
10192 => "0000000100000111",
10193 => "0000000100000111",
10194 => "0000000100000111",
10195 => "0000000100000111",
10196 => "0000000100000111",
10197 => "0000000100000111",
10198 => "0000000100001000",
10199 => "0000000100001000",
10200 => "0000000100001000",
10201 => "0000000100001000",
10202 => "0000000100001000",
10203 => "0000000100001000",
10204 => "0000000100001000",
10205 => "0000000100001000",
10206 => "0000000100001000",
10207 => "0000000100001000",
10208 => "0000000100001000",
10209 => "0000000100001000",
10210 => "0000000100001000",
10211 => "0000000100001000",
10212 => "0000000100001000",
10213 => "0000000100001001",
10214 => "0000000100001001",
10215 => "0000000100001001",
10216 => "0000000100001001",
10217 => "0000000100001001",
10218 => "0000000100001001",
10219 => "0000000100001001",
10220 => "0000000100001001",
10221 => "0000000100001001",
10222 => "0000000100001001",
10223 => "0000000100001001",
10224 => "0000000100001001",
10225 => "0000000100001001",
10226 => "0000000100001001",
10227 => "0000000100001001",
10228 => "0000000100001001",
10229 => "0000000100001010",
10230 => "0000000100001010",
10231 => "0000000100001010",
10232 => "0000000100001010",
10233 => "0000000100001010",
10234 => "0000000100001010",
10235 => "0000000100001010",
10236 => "0000000100001010",
10237 => "0000000100001010",
10238 => "0000000100001010",
10239 => "0000000100001010",
10240 => "0000000100001010",
10241 => "0000000100001010",
10242 => "0000000100001010",
10243 => "0000000100001010",
10244 => "0000000100001011",
10245 => "0000000100001011",
10246 => "0000000100001011",
10247 => "0000000100001011",
10248 => "0000000100001011",
10249 => "0000000100001011",
10250 => "0000000100001011",
10251 => "0000000100001011",
10252 => "0000000100001011",
10253 => "0000000100001011",
10254 => "0000000100001011",
10255 => "0000000100001011",
10256 => "0000000100001011",
10257 => "0000000100001011",
10258 => "0000000100001011",
10259 => "0000000100001011",
10260 => "0000000100001100",
10261 => "0000000100001100",
10262 => "0000000100001100",
10263 => "0000000100001100",
10264 => "0000000100001100",
10265 => "0000000100001100",
10266 => "0000000100001100",
10267 => "0000000100001100",
10268 => "0000000100001100",
10269 => "0000000100001100",
10270 => "0000000100001100",
10271 => "0000000100001100",
10272 => "0000000100001100",
10273 => "0000000100001100",
10274 => "0000000100001100",
10275 => "0000000100001101",
10276 => "0000000100001101",
10277 => "0000000100001101",
10278 => "0000000100001101",
10279 => "0000000100001101",
10280 => "0000000100001101",
10281 => "0000000100001101",
10282 => "0000000100001101",
10283 => "0000000100001101",
10284 => "0000000100001101",
10285 => "0000000100001101",
10286 => "0000000100001101",
10287 => "0000000100001101",
10288 => "0000000100001101",
10289 => "0000000100001101",
10290 => "0000000100001110",
10291 => "0000000100001110",
10292 => "0000000100001110",
10293 => "0000000100001110",
10294 => "0000000100001110",
10295 => "0000000100001110",
10296 => "0000000100001110",
10297 => "0000000100001110",
10298 => "0000000100001110",
10299 => "0000000100001110",
10300 => "0000000100001110",
10301 => "0000000100001110",
10302 => "0000000100001110",
10303 => "0000000100001110",
10304 => "0000000100001110",
10305 => "0000000100001110",
10306 => "0000000100001111",
10307 => "0000000100001111",
10308 => "0000000100001111",
10309 => "0000000100001111",
10310 => "0000000100001111",
10311 => "0000000100001111",
10312 => "0000000100001111",
10313 => "0000000100001111",
10314 => "0000000100001111",
10315 => "0000000100001111",
10316 => "0000000100001111",
10317 => "0000000100001111",
10318 => "0000000100001111",
10319 => "0000000100001111",
10320 => "0000000100001111",
10321 => "0000000100010000",
10322 => "0000000100010000",
10323 => "0000000100010000",
10324 => "0000000100010000",
10325 => "0000000100010000",
10326 => "0000000100010000",
10327 => "0000000100010000",
10328 => "0000000100010000",
10329 => "0000000100010000",
10330 => "0000000100010000",
10331 => "0000000100010000",
10332 => "0000000100010000",
10333 => "0000000100010000",
10334 => "0000000100010000",
10335 => "0000000100010000",
10336 => "0000000100010001",
10337 => "0000000100010001",
10338 => "0000000100010001",
10339 => "0000000100010001",
10340 => "0000000100010001",
10341 => "0000000100010001",
10342 => "0000000100010001",
10343 => "0000000100010001",
10344 => "0000000100010001",
10345 => "0000000100010001",
10346 => "0000000100010001",
10347 => "0000000100010001",
10348 => "0000000100010001",
10349 => "0000000100010001",
10350 => "0000000100010001",
10351 => "0000000100010010",
10352 => "0000000100010010",
10353 => "0000000100010010",
10354 => "0000000100010010",
10355 => "0000000100010010",
10356 => "0000000100010010",
10357 => "0000000100010010",
10358 => "0000000100010010",
10359 => "0000000100010010",
10360 => "0000000100010010",
10361 => "0000000100010010",
10362 => "0000000100010010",
10363 => "0000000100010010",
10364 => "0000000100010010",
10365 => "0000000100010010",
10366 => "0000000100010011",
10367 => "0000000100010011",
10368 => "0000000100010011",
10369 => "0000000100010011",
10370 => "0000000100010011",
10371 => "0000000100010011",
10372 => "0000000100010011",
10373 => "0000000100010011",
10374 => "0000000100010011",
10375 => "0000000100010011",
10376 => "0000000100010011",
10377 => "0000000100010011",
10378 => "0000000100010011",
10379 => "0000000100010011",
10380 => "0000000100010011",
10381 => "0000000100010100",
10382 => "0000000100010100",
10383 => "0000000100010100",
10384 => "0000000100010100",
10385 => "0000000100010100",
10386 => "0000000100010100",
10387 => "0000000100010100",
10388 => "0000000100010100",
10389 => "0000000100010100",
10390 => "0000000100010100",
10391 => "0000000100010100",
10392 => "0000000100010100",
10393 => "0000000100010100",
10394 => "0000000100010100",
10395 => "0000000100010100",
10396 => "0000000100010101",
10397 => "0000000100010101",
10398 => "0000000100010101",
10399 => "0000000100010101",
10400 => "0000000100010101",
10401 => "0000000100010101",
10402 => "0000000100010101",
10403 => "0000000100010101",
10404 => "0000000100010101",
10405 => "0000000100010101",
10406 => "0000000100010101",
10407 => "0000000100010101",
10408 => "0000000100010101",
10409 => "0000000100010101",
10410 => "0000000100010110",
10411 => "0000000100010110",
10412 => "0000000100010110",
10413 => "0000000100010110",
10414 => "0000000100010110",
10415 => "0000000100010110",
10416 => "0000000100010110",
10417 => "0000000100010110",
10418 => "0000000100010110",
10419 => "0000000100010110",
10420 => "0000000100010110",
10421 => "0000000100010110",
10422 => "0000000100010110",
10423 => "0000000100010110",
10424 => "0000000100010110",
10425 => "0000000100010111",
10426 => "0000000100010111",
10427 => "0000000100010111",
10428 => "0000000100010111",
10429 => "0000000100010111",
10430 => "0000000100010111",
10431 => "0000000100010111",
10432 => "0000000100010111",
10433 => "0000000100010111",
10434 => "0000000100010111",
10435 => "0000000100010111",
10436 => "0000000100010111",
10437 => "0000000100010111",
10438 => "0000000100010111",
10439 => "0000000100010111",
10440 => "0000000100011000",
10441 => "0000000100011000",
10442 => "0000000100011000",
10443 => "0000000100011000",
10444 => "0000000100011000",
10445 => "0000000100011000",
10446 => "0000000100011000",
10447 => "0000000100011000",
10448 => "0000000100011000",
10449 => "0000000100011000",
10450 => "0000000100011000",
10451 => "0000000100011000",
10452 => "0000000100011000",
10453 => "0000000100011000",
10454 => "0000000100011000",
10455 => "0000000100011001",
10456 => "0000000100011001",
10457 => "0000000100011001",
10458 => "0000000100011001",
10459 => "0000000100011001",
10460 => "0000000100011001",
10461 => "0000000100011001",
10462 => "0000000100011001",
10463 => "0000000100011001",
10464 => "0000000100011001",
10465 => "0000000100011001",
10466 => "0000000100011001",
10467 => "0000000100011001",
10468 => "0000000100011001",
10469 => "0000000100011010",
10470 => "0000000100011010",
10471 => "0000000100011010",
10472 => "0000000100011010",
10473 => "0000000100011010",
10474 => "0000000100011010",
10475 => "0000000100011010",
10476 => "0000000100011010",
10477 => "0000000100011010",
10478 => "0000000100011010",
10479 => "0000000100011010",
10480 => "0000000100011010",
10481 => "0000000100011010",
10482 => "0000000100011010",
10483 => "0000000100011010",
10484 => "0000000100011011",
10485 => "0000000100011011",
10486 => "0000000100011011",
10487 => "0000000100011011",
10488 => "0000000100011011",
10489 => "0000000100011011",
10490 => "0000000100011011",
10491 => "0000000100011011",
10492 => "0000000100011011",
10493 => "0000000100011011",
10494 => "0000000100011011",
10495 => "0000000100011011",
10496 => "0000000100011011",
10497 => "0000000100011011",
10498 => "0000000100011100",
10499 => "0000000100011100",
10500 => "0000000100011100",
10501 => "0000000100011100",
10502 => "0000000100011100",
10503 => "0000000100011100",
10504 => "0000000100011100",
10505 => "0000000100011100",
10506 => "0000000100011100",
10507 => "0000000100011100",
10508 => "0000000100011100",
10509 => "0000000100011100",
10510 => "0000000100011100",
10511 => "0000000100011100",
10512 => "0000000100011100",
10513 => "0000000100011101",
10514 => "0000000100011101",
10515 => "0000000100011101",
10516 => "0000000100011101",
10517 => "0000000100011101",
10518 => "0000000100011101",
10519 => "0000000100011101",
10520 => "0000000100011101",
10521 => "0000000100011101",
10522 => "0000000100011101",
10523 => "0000000100011101",
10524 => "0000000100011101",
10525 => "0000000100011101",
10526 => "0000000100011101",
10527 => "0000000100011110",
10528 => "0000000100011110",
10529 => "0000000100011110",
10530 => "0000000100011110",
10531 => "0000000100011110",
10532 => "0000000100011110",
10533 => "0000000100011110",
10534 => "0000000100011110",
10535 => "0000000100011110",
10536 => "0000000100011110",
10537 => "0000000100011110",
10538 => "0000000100011110",
10539 => "0000000100011110",
10540 => "0000000100011110",
10541 => "0000000100011111",
10542 => "0000000100011111",
10543 => "0000000100011111",
10544 => "0000000100011111",
10545 => "0000000100011111",
10546 => "0000000100011111",
10547 => "0000000100011111",
10548 => "0000000100011111",
10549 => "0000000100011111",
10550 => "0000000100011111",
10551 => "0000000100011111",
10552 => "0000000100011111",
10553 => "0000000100011111",
10554 => "0000000100011111",
10555 => "0000000100011111",
10556 => "0000000100100000",
10557 => "0000000100100000",
10558 => "0000000100100000",
10559 => "0000000100100000",
10560 => "0000000100100000",
10561 => "0000000100100000",
10562 => "0000000100100000",
10563 => "0000000100100000",
10564 => "0000000100100000",
10565 => "0000000100100000",
10566 => "0000000100100000",
10567 => "0000000100100000",
10568 => "0000000100100000",
10569 => "0000000100100000",
10570 => "0000000100100001",
10571 => "0000000100100001",
10572 => "0000000100100001",
10573 => "0000000100100001",
10574 => "0000000100100001",
10575 => "0000000100100001",
10576 => "0000000100100001",
10577 => "0000000100100001",
10578 => "0000000100100001",
10579 => "0000000100100001",
10580 => "0000000100100001",
10581 => "0000000100100001",
10582 => "0000000100100001",
10583 => "0000000100100001",
10584 => "0000000100100010",
10585 => "0000000100100010",
10586 => "0000000100100010",
10587 => "0000000100100010",
10588 => "0000000100100010",
10589 => "0000000100100010",
10590 => "0000000100100010",
10591 => "0000000100100010",
10592 => "0000000100100010",
10593 => "0000000100100010",
10594 => "0000000100100010",
10595 => "0000000100100010",
10596 => "0000000100100010",
10597 => "0000000100100010",
10598 => "0000000100100011",
10599 => "0000000100100011",
10600 => "0000000100100011",
10601 => "0000000100100011",
10602 => "0000000100100011",
10603 => "0000000100100011",
10604 => "0000000100100011",
10605 => "0000000100100011",
10606 => "0000000100100011",
10607 => "0000000100100011",
10608 => "0000000100100011",
10609 => "0000000100100011",
10610 => "0000000100100011",
10611 => "0000000100100011",
10612 => "0000000100100011",
10613 => "0000000100100100",
10614 => "0000000100100100",
10615 => "0000000100100100",
10616 => "0000000100100100",
10617 => "0000000100100100",
10618 => "0000000100100100",
10619 => "0000000100100100",
10620 => "0000000100100100",
10621 => "0000000100100100",
10622 => "0000000100100100",
10623 => "0000000100100100",
10624 => "0000000100100100",
10625 => "0000000100100100",
10626 => "0000000100100100",
10627 => "0000000100100101",
10628 => "0000000100100101",
10629 => "0000000100100101",
10630 => "0000000100100101",
10631 => "0000000100100101",
10632 => "0000000100100101",
10633 => "0000000100100101",
10634 => "0000000100100101",
10635 => "0000000100100101",
10636 => "0000000100100101",
10637 => "0000000100100101",
10638 => "0000000100100101",
10639 => "0000000100100101",
10640 => "0000000100100101",
10641 => "0000000100100110",
10642 => "0000000100100110",
10643 => "0000000100100110",
10644 => "0000000100100110",
10645 => "0000000100100110",
10646 => "0000000100100110",
10647 => "0000000100100110",
10648 => "0000000100100110",
10649 => "0000000100100110",
10650 => "0000000100100110",
10651 => "0000000100100110",
10652 => "0000000100100110",
10653 => "0000000100100110",
10654 => "0000000100100110",
10655 => "0000000100100111",
10656 => "0000000100100111",
10657 => "0000000100100111",
10658 => "0000000100100111",
10659 => "0000000100100111",
10660 => "0000000100100111",
10661 => "0000000100100111",
10662 => "0000000100100111",
10663 => "0000000100100111",
10664 => "0000000100100111",
10665 => "0000000100100111",
10666 => "0000000100100111",
10667 => "0000000100100111",
10668 => "0000000100101000",
10669 => "0000000100101000",
10670 => "0000000100101000",
10671 => "0000000100101000",
10672 => "0000000100101000",
10673 => "0000000100101000",
10674 => "0000000100101000",
10675 => "0000000100101000",
10676 => "0000000100101000",
10677 => "0000000100101000",
10678 => "0000000100101000",
10679 => "0000000100101000",
10680 => "0000000100101000",
10681 => "0000000100101000",
10682 => "0000000100101001",
10683 => "0000000100101001",
10684 => "0000000100101001",
10685 => "0000000100101001",
10686 => "0000000100101001",
10687 => "0000000100101001",
10688 => "0000000100101001",
10689 => "0000000100101001",
10690 => "0000000100101001",
10691 => "0000000100101001",
10692 => "0000000100101001",
10693 => "0000000100101001",
10694 => "0000000100101001",
10695 => "0000000100101001",
10696 => "0000000100101010",
10697 => "0000000100101010",
10698 => "0000000100101010",
10699 => "0000000100101010",
10700 => "0000000100101010",
10701 => "0000000100101010",
10702 => "0000000100101010",
10703 => "0000000100101010",
10704 => "0000000100101010",
10705 => "0000000100101010",
10706 => "0000000100101010",
10707 => "0000000100101010",
10708 => "0000000100101010",
10709 => "0000000100101010",
10710 => "0000000100101011",
10711 => "0000000100101011",
10712 => "0000000100101011",
10713 => "0000000100101011",
10714 => "0000000100101011",
10715 => "0000000100101011",
10716 => "0000000100101011",
10717 => "0000000100101011",
10718 => "0000000100101011",
10719 => "0000000100101011",
10720 => "0000000100101011",
10721 => "0000000100101011",
10722 => "0000000100101011",
10723 => "0000000100101011",
10724 => "0000000100101100",
10725 => "0000000100101100",
10726 => "0000000100101100",
10727 => "0000000100101100",
10728 => "0000000100101100",
10729 => "0000000100101100",
10730 => "0000000100101100",
10731 => "0000000100101100",
10732 => "0000000100101100",
10733 => "0000000100101100",
10734 => "0000000100101100",
10735 => "0000000100101100",
10736 => "0000000100101100",
10737 => "0000000100101101",
10738 => "0000000100101101",
10739 => "0000000100101101",
10740 => "0000000100101101",
10741 => "0000000100101101",
10742 => "0000000100101101",
10743 => "0000000100101101",
10744 => "0000000100101101",
10745 => "0000000100101101",
10746 => "0000000100101101",
10747 => "0000000100101101",
10748 => "0000000100101101",
10749 => "0000000100101101",
10750 => "0000000100101101",
10751 => "0000000100101110",
10752 => "0000000100101110",
10753 => "0000000100101110",
10754 => "0000000100101110",
10755 => "0000000100101110",
10756 => "0000000100101110",
10757 => "0000000100101110",
10758 => "0000000100101110",
10759 => "0000000100101110",
10760 => "0000000100101110",
10761 => "0000000100101110",
10762 => "0000000100101110",
10763 => "0000000100101110",
10764 => "0000000100101110",
10765 => "0000000100101111",
10766 => "0000000100101111",
10767 => "0000000100101111",
10768 => "0000000100101111",
10769 => "0000000100101111",
10770 => "0000000100101111",
10771 => "0000000100101111",
10772 => "0000000100101111",
10773 => "0000000100101111",
10774 => "0000000100101111",
10775 => "0000000100101111",
10776 => "0000000100101111",
10777 => "0000000100101111",
10778 => "0000000100110000",
10779 => "0000000100110000",
10780 => "0000000100110000",
10781 => "0000000100110000",
10782 => "0000000100110000",
10783 => "0000000100110000",
10784 => "0000000100110000",
10785 => "0000000100110000",
10786 => "0000000100110000",
10787 => "0000000100110000",
10788 => "0000000100110000",
10789 => "0000000100110000",
10790 => "0000000100110000",
10791 => "0000000100110000",
10792 => "0000000100110001",
10793 => "0000000100110001",
10794 => "0000000100110001",
10795 => "0000000100110001",
10796 => "0000000100110001",
10797 => "0000000100110001",
10798 => "0000000100110001",
10799 => "0000000100110001",
10800 => "0000000100110001",
10801 => "0000000100110001",
10802 => "0000000100110001",
10803 => "0000000100110001",
10804 => "0000000100110001",
10805 => "0000000100110010",
10806 => "0000000100110010",
10807 => "0000000100110010",
10808 => "0000000100110010",
10809 => "0000000100110010",
10810 => "0000000100110010",
10811 => "0000000100110010",
10812 => "0000000100110010",
10813 => "0000000100110010",
10814 => "0000000100110010",
10815 => "0000000100110010",
10816 => "0000000100110010",
10817 => "0000000100110010",
10818 => "0000000100110010",
10819 => "0000000100110011",
10820 => "0000000100110011",
10821 => "0000000100110011",
10822 => "0000000100110011",
10823 => "0000000100110011",
10824 => "0000000100110011",
10825 => "0000000100110011",
10826 => "0000000100110011",
10827 => "0000000100110011",
10828 => "0000000100110011",
10829 => "0000000100110011",
10830 => "0000000100110011",
10831 => "0000000100110011",
10832 => "0000000100110100",
10833 => "0000000100110100",
10834 => "0000000100110100",
10835 => "0000000100110100",
10836 => "0000000100110100",
10837 => "0000000100110100",
10838 => "0000000100110100",
10839 => "0000000100110100",
10840 => "0000000100110100",
10841 => "0000000100110100",
10842 => "0000000100110100",
10843 => "0000000100110100",
10844 => "0000000100110100",
10845 => "0000000100110101",
10846 => "0000000100110101",
10847 => "0000000100110101",
10848 => "0000000100110101",
10849 => "0000000100110101",
10850 => "0000000100110101",
10851 => "0000000100110101",
10852 => "0000000100110101",
10853 => "0000000100110101",
10854 => "0000000100110101",
10855 => "0000000100110101",
10856 => "0000000100110101",
10857 => "0000000100110101",
10858 => "0000000100110101",
10859 => "0000000100110110",
10860 => "0000000100110110",
10861 => "0000000100110110",
10862 => "0000000100110110",
10863 => "0000000100110110",
10864 => "0000000100110110",
10865 => "0000000100110110",
10866 => "0000000100110110",
10867 => "0000000100110110",
10868 => "0000000100110110",
10869 => "0000000100110110",
10870 => "0000000100110110",
10871 => "0000000100110110",
10872 => "0000000100110111",
10873 => "0000000100110111",
10874 => "0000000100110111",
10875 => "0000000100110111",
10876 => "0000000100110111",
10877 => "0000000100110111",
10878 => "0000000100110111",
10879 => "0000000100110111",
10880 => "0000000100110111",
10881 => "0000000100110111",
10882 => "0000000100110111",
10883 => "0000000100110111",
10884 => "0000000100110111",
10885 => "0000000100111000",
10886 => "0000000100111000",
10887 => "0000000100111000",
10888 => "0000000100111000",
10889 => "0000000100111000",
10890 => "0000000100111000",
10891 => "0000000100111000",
10892 => "0000000100111000",
10893 => "0000000100111000",
10894 => "0000000100111000",
10895 => "0000000100111000",
10896 => "0000000100111000",
10897 => "0000000100111000",
10898 => "0000000100111001",
10899 => "0000000100111001",
10900 => "0000000100111001",
10901 => "0000000100111001",
10902 => "0000000100111001",
10903 => "0000000100111001",
10904 => "0000000100111001",
10905 => "0000000100111001",
10906 => "0000000100111001",
10907 => "0000000100111001",
10908 => "0000000100111001",
10909 => "0000000100111001",
10910 => "0000000100111001",
10911 => "0000000100111010",
10912 => "0000000100111010",
10913 => "0000000100111010",
10914 => "0000000100111010",
10915 => "0000000100111010",
10916 => "0000000100111010",
10917 => "0000000100111010",
10918 => "0000000100111010",
10919 => "0000000100111010",
10920 => "0000000100111010",
10921 => "0000000100111010",
10922 => "0000000100111010",
10923 => "0000000100111010",
10924 => "0000000100111010",
10925 => "0000000100111011",
10926 => "0000000100111011",
10927 => "0000000100111011",
10928 => "0000000100111011",
10929 => "0000000100111011",
10930 => "0000000100111011",
10931 => "0000000100111011",
10932 => "0000000100111011",
10933 => "0000000100111011",
10934 => "0000000100111011",
10935 => "0000000100111011",
10936 => "0000000100111011",
10937 => "0000000100111011",
10938 => "0000000100111100",
10939 => "0000000100111100",
10940 => "0000000100111100",
10941 => "0000000100111100",
10942 => "0000000100111100",
10943 => "0000000100111100",
10944 => "0000000100111100",
10945 => "0000000100111100",
10946 => "0000000100111100",
10947 => "0000000100111100",
10948 => "0000000100111100",
10949 => "0000000100111100",
10950 => "0000000100111100",
10951 => "0000000100111101",
10952 => "0000000100111101",
10953 => "0000000100111101",
10954 => "0000000100111101",
10955 => "0000000100111101",
10956 => "0000000100111101",
10957 => "0000000100111101",
10958 => "0000000100111101",
10959 => "0000000100111101",
10960 => "0000000100111101",
10961 => "0000000100111101",
10962 => "0000000100111101",
10963 => "0000000100111101",
10964 => "0000000100111110",
10965 => "0000000100111110",
10966 => "0000000100111110",
10967 => "0000000100111110",
10968 => "0000000100111110",
10969 => "0000000100111110",
10970 => "0000000100111110",
10971 => "0000000100111110",
10972 => "0000000100111110",
10973 => "0000000100111110",
10974 => "0000000100111110",
10975 => "0000000100111110",
10976 => "0000000100111111",
10977 => "0000000100111111",
10978 => "0000000100111111",
10979 => "0000000100111111",
10980 => "0000000100111111",
10981 => "0000000100111111",
10982 => "0000000100111111",
10983 => "0000000100111111",
10984 => "0000000100111111",
10985 => "0000000100111111",
10986 => "0000000100111111",
10987 => "0000000100111111",
10988 => "0000000100111111",
10989 => "0000000101000000",
10990 => "0000000101000000",
10991 => "0000000101000000",
10992 => "0000000101000000",
10993 => "0000000101000000",
10994 => "0000000101000000",
10995 => "0000000101000000",
10996 => "0000000101000000",
10997 => "0000000101000000",
10998 => "0000000101000000",
10999 => "0000000101000000",
11000 => "0000000101000000",
11001 => "0000000101000000",
11002 => "0000000101000001",
11003 => "0000000101000001",
11004 => "0000000101000001",
11005 => "0000000101000001",
11006 => "0000000101000001",
11007 => "0000000101000001",
11008 => "0000000101000001",
11009 => "0000000101000001",
11010 => "0000000101000001",
11011 => "0000000101000001",
11012 => "0000000101000001",
11013 => "0000000101000001",
11014 => "0000000101000001",
11015 => "0000000101000010",
11016 => "0000000101000010",
11017 => "0000000101000010",
11018 => "0000000101000010",
11019 => "0000000101000010",
11020 => "0000000101000010",
11021 => "0000000101000010",
11022 => "0000000101000010",
11023 => "0000000101000010",
11024 => "0000000101000010",
11025 => "0000000101000010",
11026 => "0000000101000010",
11027 => "0000000101000010",
11028 => "0000000101000011",
11029 => "0000000101000011",
11030 => "0000000101000011",
11031 => "0000000101000011",
11032 => "0000000101000011",
11033 => "0000000101000011",
11034 => "0000000101000011",
11035 => "0000000101000011",
11036 => "0000000101000011",
11037 => "0000000101000011",
11038 => "0000000101000011",
11039 => "0000000101000011",
11040 => "0000000101000100",
11041 => "0000000101000100",
11042 => "0000000101000100",
11043 => "0000000101000100",
11044 => "0000000101000100",
11045 => "0000000101000100",
11046 => "0000000101000100",
11047 => "0000000101000100",
11048 => "0000000101000100",
11049 => "0000000101000100",
11050 => "0000000101000100",
11051 => "0000000101000100",
11052 => "0000000101000100",
11053 => "0000000101000101",
11054 => "0000000101000101",
11055 => "0000000101000101",
11056 => "0000000101000101",
11057 => "0000000101000101",
11058 => "0000000101000101",
11059 => "0000000101000101",
11060 => "0000000101000101",
11061 => "0000000101000101",
11062 => "0000000101000101",
11063 => "0000000101000101",
11064 => "0000000101000101",
11065 => "0000000101000101",
11066 => "0000000101000110",
11067 => "0000000101000110",
11068 => "0000000101000110",
11069 => "0000000101000110",
11070 => "0000000101000110",
11071 => "0000000101000110",
11072 => "0000000101000110",
11073 => "0000000101000110",
11074 => "0000000101000110",
11075 => "0000000101000110",
11076 => "0000000101000110",
11077 => "0000000101000110",
11078 => "0000000101000111",
11079 => "0000000101000111",
11080 => "0000000101000111",
11081 => "0000000101000111",
11082 => "0000000101000111",
11083 => "0000000101000111",
11084 => "0000000101000111",
11085 => "0000000101000111",
11086 => "0000000101000111",
11087 => "0000000101000111",
11088 => "0000000101000111",
11089 => "0000000101000111",
11090 => "0000000101000111",
11091 => "0000000101001000",
11092 => "0000000101001000",
11093 => "0000000101001000",
11094 => "0000000101001000",
11095 => "0000000101001000",
11096 => "0000000101001000",
11097 => "0000000101001000",
11098 => "0000000101001000",
11099 => "0000000101001000",
11100 => "0000000101001000",
11101 => "0000000101001000",
11102 => "0000000101001000",
11103 => "0000000101001000",
11104 => "0000000101001001",
11105 => "0000000101001001",
11106 => "0000000101001001",
11107 => "0000000101001001",
11108 => "0000000101001001",
11109 => "0000000101001001",
11110 => "0000000101001001",
11111 => "0000000101001001",
11112 => "0000000101001001",
11113 => "0000000101001001",
11114 => "0000000101001001",
11115 => "0000000101001001",
11116 => "0000000101001010",
11117 => "0000000101001010",
11118 => "0000000101001010",
11119 => "0000000101001010",
11120 => "0000000101001010",
11121 => "0000000101001010",
11122 => "0000000101001010",
11123 => "0000000101001010",
11124 => "0000000101001010",
11125 => "0000000101001010",
11126 => "0000000101001010",
11127 => "0000000101001010",
11128 => "0000000101001011",
11129 => "0000000101001011",
11130 => "0000000101001011",
11131 => "0000000101001011",
11132 => "0000000101001011",
11133 => "0000000101001011",
11134 => "0000000101001011",
11135 => "0000000101001011",
11136 => "0000000101001011",
11137 => "0000000101001011",
11138 => "0000000101001011",
11139 => "0000000101001011",
11140 => "0000000101001011",
11141 => "0000000101001100",
11142 => "0000000101001100",
11143 => "0000000101001100",
11144 => "0000000101001100",
11145 => "0000000101001100",
11146 => "0000000101001100",
11147 => "0000000101001100",
11148 => "0000000101001100",
11149 => "0000000101001100",
11150 => "0000000101001100",
11151 => "0000000101001100",
11152 => "0000000101001100",
11153 => "0000000101001101",
11154 => "0000000101001101",
11155 => "0000000101001101",
11156 => "0000000101001101",
11157 => "0000000101001101",
11158 => "0000000101001101",
11159 => "0000000101001101",
11160 => "0000000101001101",
11161 => "0000000101001101",
11162 => "0000000101001101",
11163 => "0000000101001101",
11164 => "0000000101001101",
11165 => "0000000101001101",
11166 => "0000000101001110",
11167 => "0000000101001110",
11168 => "0000000101001110",
11169 => "0000000101001110",
11170 => "0000000101001110",
11171 => "0000000101001110",
11172 => "0000000101001110",
11173 => "0000000101001110",
11174 => "0000000101001110",
11175 => "0000000101001110",
11176 => "0000000101001110",
11177 => "0000000101001110",
11178 => "0000000101001111",
11179 => "0000000101001111",
11180 => "0000000101001111",
11181 => "0000000101001111",
11182 => "0000000101001111",
11183 => "0000000101001111",
11184 => "0000000101001111",
11185 => "0000000101001111",
11186 => "0000000101001111",
11187 => "0000000101001111",
11188 => "0000000101001111",
11189 => "0000000101001111",
11190 => "0000000101010000",
11191 => "0000000101010000",
11192 => "0000000101010000",
11193 => "0000000101010000",
11194 => "0000000101010000",
11195 => "0000000101010000",
11196 => "0000000101010000",
11197 => "0000000101010000",
11198 => "0000000101010000",
11199 => "0000000101010000",
11200 => "0000000101010000",
11201 => "0000000101010000",
11202 => "0000000101010001",
11203 => "0000000101010001",
11204 => "0000000101010001",
11205 => "0000000101010001",
11206 => "0000000101010001",
11207 => "0000000101010001",
11208 => "0000000101010001",
11209 => "0000000101010001",
11210 => "0000000101010001",
11211 => "0000000101010001",
11212 => "0000000101010001",
11213 => "0000000101010001",
11214 => "0000000101010001",
11215 => "0000000101010010",
11216 => "0000000101010010",
11217 => "0000000101010010",
11218 => "0000000101010010",
11219 => "0000000101010010",
11220 => "0000000101010010",
11221 => "0000000101010010",
11222 => "0000000101010010",
11223 => "0000000101010010",
11224 => "0000000101010010",
11225 => "0000000101010010",
11226 => "0000000101010010",
11227 => "0000000101010011",
11228 => "0000000101010011",
11229 => "0000000101010011",
11230 => "0000000101010011",
11231 => "0000000101010011",
11232 => "0000000101010011",
11233 => "0000000101010011",
11234 => "0000000101010011",
11235 => "0000000101010011",
11236 => "0000000101010011",
11237 => "0000000101010011",
11238 => "0000000101010011",
11239 => "0000000101010100",
11240 => "0000000101010100",
11241 => "0000000101010100",
11242 => "0000000101010100",
11243 => "0000000101010100",
11244 => "0000000101010100",
11245 => "0000000101010100",
11246 => "0000000101010100",
11247 => "0000000101010100",
11248 => "0000000101010100",
11249 => "0000000101010100",
11250 => "0000000101010100",
11251 => "0000000101010101",
11252 => "0000000101010101",
11253 => "0000000101010101",
11254 => "0000000101010101",
11255 => "0000000101010101",
11256 => "0000000101010101",
11257 => "0000000101010101",
11258 => "0000000101010101",
11259 => "0000000101010101",
11260 => "0000000101010101",
11261 => "0000000101010101",
11262 => "0000000101010101",
11263 => "0000000101010110",
11264 => "0000000101010110",
11265 => "0000000101010110",
11266 => "0000000101010110",
11267 => "0000000101010110",
11268 => "0000000101010110",
11269 => "0000000101010110",
11270 => "0000000101010110",
11271 => "0000000101010110",
11272 => "0000000101010110",
11273 => "0000000101010110",
11274 => "0000000101010110",
11275 => "0000000101010111",
11276 => "0000000101010111",
11277 => "0000000101010111",
11278 => "0000000101010111",
11279 => "0000000101010111",
11280 => "0000000101010111",
11281 => "0000000101010111",
11282 => "0000000101010111",
11283 => "0000000101010111",
11284 => "0000000101010111",
11285 => "0000000101010111",
11286 => "0000000101010111",
11287 => "0000000101011000",
11288 => "0000000101011000",
11289 => "0000000101011000",
11290 => "0000000101011000",
11291 => "0000000101011000",
11292 => "0000000101011000",
11293 => "0000000101011000",
11294 => "0000000101011000",
11295 => "0000000101011000",
11296 => "0000000101011000",
11297 => "0000000101011000",
11298 => "0000000101011000",
11299 => "0000000101011001",
11300 => "0000000101011001",
11301 => "0000000101011001",
11302 => "0000000101011001",
11303 => "0000000101011001",
11304 => "0000000101011001",
11305 => "0000000101011001",
11306 => "0000000101011001",
11307 => "0000000101011001",
11308 => "0000000101011001",
11309 => "0000000101011001",
11310 => "0000000101011001",
11311 => "0000000101011010",
11312 => "0000000101011010",
11313 => "0000000101011010",
11314 => "0000000101011010",
11315 => "0000000101011010",
11316 => "0000000101011010",
11317 => "0000000101011010",
11318 => "0000000101011010",
11319 => "0000000101011010",
11320 => "0000000101011010",
11321 => "0000000101011010",
11322 => "0000000101011010",
11323 => "0000000101011011",
11324 => "0000000101011011",
11325 => "0000000101011011",
11326 => "0000000101011011",
11327 => "0000000101011011",
11328 => "0000000101011011",
11329 => "0000000101011011",
11330 => "0000000101011011",
11331 => "0000000101011011",
11332 => "0000000101011011",
11333 => "0000000101011011",
11334 => "0000000101011011",
11335 => "0000000101011100",
11336 => "0000000101011100",
11337 => "0000000101011100",
11338 => "0000000101011100",
11339 => "0000000101011100",
11340 => "0000000101011100",
11341 => "0000000101011100",
11342 => "0000000101011100",
11343 => "0000000101011100",
11344 => "0000000101011100",
11345 => "0000000101011100",
11346 => "0000000101011101",
11347 => "0000000101011101",
11348 => "0000000101011101",
11349 => "0000000101011101",
11350 => "0000000101011101",
11351 => "0000000101011101",
11352 => "0000000101011101",
11353 => "0000000101011101",
11354 => "0000000101011101",
11355 => "0000000101011101",
11356 => "0000000101011101",
11357 => "0000000101011101",
11358 => "0000000101011110",
11359 => "0000000101011110",
11360 => "0000000101011110",
11361 => "0000000101011110",
11362 => "0000000101011110",
11363 => "0000000101011110",
11364 => "0000000101011110",
11365 => "0000000101011110",
11366 => "0000000101011110",
11367 => "0000000101011110",
11368 => "0000000101011110",
11369 => "0000000101011110",
11370 => "0000000101011111",
11371 => "0000000101011111",
11372 => "0000000101011111",
11373 => "0000000101011111",
11374 => "0000000101011111",
11375 => "0000000101011111",
11376 => "0000000101011111",
11377 => "0000000101011111",
11378 => "0000000101011111",
11379 => "0000000101011111",
11380 => "0000000101011111",
11381 => "0000000101011111",
11382 => "0000000101100000",
11383 => "0000000101100000",
11384 => "0000000101100000",
11385 => "0000000101100000",
11386 => "0000000101100000",
11387 => "0000000101100000",
11388 => "0000000101100000",
11389 => "0000000101100000",
11390 => "0000000101100000",
11391 => "0000000101100000",
11392 => "0000000101100000",
11393 => "0000000101100001",
11394 => "0000000101100001",
11395 => "0000000101100001",
11396 => "0000000101100001",
11397 => "0000000101100001",
11398 => "0000000101100001",
11399 => "0000000101100001",
11400 => "0000000101100001",
11401 => "0000000101100001",
11402 => "0000000101100001",
11403 => "0000000101100001",
11404 => "0000000101100001",
11405 => "0000000101100010",
11406 => "0000000101100010",
11407 => "0000000101100010",
11408 => "0000000101100010",
11409 => "0000000101100010",
11410 => "0000000101100010",
11411 => "0000000101100010",
11412 => "0000000101100010",
11413 => "0000000101100010",
11414 => "0000000101100010",
11415 => "0000000101100010",
11416 => "0000000101100010",
11417 => "0000000101100011",
11418 => "0000000101100011",
11419 => "0000000101100011",
11420 => "0000000101100011",
11421 => "0000000101100011",
11422 => "0000000101100011",
11423 => "0000000101100011",
11424 => "0000000101100011",
11425 => "0000000101100011",
11426 => "0000000101100011",
11427 => "0000000101100011",
11428 => "0000000101100100",
11429 => "0000000101100100",
11430 => "0000000101100100",
11431 => "0000000101100100",
11432 => "0000000101100100",
11433 => "0000000101100100",
11434 => "0000000101100100",
11435 => "0000000101100100",
11436 => "0000000101100100",
11437 => "0000000101100100",
11438 => "0000000101100100",
11439 => "0000000101100100",
11440 => "0000000101100101",
11441 => "0000000101100101",
11442 => "0000000101100101",
11443 => "0000000101100101",
11444 => "0000000101100101",
11445 => "0000000101100101",
11446 => "0000000101100101",
11447 => "0000000101100101",
11448 => "0000000101100101",
11449 => "0000000101100101",
11450 => "0000000101100101",
11451 => "0000000101100110",
11452 => "0000000101100110",
11453 => "0000000101100110",
11454 => "0000000101100110",
11455 => "0000000101100110",
11456 => "0000000101100110",
11457 => "0000000101100110",
11458 => "0000000101100110",
11459 => "0000000101100110",
11460 => "0000000101100110",
11461 => "0000000101100110",
11462 => "0000000101100110",
11463 => "0000000101100111",
11464 => "0000000101100111",
11465 => "0000000101100111",
11466 => "0000000101100111",
11467 => "0000000101100111",
11468 => "0000000101100111",
11469 => "0000000101100111",
11470 => "0000000101100111",
11471 => "0000000101100111",
11472 => "0000000101100111",
11473 => "0000000101100111",
11474 => "0000000101101000",
11475 => "0000000101101000",
11476 => "0000000101101000",
11477 => "0000000101101000",
11478 => "0000000101101000",
11479 => "0000000101101000",
11480 => "0000000101101000",
11481 => "0000000101101000",
11482 => "0000000101101000",
11483 => "0000000101101000",
11484 => "0000000101101000",
11485 => "0000000101101000",
11486 => "0000000101101001",
11487 => "0000000101101001",
11488 => "0000000101101001",
11489 => "0000000101101001",
11490 => "0000000101101001",
11491 => "0000000101101001",
11492 => "0000000101101001",
11493 => "0000000101101001",
11494 => "0000000101101001",
11495 => "0000000101101001",
11496 => "0000000101101001",
11497 => "0000000101101010",
11498 => "0000000101101010",
11499 => "0000000101101010",
11500 => "0000000101101010",
11501 => "0000000101101010",
11502 => "0000000101101010",
11503 => "0000000101101010",
11504 => "0000000101101010",
11505 => "0000000101101010",
11506 => "0000000101101010",
11507 => "0000000101101010",
11508 => "0000000101101011",
11509 => "0000000101101011",
11510 => "0000000101101011",
11511 => "0000000101101011",
11512 => "0000000101101011",
11513 => "0000000101101011",
11514 => "0000000101101011",
11515 => "0000000101101011",
11516 => "0000000101101011",
11517 => "0000000101101011",
11518 => "0000000101101011",
11519 => "0000000101101011",
11520 => "0000000101101100",
11521 => "0000000101101100",
11522 => "0000000101101100",
11523 => "0000000101101100",
11524 => "0000000101101100",
11525 => "0000000101101100",
11526 => "0000000101101100",
11527 => "0000000101101100",
11528 => "0000000101101100",
11529 => "0000000101101100",
11530 => "0000000101101100",
11531 => "0000000101101101",
11532 => "0000000101101101",
11533 => "0000000101101101",
11534 => "0000000101101101",
11535 => "0000000101101101",
11536 => "0000000101101101",
11537 => "0000000101101101",
11538 => "0000000101101101",
11539 => "0000000101101101",
11540 => "0000000101101101",
11541 => "0000000101101101",
11542 => "0000000101101110",
11543 => "0000000101101110",
11544 => "0000000101101110",
11545 => "0000000101101110",
11546 => "0000000101101110",
11547 => "0000000101101110",
11548 => "0000000101101110",
11549 => "0000000101101110",
11550 => "0000000101101110",
11551 => "0000000101101110",
11552 => "0000000101101110",
11553 => "0000000101101110",
11554 => "0000000101101111",
11555 => "0000000101101111",
11556 => "0000000101101111",
11557 => "0000000101101111",
11558 => "0000000101101111",
11559 => "0000000101101111",
11560 => "0000000101101111",
11561 => "0000000101101111",
11562 => "0000000101101111",
11563 => "0000000101101111",
11564 => "0000000101101111",
11565 => "0000000101110000",
11566 => "0000000101110000",
11567 => "0000000101110000",
11568 => "0000000101110000",
11569 => "0000000101110000",
11570 => "0000000101110000",
11571 => "0000000101110000",
11572 => "0000000101110000",
11573 => "0000000101110000",
11574 => "0000000101110000",
11575 => "0000000101110000",
11576 => "0000000101110001",
11577 => "0000000101110001",
11578 => "0000000101110001",
11579 => "0000000101110001",
11580 => "0000000101110001",
11581 => "0000000101110001",
11582 => "0000000101110001",
11583 => "0000000101110001",
11584 => "0000000101110001",
11585 => "0000000101110001",
11586 => "0000000101110001",
11587 => "0000000101110010",
11588 => "0000000101110010",
11589 => "0000000101110010",
11590 => "0000000101110010",
11591 => "0000000101110010",
11592 => "0000000101110010",
11593 => "0000000101110010",
11594 => "0000000101110010",
11595 => "0000000101110010",
11596 => "0000000101110010",
11597 => "0000000101110010",
11598 => "0000000101110011",
11599 => "0000000101110011",
11600 => "0000000101110011",
11601 => "0000000101110011",
11602 => "0000000101110011",
11603 => "0000000101110011",
11604 => "0000000101110011",
11605 => "0000000101110011",
11606 => "0000000101110011",
11607 => "0000000101110011",
11608 => "0000000101110011",
11609 => "0000000101110100",
11610 => "0000000101110100",
11611 => "0000000101110100",
11612 => "0000000101110100",
11613 => "0000000101110100",
11614 => "0000000101110100",
11615 => "0000000101110100",
11616 => "0000000101110100",
11617 => "0000000101110100",
11618 => "0000000101110100",
11619 => "0000000101110100",
11620 => "0000000101110101",
11621 => "0000000101110101",
11622 => "0000000101110101",
11623 => "0000000101110101",
11624 => "0000000101110101",
11625 => "0000000101110101",
11626 => "0000000101110101",
11627 => "0000000101110101",
11628 => "0000000101110101",
11629 => "0000000101110101",
11630 => "0000000101110101",
11631 => "0000000101110110",
11632 => "0000000101110110",
11633 => "0000000101110110",
11634 => "0000000101110110",
11635 => "0000000101110110",
11636 => "0000000101110110",
11637 => "0000000101110110",
11638 => "0000000101110110",
11639 => "0000000101110110",
11640 => "0000000101110110",
11641 => "0000000101110110",
11642 => "0000000101110111",
11643 => "0000000101110111",
11644 => "0000000101110111",
11645 => "0000000101110111",
11646 => "0000000101110111",
11647 => "0000000101110111",
11648 => "0000000101110111",
11649 => "0000000101110111",
11650 => "0000000101110111",
11651 => "0000000101110111",
11652 => "0000000101110111",
11653 => "0000000101111000",
11654 => "0000000101111000",
11655 => "0000000101111000",
11656 => "0000000101111000",
11657 => "0000000101111000",
11658 => "0000000101111000",
11659 => "0000000101111000",
11660 => "0000000101111000",
11661 => "0000000101111000",
11662 => "0000000101111000",
11663 => "0000000101111000",
11664 => "0000000101111001",
11665 => "0000000101111001",
11666 => "0000000101111001",
11667 => "0000000101111001",
11668 => "0000000101111001",
11669 => "0000000101111001",
11670 => "0000000101111001",
11671 => "0000000101111001",
11672 => "0000000101111001",
11673 => "0000000101111001",
11674 => "0000000101111001",
11675 => "0000000101111010",
11676 => "0000000101111010",
11677 => "0000000101111010",
11678 => "0000000101111010",
11679 => "0000000101111010",
11680 => "0000000101111010",
11681 => "0000000101111010",
11682 => "0000000101111010",
11683 => "0000000101111010",
11684 => "0000000101111010",
11685 => "0000000101111010",
11686 => "0000000101111011",
11687 => "0000000101111011",
11688 => "0000000101111011",
11689 => "0000000101111011",
11690 => "0000000101111011",
11691 => "0000000101111011",
11692 => "0000000101111011",
11693 => "0000000101111011",
11694 => "0000000101111011",
11695 => "0000000101111011",
11696 => "0000000101111011",
11697 => "0000000101111100",
11698 => "0000000101111100",
11699 => "0000000101111100",
11700 => "0000000101111100",
11701 => "0000000101111100",
11702 => "0000000101111100",
11703 => "0000000101111100",
11704 => "0000000101111100",
11705 => "0000000101111100",
11706 => "0000000101111100",
11707 => "0000000101111100",
11708 => "0000000101111101",
11709 => "0000000101111101",
11710 => "0000000101111101",
11711 => "0000000101111101",
11712 => "0000000101111101",
11713 => "0000000101111101",
11714 => "0000000101111101",
11715 => "0000000101111101",
11716 => "0000000101111101",
11717 => "0000000101111101",
11718 => "0000000101111101",
11719 => "0000000101111110",
11720 => "0000000101111110",
11721 => "0000000101111110",
11722 => "0000000101111110",
11723 => "0000000101111110",
11724 => "0000000101111110",
11725 => "0000000101111110",
11726 => "0000000101111110",
11727 => "0000000101111110",
11728 => "0000000101111110",
11729 => "0000000101111111",
11730 => "0000000101111111",
11731 => "0000000101111111",
11732 => "0000000101111111",
11733 => "0000000101111111",
11734 => "0000000101111111",
11735 => "0000000101111111",
11736 => "0000000101111111",
11737 => "0000000101111111",
11738 => "0000000101111111",
11739 => "0000000101111111",
11740 => "0000000110000000",
11741 => "0000000110000000",
11742 => "0000000110000000",
11743 => "0000000110000000",
11744 => "0000000110000000",
11745 => "0000000110000000",
11746 => "0000000110000000",
11747 => "0000000110000000",
11748 => "0000000110000000",
11749 => "0000000110000000",
11750 => "0000000110000000",
11751 => "0000000110000001",
11752 => "0000000110000001",
11753 => "0000000110000001",
11754 => "0000000110000001",
11755 => "0000000110000001",
11756 => "0000000110000001",
11757 => "0000000110000001",
11758 => "0000000110000001",
11759 => "0000000110000001",
11760 => "0000000110000001",
11761 => "0000000110000001",
11762 => "0000000110000010",
11763 => "0000000110000010",
11764 => "0000000110000010",
11765 => "0000000110000010",
11766 => "0000000110000010",
11767 => "0000000110000010",
11768 => "0000000110000010",
11769 => "0000000110000010",
11770 => "0000000110000010",
11771 => "0000000110000010",
11772 => "0000000110000011",
11773 => "0000000110000011",
11774 => "0000000110000011",
11775 => "0000000110000011",
11776 => "0000000110000011",
11777 => "0000000110000011",
11778 => "0000000110000011",
11779 => "0000000110000011",
11780 => "0000000110000011",
11781 => "0000000110000011",
11782 => "0000000110000011",
11783 => "0000000110000100",
11784 => "0000000110000100",
11785 => "0000000110000100",
11786 => "0000000110000100",
11787 => "0000000110000100",
11788 => "0000000110000100",
11789 => "0000000110000100",
11790 => "0000000110000100",
11791 => "0000000110000100",
11792 => "0000000110000100",
11793 => "0000000110000101",
11794 => "0000000110000101",
11795 => "0000000110000101",
11796 => "0000000110000101",
11797 => "0000000110000101",
11798 => "0000000110000101",
11799 => "0000000110000101",
11800 => "0000000110000101",
11801 => "0000000110000101",
11802 => "0000000110000101",
11803 => "0000000110000101",
11804 => "0000000110000110",
11805 => "0000000110000110",
11806 => "0000000110000110",
11807 => "0000000110000110",
11808 => "0000000110000110",
11809 => "0000000110000110",
11810 => "0000000110000110",
11811 => "0000000110000110",
11812 => "0000000110000110",
11813 => "0000000110000110",
11814 => "0000000110000110",
11815 => "0000000110000111",
11816 => "0000000110000111",
11817 => "0000000110000111",
11818 => "0000000110000111",
11819 => "0000000110000111",
11820 => "0000000110000111",
11821 => "0000000110000111",
11822 => "0000000110000111",
11823 => "0000000110000111",
11824 => "0000000110000111",
11825 => "0000000110001000",
11826 => "0000000110001000",
11827 => "0000000110001000",
11828 => "0000000110001000",
11829 => "0000000110001000",
11830 => "0000000110001000",
11831 => "0000000110001000",
11832 => "0000000110001000",
11833 => "0000000110001000",
11834 => "0000000110001000",
11835 => "0000000110001000",
11836 => "0000000110001001",
11837 => "0000000110001001",
11838 => "0000000110001001",
11839 => "0000000110001001",
11840 => "0000000110001001",
11841 => "0000000110001001",
11842 => "0000000110001001",
11843 => "0000000110001001",
11844 => "0000000110001001",
11845 => "0000000110001001",
11846 => "0000000110001010",
11847 => "0000000110001010",
11848 => "0000000110001010",
11849 => "0000000110001010",
11850 => "0000000110001010",
11851 => "0000000110001010",
11852 => "0000000110001010",
11853 => "0000000110001010",
11854 => "0000000110001010",
11855 => "0000000110001010",
11856 => "0000000110001010",
11857 => "0000000110001011",
11858 => "0000000110001011",
11859 => "0000000110001011",
11860 => "0000000110001011",
11861 => "0000000110001011",
11862 => "0000000110001011",
11863 => "0000000110001011",
11864 => "0000000110001011",
11865 => "0000000110001011",
11866 => "0000000110001011",
11867 => "0000000110001100",
11868 => "0000000110001100",
11869 => "0000000110001100",
11870 => "0000000110001100",
11871 => "0000000110001100",
11872 => "0000000110001100",
11873 => "0000000110001100",
11874 => "0000000110001100",
11875 => "0000000110001100",
11876 => "0000000110001100",
11877 => "0000000110001101",
11878 => "0000000110001101",
11879 => "0000000110001101",
11880 => "0000000110001101",
11881 => "0000000110001101",
11882 => "0000000110001101",
11883 => "0000000110001101",
11884 => "0000000110001101",
11885 => "0000000110001101",
11886 => "0000000110001101",
11887 => "0000000110001101",
11888 => "0000000110001110",
11889 => "0000000110001110",
11890 => "0000000110001110",
11891 => "0000000110001110",
11892 => "0000000110001110",
11893 => "0000000110001110",
11894 => "0000000110001110",
11895 => "0000000110001110",
11896 => "0000000110001110",
11897 => "0000000110001110",
11898 => "0000000110001111",
11899 => "0000000110001111",
11900 => "0000000110001111",
11901 => "0000000110001111",
11902 => "0000000110001111",
11903 => "0000000110001111",
11904 => "0000000110001111",
11905 => "0000000110001111",
11906 => "0000000110001111",
11907 => "0000000110001111",
11908 => "0000000110010000",
11909 => "0000000110010000",
11910 => "0000000110010000",
11911 => "0000000110010000",
11912 => "0000000110010000",
11913 => "0000000110010000",
11914 => "0000000110010000",
11915 => "0000000110010000",
11916 => "0000000110010000",
11917 => "0000000110010000",
11918 => "0000000110010000",
11919 => "0000000110010001",
11920 => "0000000110010001",
11921 => "0000000110010001",
11922 => "0000000110010001",
11923 => "0000000110010001",
11924 => "0000000110010001",
11925 => "0000000110010001",
11926 => "0000000110010001",
11927 => "0000000110010001",
11928 => "0000000110010001",
11929 => "0000000110010010",
11930 => "0000000110010010",
11931 => "0000000110010010",
11932 => "0000000110010010",
11933 => "0000000110010010",
11934 => "0000000110010010",
11935 => "0000000110010010",
11936 => "0000000110010010",
11937 => "0000000110010010",
11938 => "0000000110010010",
11939 => "0000000110010011",
11940 => "0000000110010011",
11941 => "0000000110010011",
11942 => "0000000110010011",
11943 => "0000000110010011",
11944 => "0000000110010011",
11945 => "0000000110010011",
11946 => "0000000110010011",
11947 => "0000000110010011",
11948 => "0000000110010011",
11949 => "0000000110010100",
11950 => "0000000110010100",
11951 => "0000000110010100",
11952 => "0000000110010100",
11953 => "0000000110010100",
11954 => "0000000110010100",
11955 => "0000000110010100",
11956 => "0000000110010100",
11957 => "0000000110010100",
11958 => "0000000110010100",
11959 => "0000000110010100",
11960 => "0000000110010101",
11961 => "0000000110010101",
11962 => "0000000110010101",
11963 => "0000000110010101",
11964 => "0000000110010101",
11965 => "0000000110010101",
11966 => "0000000110010101",
11967 => "0000000110010101",
11968 => "0000000110010101",
11969 => "0000000110010101",
11970 => "0000000110010110",
11971 => "0000000110010110",
11972 => "0000000110010110",
11973 => "0000000110010110",
11974 => "0000000110010110",
11975 => "0000000110010110",
11976 => "0000000110010110",
11977 => "0000000110010110",
11978 => "0000000110010110",
11979 => "0000000110010110",
11980 => "0000000110010111",
11981 => "0000000110010111",
11982 => "0000000110010111",
11983 => "0000000110010111",
11984 => "0000000110010111",
11985 => "0000000110010111",
11986 => "0000000110010111",
11987 => "0000000110010111",
11988 => "0000000110010111",
11989 => "0000000110010111",
11990 => "0000000110011000",
11991 => "0000000110011000",
11992 => "0000000110011000",
11993 => "0000000110011000",
11994 => "0000000110011000",
11995 => "0000000110011000",
11996 => "0000000110011000",
11997 => "0000000110011000",
11998 => "0000000110011000",
11999 => "0000000110011000",
12000 => "0000000110011001",
12001 => "0000000110011001",
12002 => "0000000110011001",
12003 => "0000000110011001",
12004 => "0000000110011001",
12005 => "0000000110011001",
12006 => "0000000110011001",
12007 => "0000000110011001",
12008 => "0000000110011001",
12009 => "0000000110011001",
12010 => "0000000110011010",
12011 => "0000000110011010",
12012 => "0000000110011010",
12013 => "0000000110011010",
12014 => "0000000110011010",
12015 => "0000000110011010",
12016 => "0000000110011010",
12017 => "0000000110011010",
12018 => "0000000110011010",
12019 => "0000000110011010",
12020 => "0000000110011011",
12021 => "0000000110011011",
12022 => "0000000110011011",
12023 => "0000000110011011",
12024 => "0000000110011011",
12025 => "0000000110011011",
12026 => "0000000110011011",
12027 => "0000000110011011",
12028 => "0000000110011011",
12029 => "0000000110011011",
12030 => "0000000110011100",
12031 => "0000000110011100",
12032 => "0000000110011100",
12033 => "0000000110011100",
12034 => "0000000110011100",
12035 => "0000000110011100",
12036 => "0000000110011100",
12037 => "0000000110011100",
12038 => "0000000110011100",
12039 => "0000000110011100",
12040 => "0000000110011101",
12041 => "0000000110011101",
12042 => "0000000110011101",
12043 => "0000000110011101",
12044 => "0000000110011101",
12045 => "0000000110011101",
12046 => "0000000110011101",
12047 => "0000000110011101",
12048 => "0000000110011101",
12049 => "0000000110011101",
12050 => "0000000110011110",
12051 => "0000000110011110",
12052 => "0000000110011110",
12053 => "0000000110011110",
12054 => "0000000110011110",
12055 => "0000000110011110",
12056 => "0000000110011110",
12057 => "0000000110011110",
12058 => "0000000110011110",
12059 => "0000000110011110",
12060 => "0000000110011111",
12061 => "0000000110011111",
12062 => "0000000110011111",
12063 => "0000000110011111",
12064 => "0000000110011111",
12065 => "0000000110011111",
12066 => "0000000110011111",
12067 => "0000000110011111",
12068 => "0000000110011111",
12069 => "0000000110011111",
12070 => "0000000110100000",
12071 => "0000000110100000",
12072 => "0000000110100000",
12073 => "0000000110100000",
12074 => "0000000110100000",
12075 => "0000000110100000",
12076 => "0000000110100000",
12077 => "0000000110100000",
12078 => "0000000110100000",
12079 => "0000000110100000",
12080 => "0000000110100001",
12081 => "0000000110100001",
12082 => "0000000110100001",
12083 => "0000000110100001",
12084 => "0000000110100001",
12085 => "0000000110100001",
12086 => "0000000110100001",
12087 => "0000000110100001",
12088 => "0000000110100001",
12089 => "0000000110100001",
12090 => "0000000110100010",
12091 => "0000000110100010",
12092 => "0000000110100010",
12093 => "0000000110100010",
12094 => "0000000110100010",
12095 => "0000000110100010",
12096 => "0000000110100010",
12097 => "0000000110100010",
12098 => "0000000110100010",
12099 => "0000000110100010",
12100 => "0000000110100011",
12101 => "0000000110100011",
12102 => "0000000110100011",
12103 => "0000000110100011",
12104 => "0000000110100011",
12105 => "0000000110100011",
12106 => "0000000110100011",
12107 => "0000000110100011",
12108 => "0000000110100011",
12109 => "0000000110100100",
12110 => "0000000110100100",
12111 => "0000000110100100",
12112 => "0000000110100100",
12113 => "0000000110100100",
12114 => "0000000110100100",
12115 => "0000000110100100",
12116 => "0000000110100100",
12117 => "0000000110100100",
12118 => "0000000110100100",
12119 => "0000000110100101",
12120 => "0000000110100101",
12121 => "0000000110100101",
12122 => "0000000110100101",
12123 => "0000000110100101",
12124 => "0000000110100101",
12125 => "0000000110100101",
12126 => "0000000110100101",
12127 => "0000000110100101",
12128 => "0000000110100101",
12129 => "0000000110100110",
12130 => "0000000110100110",
12131 => "0000000110100110",
12132 => "0000000110100110",
12133 => "0000000110100110",
12134 => "0000000110100110",
12135 => "0000000110100110",
12136 => "0000000110100110",
12137 => "0000000110100110",
12138 => "0000000110100110",
12139 => "0000000110100111",
12140 => "0000000110100111",
12141 => "0000000110100111",
12142 => "0000000110100111",
12143 => "0000000110100111",
12144 => "0000000110100111",
12145 => "0000000110100111",
12146 => "0000000110100111",
12147 => "0000000110100111",
12148 => "0000000110100111",
12149 => "0000000110101000",
12150 => "0000000110101000",
12151 => "0000000110101000",
12152 => "0000000110101000",
12153 => "0000000110101000",
12154 => "0000000110101000",
12155 => "0000000110101000",
12156 => "0000000110101000",
12157 => "0000000110101000",
12158 => "0000000110101001",
12159 => "0000000110101001",
12160 => "0000000110101001",
12161 => "0000000110101001",
12162 => "0000000110101001",
12163 => "0000000110101001",
12164 => "0000000110101001",
12165 => "0000000110101001",
12166 => "0000000110101001",
12167 => "0000000110101001",
12168 => "0000000110101010",
12169 => "0000000110101010",
12170 => "0000000110101010",
12171 => "0000000110101010",
12172 => "0000000110101010",
12173 => "0000000110101010",
12174 => "0000000110101010",
12175 => "0000000110101010",
12176 => "0000000110101010",
12177 => "0000000110101010",
12178 => "0000000110101011",
12179 => "0000000110101011",
12180 => "0000000110101011",
12181 => "0000000110101011",
12182 => "0000000110101011",
12183 => "0000000110101011",
12184 => "0000000110101011",
12185 => "0000000110101011",
12186 => "0000000110101011",
12187 => "0000000110101100",
12188 => "0000000110101100",
12189 => "0000000110101100",
12190 => "0000000110101100",
12191 => "0000000110101100",
12192 => "0000000110101100",
12193 => "0000000110101100",
12194 => "0000000110101100",
12195 => "0000000110101100",
12196 => "0000000110101100",
12197 => "0000000110101101",
12198 => "0000000110101101",
12199 => "0000000110101101",
12200 => "0000000110101101",
12201 => "0000000110101101",
12202 => "0000000110101101",
12203 => "0000000110101101",
12204 => "0000000110101101",
12205 => "0000000110101101",
12206 => "0000000110101110",
12207 => "0000000110101110",
12208 => "0000000110101110",
12209 => "0000000110101110",
12210 => "0000000110101110",
12211 => "0000000110101110",
12212 => "0000000110101110",
12213 => "0000000110101110",
12214 => "0000000110101110",
12215 => "0000000110101110",
12216 => "0000000110101111",
12217 => "0000000110101111",
12218 => "0000000110101111",
12219 => "0000000110101111",
12220 => "0000000110101111",
12221 => "0000000110101111",
12222 => "0000000110101111",
12223 => "0000000110101111",
12224 => "0000000110101111",
12225 => "0000000110101111",
12226 => "0000000110110000",
12227 => "0000000110110000",
12228 => "0000000110110000",
12229 => "0000000110110000",
12230 => "0000000110110000",
12231 => "0000000110110000",
12232 => "0000000110110000",
12233 => "0000000110110000",
12234 => "0000000110110000",
12235 => "0000000110110001",
12236 => "0000000110110001",
12237 => "0000000110110001",
12238 => "0000000110110001",
12239 => "0000000110110001",
12240 => "0000000110110001",
12241 => "0000000110110001",
12242 => "0000000110110001",
12243 => "0000000110110001",
12244 => "0000000110110001",
12245 => "0000000110110010",
12246 => "0000000110110010",
12247 => "0000000110110010",
12248 => "0000000110110010",
12249 => "0000000110110010",
12250 => "0000000110110010",
12251 => "0000000110110010",
12252 => "0000000110110010",
12253 => "0000000110110010",
12254 => "0000000110110011",
12255 => "0000000110110011",
12256 => "0000000110110011",
12257 => "0000000110110011",
12258 => "0000000110110011",
12259 => "0000000110110011",
12260 => "0000000110110011",
12261 => "0000000110110011",
12262 => "0000000110110011",
12263 => "0000000110110011",
12264 => "0000000110110100",
12265 => "0000000110110100",
12266 => "0000000110110100",
12267 => "0000000110110100",
12268 => "0000000110110100",
12269 => "0000000110110100",
12270 => "0000000110110100",
12271 => "0000000110110100",
12272 => "0000000110110100",
12273 => "0000000110110101",
12274 => "0000000110110101",
12275 => "0000000110110101",
12276 => "0000000110110101",
12277 => "0000000110110101",
12278 => "0000000110110101",
12279 => "0000000110110101",
12280 => "0000000110110101",
12281 => "0000000110110101",
12282 => "0000000110110110",
12283 => "0000000110110110",
12284 => "0000000110110110",
12285 => "0000000110110110",
12286 => "0000000110110110",
12287 => "0000000110110110",
12288 => "0000000110110110",
12289 => "0000000110110110",
12290 => "0000000110110110",
12291 => "0000000110110110",
12292 => "0000000110110111",
12293 => "0000000110110111",
12294 => "0000000110110111",
12295 => "0000000110110111",
12296 => "0000000110110111",
12297 => "0000000110110111",
12298 => "0000000110110111",
12299 => "0000000110110111",
12300 => "0000000110110111",
12301 => "0000000110111000",
12302 => "0000000110111000",
12303 => "0000000110111000",
12304 => "0000000110111000",
12305 => "0000000110111000",
12306 => "0000000110111000",
12307 => "0000000110111000",
12308 => "0000000110111000",
12309 => "0000000110111000",
12310 => "0000000110111000",
12311 => "0000000110111001",
12312 => "0000000110111001",
12313 => "0000000110111001",
12314 => "0000000110111001",
12315 => "0000000110111001",
12316 => "0000000110111001",
12317 => "0000000110111001",
12318 => "0000000110111001",
12319 => "0000000110111001",
12320 => "0000000110111010",
12321 => "0000000110111010",
12322 => "0000000110111010",
12323 => "0000000110111010",
12324 => "0000000110111010",
12325 => "0000000110111010",
12326 => "0000000110111010",
12327 => "0000000110111010",
12328 => "0000000110111010",
12329 => "0000000110111011",
12330 => "0000000110111011",
12331 => "0000000110111011",
12332 => "0000000110111011",
12333 => "0000000110111011",
12334 => "0000000110111011",
12335 => "0000000110111011",
12336 => "0000000110111011",
12337 => "0000000110111011",
12338 => "0000000110111011",
12339 => "0000000110111100",
12340 => "0000000110111100",
12341 => "0000000110111100",
12342 => "0000000110111100",
12343 => "0000000110111100",
12344 => "0000000110111100",
12345 => "0000000110111100",
12346 => "0000000110111100",
12347 => "0000000110111100",
12348 => "0000000110111101",
12349 => "0000000110111101",
12350 => "0000000110111101",
12351 => "0000000110111101",
12352 => "0000000110111101",
12353 => "0000000110111101",
12354 => "0000000110111101",
12355 => "0000000110111101",
12356 => "0000000110111101",
12357 => "0000000110111110",
12358 => "0000000110111110",
12359 => "0000000110111110",
12360 => "0000000110111110",
12361 => "0000000110111110",
12362 => "0000000110111110",
12363 => "0000000110111110",
12364 => "0000000110111110",
12365 => "0000000110111110",
12366 => "0000000110111111",
12367 => "0000000110111111",
12368 => "0000000110111111",
12369 => "0000000110111111",
12370 => "0000000110111111",
12371 => "0000000110111111",
12372 => "0000000110111111",
12373 => "0000000110111111",
12374 => "0000000110111111",
12375 => "0000000110111111",
12376 => "0000000111000000",
12377 => "0000000111000000",
12378 => "0000000111000000",
12379 => "0000000111000000",
12380 => "0000000111000000",
12381 => "0000000111000000",
12382 => "0000000111000000",
12383 => "0000000111000000",
12384 => "0000000111000000",
12385 => "0000000111000001",
12386 => "0000000111000001",
12387 => "0000000111000001",
12388 => "0000000111000001",
12389 => "0000000111000001",
12390 => "0000000111000001",
12391 => "0000000111000001",
12392 => "0000000111000001",
12393 => "0000000111000001",
12394 => "0000000111000010",
12395 => "0000000111000010",
12396 => "0000000111000010",
12397 => "0000000111000010",
12398 => "0000000111000010",
12399 => "0000000111000010",
12400 => "0000000111000010",
12401 => "0000000111000010",
12402 => "0000000111000010",
12403 => "0000000111000011",
12404 => "0000000111000011",
12405 => "0000000111000011",
12406 => "0000000111000011",
12407 => "0000000111000011",
12408 => "0000000111000011",
12409 => "0000000111000011",
12410 => "0000000111000011",
12411 => "0000000111000011",
12412 => "0000000111000100",
12413 => "0000000111000100",
12414 => "0000000111000100",
12415 => "0000000111000100",
12416 => "0000000111000100",
12417 => "0000000111000100",
12418 => "0000000111000100",
12419 => "0000000111000100",
12420 => "0000000111000100",
12421 => "0000000111000101",
12422 => "0000000111000101",
12423 => "0000000111000101",
12424 => "0000000111000101",
12425 => "0000000111000101",
12426 => "0000000111000101",
12427 => "0000000111000101",
12428 => "0000000111000101",
12429 => "0000000111000101",
12430 => "0000000111000110",
12431 => "0000000111000110",
12432 => "0000000111000110",
12433 => "0000000111000110",
12434 => "0000000111000110",
12435 => "0000000111000110",
12436 => "0000000111000110",
12437 => "0000000111000110",
12438 => "0000000111000110",
12439 => "0000000111000111",
12440 => "0000000111000111",
12441 => "0000000111000111",
12442 => "0000000111000111",
12443 => "0000000111000111",
12444 => "0000000111000111",
12445 => "0000000111000111",
12446 => "0000000111000111",
12447 => "0000000111000111",
12448 => "0000000111000111",
12449 => "0000000111001000",
12450 => "0000000111001000",
12451 => "0000000111001000",
12452 => "0000000111001000",
12453 => "0000000111001000",
12454 => "0000000111001000",
12455 => "0000000111001000",
12456 => "0000000111001000",
12457 => "0000000111001000",
12458 => "0000000111001001",
12459 => "0000000111001001",
12460 => "0000000111001001",
12461 => "0000000111001001",
12462 => "0000000111001001",
12463 => "0000000111001001",
12464 => "0000000111001001",
12465 => "0000000111001001",
12466 => "0000000111001001",
12467 => "0000000111001010",
12468 => "0000000111001010",
12469 => "0000000111001010",
12470 => "0000000111001010",
12471 => "0000000111001010",
12472 => "0000000111001010",
12473 => "0000000111001010",
12474 => "0000000111001010",
12475 => "0000000111001010",
12476 => "0000000111001011",
12477 => "0000000111001011",
12478 => "0000000111001011",
12479 => "0000000111001011",
12480 => "0000000111001011",
12481 => "0000000111001011",
12482 => "0000000111001011",
12483 => "0000000111001011",
12484 => "0000000111001011",
12485 => "0000000111001100",
12486 => "0000000111001100",
12487 => "0000000111001100",
12488 => "0000000111001100",
12489 => "0000000111001100",
12490 => "0000000111001100",
12491 => "0000000111001100",
12492 => "0000000111001100",
12493 => "0000000111001100",
12494 => "0000000111001101",
12495 => "0000000111001101",
12496 => "0000000111001101",
12497 => "0000000111001101",
12498 => "0000000111001101",
12499 => "0000000111001101",
12500 => "0000000111001101",
12501 => "0000000111001101",
12502 => "0000000111001110",
12503 => "0000000111001110",
12504 => "0000000111001110",
12505 => "0000000111001110",
12506 => "0000000111001110",
12507 => "0000000111001110",
12508 => "0000000111001110",
12509 => "0000000111001110",
12510 => "0000000111001110",
12511 => "0000000111001111",
12512 => "0000000111001111",
12513 => "0000000111001111",
12514 => "0000000111001111",
12515 => "0000000111001111",
12516 => "0000000111001111",
12517 => "0000000111001111",
12518 => "0000000111001111",
12519 => "0000000111001111",
12520 => "0000000111010000",
12521 => "0000000111010000",
12522 => "0000000111010000",
12523 => "0000000111010000",
12524 => "0000000111010000",
12525 => "0000000111010000",
12526 => "0000000111010000",
12527 => "0000000111010000",
12528 => "0000000111010000",
12529 => "0000000111010001",
12530 => "0000000111010001",
12531 => "0000000111010001",
12532 => "0000000111010001",
12533 => "0000000111010001",
12534 => "0000000111010001",
12535 => "0000000111010001",
12536 => "0000000111010001",
12537 => "0000000111010001",
12538 => "0000000111010010",
12539 => "0000000111010010",
12540 => "0000000111010010",
12541 => "0000000111010010",
12542 => "0000000111010010",
12543 => "0000000111010010",
12544 => "0000000111010010",
12545 => "0000000111010010",
12546 => "0000000111010010",
12547 => "0000000111010011",
12548 => "0000000111010011",
12549 => "0000000111010011",
12550 => "0000000111010011",
12551 => "0000000111010011",
12552 => "0000000111010011",
12553 => "0000000111010011",
12554 => "0000000111010011",
12555 => "0000000111010011",
12556 => "0000000111010100",
12557 => "0000000111010100",
12558 => "0000000111010100",
12559 => "0000000111010100",
12560 => "0000000111010100",
12561 => "0000000111010100",
12562 => "0000000111010100",
12563 => "0000000111010100",
12564 => "0000000111010100",
12565 => "0000000111010101",
12566 => "0000000111010101",
12567 => "0000000111010101",
12568 => "0000000111010101",
12569 => "0000000111010101",
12570 => "0000000111010101",
12571 => "0000000111010101",
12572 => "0000000111010101",
12573 => "0000000111010110",
12574 => "0000000111010110",
12575 => "0000000111010110",
12576 => "0000000111010110",
12577 => "0000000111010110",
12578 => "0000000111010110",
12579 => "0000000111010110",
12580 => "0000000111010110",
12581 => "0000000111010110",
12582 => "0000000111010111",
12583 => "0000000111010111",
12584 => "0000000111010111",
12585 => "0000000111010111",
12586 => "0000000111010111",
12587 => "0000000111010111",
12588 => "0000000111010111",
12589 => "0000000111010111",
12590 => "0000000111010111",
12591 => "0000000111011000",
12592 => "0000000111011000",
12593 => "0000000111011000",
12594 => "0000000111011000",
12595 => "0000000111011000",
12596 => "0000000111011000",
12597 => "0000000111011000",
12598 => "0000000111011000",
12599 => "0000000111011000",
12600 => "0000000111011001",
12601 => "0000000111011001",
12602 => "0000000111011001",
12603 => "0000000111011001",
12604 => "0000000111011001",
12605 => "0000000111011001",
12606 => "0000000111011001",
12607 => "0000000111011001",
12608 => "0000000111011010",
12609 => "0000000111011010",
12610 => "0000000111011010",
12611 => "0000000111011010",
12612 => "0000000111011010",
12613 => "0000000111011010",
12614 => "0000000111011010",
12615 => "0000000111011010",
12616 => "0000000111011010",
12617 => "0000000111011011",
12618 => "0000000111011011",
12619 => "0000000111011011",
12620 => "0000000111011011",
12621 => "0000000111011011",
12622 => "0000000111011011",
12623 => "0000000111011011",
12624 => "0000000111011011",
12625 => "0000000111011011",
12626 => "0000000111011100",
12627 => "0000000111011100",
12628 => "0000000111011100",
12629 => "0000000111011100",
12630 => "0000000111011100",
12631 => "0000000111011100",
12632 => "0000000111011100",
12633 => "0000000111011100",
12634 => "0000000111011101",
12635 => "0000000111011101",
12636 => "0000000111011101",
12637 => "0000000111011101",
12638 => "0000000111011101",
12639 => "0000000111011101",
12640 => "0000000111011101",
12641 => "0000000111011101",
12642 => "0000000111011101",
12643 => "0000000111011110",
12644 => "0000000111011110",
12645 => "0000000111011110",
12646 => "0000000111011110",
12647 => "0000000111011110",
12648 => "0000000111011110",
12649 => "0000000111011110",
12650 => "0000000111011110",
12651 => "0000000111011110",
12652 => "0000000111011111",
12653 => "0000000111011111",
12654 => "0000000111011111",
12655 => "0000000111011111",
12656 => "0000000111011111",
12657 => "0000000111011111",
12658 => "0000000111011111",
12659 => "0000000111011111",
12660 => "0000000111100000",
12661 => "0000000111100000",
12662 => "0000000111100000",
12663 => "0000000111100000",
12664 => "0000000111100000",
12665 => "0000000111100000",
12666 => "0000000111100000",
12667 => "0000000111100000",
12668 => "0000000111100000",
12669 => "0000000111100001",
12670 => "0000000111100001",
12671 => "0000000111100001",
12672 => "0000000111100001",
12673 => "0000000111100001",
12674 => "0000000111100001",
12675 => "0000000111100001",
12676 => "0000000111100001",
12677 => "0000000111100010",
12678 => "0000000111100010",
12679 => "0000000111100010",
12680 => "0000000111100010",
12681 => "0000000111100010",
12682 => "0000000111100010",
12683 => "0000000111100010",
12684 => "0000000111100010",
12685 => "0000000111100010",
12686 => "0000000111100011",
12687 => "0000000111100011",
12688 => "0000000111100011",
12689 => "0000000111100011",
12690 => "0000000111100011",
12691 => "0000000111100011",
12692 => "0000000111100011",
12693 => "0000000111100011",
12694 => "0000000111100100",
12695 => "0000000111100100",
12696 => "0000000111100100",
12697 => "0000000111100100",
12698 => "0000000111100100",
12699 => "0000000111100100",
12700 => "0000000111100100",
12701 => "0000000111100100",
12702 => "0000000111100100",
12703 => "0000000111100101",
12704 => "0000000111100101",
12705 => "0000000111100101",
12706 => "0000000111100101",
12707 => "0000000111100101",
12708 => "0000000111100101",
12709 => "0000000111100101",
12710 => "0000000111100101",
12711 => "0000000111100110",
12712 => "0000000111100110",
12713 => "0000000111100110",
12714 => "0000000111100110",
12715 => "0000000111100110",
12716 => "0000000111100110",
12717 => "0000000111100110",
12718 => "0000000111100110",
12719 => "0000000111100110",
12720 => "0000000111100111",
12721 => "0000000111100111",
12722 => "0000000111100111",
12723 => "0000000111100111",
12724 => "0000000111100111",
12725 => "0000000111100111",
12726 => "0000000111100111",
12727 => "0000000111100111",
12728 => "0000000111101000",
12729 => "0000000111101000",
12730 => "0000000111101000",
12731 => "0000000111101000",
12732 => "0000000111101000",
12733 => "0000000111101000",
12734 => "0000000111101000",
12735 => "0000000111101000",
12736 => "0000000111101000",
12737 => "0000000111101001",
12738 => "0000000111101001",
12739 => "0000000111101001",
12740 => "0000000111101001",
12741 => "0000000111101001",
12742 => "0000000111101001",
12743 => "0000000111101001",
12744 => "0000000111101001",
12745 => "0000000111101010",
12746 => "0000000111101010",
12747 => "0000000111101010",
12748 => "0000000111101010",
12749 => "0000000111101010",
12750 => "0000000111101010",
12751 => "0000000111101010",
12752 => "0000000111101010",
12753 => "0000000111101010",
12754 => "0000000111101011",
12755 => "0000000111101011",
12756 => "0000000111101011",
12757 => "0000000111101011",
12758 => "0000000111101011",
12759 => "0000000111101011",
12760 => "0000000111101011",
12761 => "0000000111101011",
12762 => "0000000111101100",
12763 => "0000000111101100",
12764 => "0000000111101100",
12765 => "0000000111101100",
12766 => "0000000111101100",
12767 => "0000000111101100",
12768 => "0000000111101100",
12769 => "0000000111101100",
12770 => "0000000111101101",
12771 => "0000000111101101",
12772 => "0000000111101101",
12773 => "0000000111101101",
12774 => "0000000111101101",
12775 => "0000000111101101",
12776 => "0000000111101101",
12777 => "0000000111101101",
12778 => "0000000111101101",
12779 => "0000000111101110",
12780 => "0000000111101110",
12781 => "0000000111101110",
12782 => "0000000111101110",
12783 => "0000000111101110",
12784 => "0000000111101110",
12785 => "0000000111101110",
12786 => "0000000111101110",
12787 => "0000000111101111",
12788 => "0000000111101111",
12789 => "0000000111101111",
12790 => "0000000111101111",
12791 => "0000000111101111",
12792 => "0000000111101111",
12793 => "0000000111101111",
12794 => "0000000111101111",
12795 => "0000000111110000",
12796 => "0000000111110000",
12797 => "0000000111110000",
12798 => "0000000111110000",
12799 => "0000000111110000",
12800 => "0000000111110000",
12801 => "0000000111110000",
12802 => "0000000111110000",
12803 => "0000000111110000",
12804 => "0000000111110001",
12805 => "0000000111110001",
12806 => "0000000111110001",
12807 => "0000000111110001",
12808 => "0000000111110001",
12809 => "0000000111110001",
12810 => "0000000111110001",
12811 => "0000000111110001",
12812 => "0000000111110010",
12813 => "0000000111110010",
12814 => "0000000111110010",
12815 => "0000000111110010",
12816 => "0000000111110010",
12817 => "0000000111110010",
12818 => "0000000111110010",
12819 => "0000000111110010",
12820 => "0000000111110011",
12821 => "0000000111110011",
12822 => "0000000111110011",
12823 => "0000000111110011",
12824 => "0000000111110011",
12825 => "0000000111110011",
12826 => "0000000111110011",
12827 => "0000000111110011",
12828 => "0000000111110011",
12829 => "0000000111110100",
12830 => "0000000111110100",
12831 => "0000000111110100",
12832 => "0000000111110100",
12833 => "0000000111110100",
12834 => "0000000111110100",
12835 => "0000000111110100",
12836 => "0000000111110100",
12837 => "0000000111110101",
12838 => "0000000111110101",
12839 => "0000000111110101",
12840 => "0000000111110101",
12841 => "0000000111110101",
12842 => "0000000111110101",
12843 => "0000000111110101",
12844 => "0000000111110101",
12845 => "0000000111110110",
12846 => "0000000111110110",
12847 => "0000000111110110",
12848 => "0000000111110110",
12849 => "0000000111110110",
12850 => "0000000111110110",
12851 => "0000000111110110",
12852 => "0000000111110110",
12853 => "0000000111110111",
12854 => "0000000111110111",
12855 => "0000000111110111",
12856 => "0000000111110111",
12857 => "0000000111110111",
12858 => "0000000111110111",
12859 => "0000000111110111",
12860 => "0000000111110111",
12861 => "0000000111110111",
12862 => "0000000111111000",
12863 => "0000000111111000",
12864 => "0000000111111000",
12865 => "0000000111111000",
12866 => "0000000111111000",
12867 => "0000000111111000",
12868 => "0000000111111000",
12869 => "0000000111111000",
12870 => "0000000111111001",
12871 => "0000000111111001",
12872 => "0000000111111001",
12873 => "0000000111111001",
12874 => "0000000111111001",
12875 => "0000000111111001",
12876 => "0000000111111001",
12877 => "0000000111111001",
12878 => "0000000111111010",
12879 => "0000000111111010",
12880 => "0000000111111010",
12881 => "0000000111111010",
12882 => "0000000111111010",
12883 => "0000000111111010",
12884 => "0000000111111010",
12885 => "0000000111111010",
12886 => "0000000111111011",
12887 => "0000000111111011",
12888 => "0000000111111011",
12889 => "0000000111111011",
12890 => "0000000111111011",
12891 => "0000000111111011",
12892 => "0000000111111011",
12893 => "0000000111111011",
12894 => "0000000111111100",
12895 => "0000000111111100",
12896 => "0000000111111100",
12897 => "0000000111111100",
12898 => "0000000111111100",
12899 => "0000000111111100",
12900 => "0000000111111100",
12901 => "0000000111111100",
12902 => "0000000111111101",
12903 => "0000000111111101",
12904 => "0000000111111101",
12905 => "0000000111111101",
12906 => "0000000111111101",
12907 => "0000000111111101",
12908 => "0000000111111101",
12909 => "0000000111111101",
12910 => "0000000111111110",
12911 => "0000000111111110",
12912 => "0000000111111110",
12913 => "0000000111111110",
12914 => "0000000111111110",
12915 => "0000000111111110",
12916 => "0000000111111110",
12917 => "0000000111111110",
12918 => "0000000111111111",
12919 => "0000000111111111",
12920 => "0000000111111111",
12921 => "0000000111111111",
12922 => "0000000111111111",
12923 => "0000000111111111",
12924 => "0000000111111111",
12925 => "0000000111111111",
12926 => "0000000111111111",
12927 => "0000001000000000",
12928 => "0000001000000000",
12929 => "0000001000000000",
12930 => "0000001000000000",
12931 => "0000001000000000",
12932 => "0000001000000000",
12933 => "0000001000000000",
12934 => "0000001000000000",
12935 => "0000001000000001",
12936 => "0000001000000001",
12937 => "0000001000000001",
12938 => "0000001000000001",
12939 => "0000001000000001",
12940 => "0000001000000001",
12941 => "0000001000000001",
12942 => "0000001000000001",
12943 => "0000001000000010",
12944 => "0000001000000010",
12945 => "0000001000000010",
12946 => "0000001000000010",
12947 => "0000001000000010",
12948 => "0000001000000010",
12949 => "0000001000000010",
12950 => "0000001000000010",
12951 => "0000001000000011",
12952 => "0000001000000011",
12953 => "0000001000000011",
12954 => "0000001000000011",
12955 => "0000001000000011",
12956 => "0000001000000011",
12957 => "0000001000000011",
12958 => "0000001000000011",
12959 => "0000001000000100",
12960 => "0000001000000100",
12961 => "0000001000000100",
12962 => "0000001000000100",
12963 => "0000001000000100",
12964 => "0000001000000100",
12965 => "0000001000000100",
12966 => "0000001000000100",
12967 => "0000001000000101",
12968 => "0000001000000101",
12969 => "0000001000000101",
12970 => "0000001000000101",
12971 => "0000001000000101",
12972 => "0000001000000101",
12973 => "0000001000000101",
12974 => "0000001000000101",
12975 => "0000001000000110",
12976 => "0000001000000110",
12977 => "0000001000000110",
12978 => "0000001000000110",
12979 => "0000001000000110",
12980 => "0000001000000110",
12981 => "0000001000000110",
12982 => "0000001000000110",
12983 => "0000001000000111",
12984 => "0000001000000111",
12985 => "0000001000000111",
12986 => "0000001000000111",
12987 => "0000001000000111",
12988 => "0000001000000111",
12989 => "0000001000000111",
12990 => "0000001000000111",
12991 => "0000001000001000",
12992 => "0000001000001000",
12993 => "0000001000001000",
12994 => "0000001000001000",
12995 => "0000001000001000",
12996 => "0000001000001000",
12997 => "0000001000001000",
12998 => "0000001000001001",
12999 => "0000001000001001",
13000 => "0000001000001001",
13001 => "0000001000001001",
13002 => "0000001000001001",
13003 => "0000001000001001",
13004 => "0000001000001001",
13005 => "0000001000001001",
13006 => "0000001000001010",
13007 => "0000001000001010",
13008 => "0000001000001010",
13009 => "0000001000001010",
13010 => "0000001000001010",
13011 => "0000001000001010",
13012 => "0000001000001010",
13013 => "0000001000001010",
13014 => "0000001000001011",
13015 => "0000001000001011",
13016 => "0000001000001011",
13017 => "0000001000001011",
13018 => "0000001000001011",
13019 => "0000001000001011",
13020 => "0000001000001011",
13021 => "0000001000001011",
13022 => "0000001000001100",
13023 => "0000001000001100",
13024 => "0000001000001100",
13025 => "0000001000001100",
13026 => "0000001000001100",
13027 => "0000001000001100",
13028 => "0000001000001100",
13029 => "0000001000001100",
13030 => "0000001000001101",
13031 => "0000001000001101",
13032 => "0000001000001101",
13033 => "0000001000001101",
13034 => "0000001000001101",
13035 => "0000001000001101",
13036 => "0000001000001101",
13037 => "0000001000001101",
13038 => "0000001000001110",
13039 => "0000001000001110",
13040 => "0000001000001110",
13041 => "0000001000001110",
13042 => "0000001000001110",
13043 => "0000001000001110",
13044 => "0000001000001110",
13045 => "0000001000001110",
13046 => "0000001000001111",
13047 => "0000001000001111",
13048 => "0000001000001111",
13049 => "0000001000001111",
13050 => "0000001000001111",
13051 => "0000001000001111",
13052 => "0000001000001111",
13053 => "0000001000001111",
13054 => "0000001000010000",
13055 => "0000001000010000",
13056 => "0000001000010000",
13057 => "0000001000010000",
13058 => "0000001000010000",
13059 => "0000001000010000",
13060 => "0000001000010000",
13061 => "0000001000010001",
13062 => "0000001000010001",
13063 => "0000001000010001",
13064 => "0000001000010001",
13065 => "0000001000010001",
13066 => "0000001000010001",
13067 => "0000001000010001",
13068 => "0000001000010001",
13069 => "0000001000010010",
13070 => "0000001000010010",
13071 => "0000001000010010",
13072 => "0000001000010010",
13073 => "0000001000010010",
13074 => "0000001000010010",
13075 => "0000001000010010",
13076 => "0000001000010010",
13077 => "0000001000010011",
13078 => "0000001000010011",
13079 => "0000001000010011",
13080 => "0000001000010011",
13081 => "0000001000010011",
13082 => "0000001000010011",
13083 => "0000001000010011",
13084 => "0000001000010011",
13085 => "0000001000010100",
13086 => "0000001000010100",
13087 => "0000001000010100",
13088 => "0000001000010100",
13089 => "0000001000010100",
13090 => "0000001000010100",
13091 => "0000001000010100",
13092 => "0000001000010101",
13093 => "0000001000010101",
13094 => "0000001000010101",
13095 => "0000001000010101",
13096 => "0000001000010101",
13097 => "0000001000010101",
13098 => "0000001000010101",
13099 => "0000001000010101",
13100 => "0000001000010110",
13101 => "0000001000010110",
13102 => "0000001000010110",
13103 => "0000001000010110",
13104 => "0000001000010110",
13105 => "0000001000010110",
13106 => "0000001000010110",
13107 => "0000001000010110",
13108 => "0000001000010111",
13109 => "0000001000010111",
13110 => "0000001000010111",
13111 => "0000001000010111",
13112 => "0000001000010111",
13113 => "0000001000010111",
13114 => "0000001000010111",
13115 => "0000001000010111",
13116 => "0000001000011000",
13117 => "0000001000011000",
13118 => "0000001000011000",
13119 => "0000001000011000",
13120 => "0000001000011000",
13121 => "0000001000011000",
13122 => "0000001000011000",
13123 => "0000001000011001",
13124 => "0000001000011001",
13125 => "0000001000011001",
13126 => "0000001000011001",
13127 => "0000001000011001",
13128 => "0000001000011001",
13129 => "0000001000011001",
13130 => "0000001000011001",
13131 => "0000001000011010",
13132 => "0000001000011010",
13133 => "0000001000011010",
13134 => "0000001000011010",
13135 => "0000001000011010",
13136 => "0000001000011010",
13137 => "0000001000011010",
13138 => "0000001000011010",
13139 => "0000001000011011",
13140 => "0000001000011011",
13141 => "0000001000011011",
13142 => "0000001000011011",
13143 => "0000001000011011",
13144 => "0000001000011011",
13145 => "0000001000011011",
13146 => "0000001000011100",
13147 => "0000001000011100",
13148 => "0000001000011100",
13149 => "0000001000011100",
13150 => "0000001000011100",
13151 => "0000001000011100",
13152 => "0000001000011100",
13153 => "0000001000011100",
13154 => "0000001000011101",
13155 => "0000001000011101",
13156 => "0000001000011101",
13157 => "0000001000011101",
13158 => "0000001000011101",
13159 => "0000001000011101",
13160 => "0000001000011101",
13161 => "0000001000011101",
13162 => "0000001000011110",
13163 => "0000001000011110",
13164 => "0000001000011110",
13165 => "0000001000011110",
13166 => "0000001000011110",
13167 => "0000001000011110",
13168 => "0000001000011110",
13169 => "0000001000011111",
13170 => "0000001000011111",
13171 => "0000001000011111",
13172 => "0000001000011111",
13173 => "0000001000011111",
13174 => "0000001000011111",
13175 => "0000001000011111",
13176 => "0000001000011111",
13177 => "0000001000100000",
13178 => "0000001000100000",
13179 => "0000001000100000",
13180 => "0000001000100000",
13181 => "0000001000100000",
13182 => "0000001000100000",
13183 => "0000001000100000",
13184 => "0000001000100001",
13185 => "0000001000100001",
13186 => "0000001000100001",
13187 => "0000001000100001",
13188 => "0000001000100001",
13189 => "0000001000100001",
13190 => "0000001000100001",
13191 => "0000001000100001",
13192 => "0000001000100010",
13193 => "0000001000100010",
13194 => "0000001000100010",
13195 => "0000001000100010",
13196 => "0000001000100010",
13197 => "0000001000100010",
13198 => "0000001000100010",
13199 => "0000001000100010",
13200 => "0000001000100011",
13201 => "0000001000100011",
13202 => "0000001000100011",
13203 => "0000001000100011",
13204 => "0000001000100011",
13205 => "0000001000100011",
13206 => "0000001000100011",
13207 => "0000001000100100",
13208 => "0000001000100100",
13209 => "0000001000100100",
13210 => "0000001000100100",
13211 => "0000001000100100",
13212 => "0000001000100100",
13213 => "0000001000100100",
13214 => "0000001000100100",
13215 => "0000001000100101",
13216 => "0000001000100101",
13217 => "0000001000100101",
13218 => "0000001000100101",
13219 => "0000001000100101",
13220 => "0000001000100101",
13221 => "0000001000100101",
13222 => "0000001000100110",
13223 => "0000001000100110",
13224 => "0000001000100110",
13225 => "0000001000100110",
13226 => "0000001000100110",
13227 => "0000001000100110",
13228 => "0000001000100110",
13229 => "0000001000100110",
13230 => "0000001000100111",
13231 => "0000001000100111",
13232 => "0000001000100111",
13233 => "0000001000100111",
13234 => "0000001000100111",
13235 => "0000001000100111",
13236 => "0000001000100111",
13237 => "0000001000101000",
13238 => "0000001000101000",
13239 => "0000001000101000",
13240 => "0000001000101000",
13241 => "0000001000101000",
13242 => "0000001000101000",
13243 => "0000001000101000",
13244 => "0000001000101000",
13245 => "0000001000101001",
13246 => "0000001000101001",
13247 => "0000001000101001",
13248 => "0000001000101001",
13249 => "0000001000101001",
13250 => "0000001000101001",
13251 => "0000001000101001",
13252 => "0000001000101010",
13253 => "0000001000101010",
13254 => "0000001000101010",
13255 => "0000001000101010",
13256 => "0000001000101010",
13257 => "0000001000101010",
13258 => "0000001000101010",
13259 => "0000001000101010",
13260 => "0000001000101011",
13261 => "0000001000101011",
13262 => "0000001000101011",
13263 => "0000001000101011",
13264 => "0000001000101011",
13265 => "0000001000101011",
13266 => "0000001000101011",
13267 => "0000001000101100",
13268 => "0000001000101100",
13269 => "0000001000101100",
13270 => "0000001000101100",
13271 => "0000001000101100",
13272 => "0000001000101100",
13273 => "0000001000101100",
13274 => "0000001000101101",
13275 => "0000001000101101",
13276 => "0000001000101101",
13277 => "0000001000101101",
13278 => "0000001000101101",
13279 => "0000001000101101",
13280 => "0000001000101101",
13281 => "0000001000101101",
13282 => "0000001000101110",
13283 => "0000001000101110",
13284 => "0000001000101110",
13285 => "0000001000101110",
13286 => "0000001000101110",
13287 => "0000001000101110",
13288 => "0000001000101110",
13289 => "0000001000101111",
13290 => "0000001000101111",
13291 => "0000001000101111",
13292 => "0000001000101111",
13293 => "0000001000101111",
13294 => "0000001000101111",
13295 => "0000001000101111",
13296 => "0000001000101111",
13297 => "0000001000110000",
13298 => "0000001000110000",
13299 => "0000001000110000",
13300 => "0000001000110000",
13301 => "0000001000110000",
13302 => "0000001000110000",
13303 => "0000001000110000",
13304 => "0000001000110001",
13305 => "0000001000110001",
13306 => "0000001000110001",
13307 => "0000001000110001",
13308 => "0000001000110001",
13309 => "0000001000110001",
13310 => "0000001000110001",
13311 => "0000001000110010",
13312 => "0000001000110010",
13313 => "0000001000110010",
13314 => "0000001000110010",
13315 => "0000001000110010",
13316 => "0000001000110010",
13317 => "0000001000110010",
13318 => "0000001000110010",
13319 => "0000001000110011",
13320 => "0000001000110011",
13321 => "0000001000110011",
13322 => "0000001000110011",
13323 => "0000001000110011",
13324 => "0000001000110011",
13325 => "0000001000110011",
13326 => "0000001000110100",
13327 => "0000001000110100",
13328 => "0000001000110100",
13329 => "0000001000110100",
13330 => "0000001000110100",
13331 => "0000001000110100",
13332 => "0000001000110100",
13333 => "0000001000110101",
13334 => "0000001000110101",
13335 => "0000001000110101",
13336 => "0000001000110101",
13337 => "0000001000110101",
13338 => "0000001000110101",
13339 => "0000001000110101",
13340 => "0000001000110101",
13341 => "0000001000110110",
13342 => "0000001000110110",
13343 => "0000001000110110",
13344 => "0000001000110110",
13345 => "0000001000110110",
13346 => "0000001000110110",
13347 => "0000001000110110",
13348 => "0000001000110111",
13349 => "0000001000110111",
13350 => "0000001000110111",
13351 => "0000001000110111",
13352 => "0000001000110111",
13353 => "0000001000110111",
13354 => "0000001000110111",
13355 => "0000001000111000",
13356 => "0000001000111000",
13357 => "0000001000111000",
13358 => "0000001000111000",
13359 => "0000001000111000",
13360 => "0000001000111000",
13361 => "0000001000111000",
13362 => "0000001000111001",
13363 => "0000001000111001",
13364 => "0000001000111001",
13365 => "0000001000111001",
13366 => "0000001000111001",
13367 => "0000001000111001",
13368 => "0000001000111001",
13369 => "0000001000111001",
13370 => "0000001000111010",
13371 => "0000001000111010",
13372 => "0000001000111010",
13373 => "0000001000111010",
13374 => "0000001000111010",
13375 => "0000001000111010",
13376 => "0000001000111010",
13377 => "0000001000111011",
13378 => "0000001000111011",
13379 => "0000001000111011",
13380 => "0000001000111011",
13381 => "0000001000111011",
13382 => "0000001000111011",
13383 => "0000001000111011",
13384 => "0000001000111100",
13385 => "0000001000111100",
13386 => "0000001000111100",
13387 => "0000001000111100",
13388 => "0000001000111100",
13389 => "0000001000111100",
13390 => "0000001000111100",
13391 => "0000001000111101",
13392 => "0000001000111101",
13393 => "0000001000111101",
13394 => "0000001000111101",
13395 => "0000001000111101",
13396 => "0000001000111101",
13397 => "0000001000111101",
13398 => "0000001000111101",
13399 => "0000001000111110",
13400 => "0000001000111110",
13401 => "0000001000111110",
13402 => "0000001000111110",
13403 => "0000001000111110",
13404 => "0000001000111110",
13405 => "0000001000111110",
13406 => "0000001000111111",
13407 => "0000001000111111",
13408 => "0000001000111111",
13409 => "0000001000111111",
13410 => "0000001000111111",
13411 => "0000001000111111",
13412 => "0000001000111111",
13413 => "0000001001000000",
13414 => "0000001001000000",
13415 => "0000001001000000",
13416 => "0000001001000000",
13417 => "0000001001000000",
13418 => "0000001001000000",
13419 => "0000001001000000",
13420 => "0000001001000001",
13421 => "0000001001000001",
13422 => "0000001001000001",
13423 => "0000001001000001",
13424 => "0000001001000001",
13425 => "0000001001000001",
13426 => "0000001001000001",
13427 => "0000001001000010",
13428 => "0000001001000010",
13429 => "0000001001000010",
13430 => "0000001001000010",
13431 => "0000001001000010",
13432 => "0000001001000010",
13433 => "0000001001000010",
13434 => "0000001001000011",
13435 => "0000001001000011",
13436 => "0000001001000011",
13437 => "0000001001000011",
13438 => "0000001001000011",
13439 => "0000001001000011",
13440 => "0000001001000011",
13441 => "0000001001000011",
13442 => "0000001001000100",
13443 => "0000001001000100",
13444 => "0000001001000100",
13445 => "0000001001000100",
13446 => "0000001001000100",
13447 => "0000001001000100",
13448 => "0000001001000100",
13449 => "0000001001000101",
13450 => "0000001001000101",
13451 => "0000001001000101",
13452 => "0000001001000101",
13453 => "0000001001000101",
13454 => "0000001001000101",
13455 => "0000001001000101",
13456 => "0000001001000110",
13457 => "0000001001000110",
13458 => "0000001001000110",
13459 => "0000001001000110",
13460 => "0000001001000110",
13461 => "0000001001000110",
13462 => "0000001001000110",
13463 => "0000001001000111",
13464 => "0000001001000111",
13465 => "0000001001000111",
13466 => "0000001001000111",
13467 => "0000001001000111",
13468 => "0000001001000111",
13469 => "0000001001000111",
13470 => "0000001001001000",
13471 => "0000001001001000",
13472 => "0000001001001000",
13473 => "0000001001001000",
13474 => "0000001001001000",
13475 => "0000001001001000",
13476 => "0000001001001000",
13477 => "0000001001001001",
13478 => "0000001001001001",
13479 => "0000001001001001",
13480 => "0000001001001001",
13481 => "0000001001001001",
13482 => "0000001001001001",
13483 => "0000001001001001",
13484 => "0000001001001010",
13485 => "0000001001001010",
13486 => "0000001001001010",
13487 => "0000001001001010",
13488 => "0000001001001010",
13489 => "0000001001001010",
13490 => "0000001001001010",
13491 => "0000001001001011",
13492 => "0000001001001011",
13493 => "0000001001001011",
13494 => "0000001001001011",
13495 => "0000001001001011",
13496 => "0000001001001011",
13497 => "0000001001001011",
13498 => "0000001001001100",
13499 => "0000001001001100",
13500 => "0000001001001100",
13501 => "0000001001001100",
13502 => "0000001001001100",
13503 => "0000001001001100",
13504 => "0000001001001100",
13505 => "0000001001001101",
13506 => "0000001001001101",
13507 => "0000001001001101",
13508 => "0000001001001101",
13509 => "0000001001001101",
13510 => "0000001001001101",
13511 => "0000001001001101",
13512 => "0000001001001110",
13513 => "0000001001001110",
13514 => "0000001001001110",
13515 => "0000001001001110",
13516 => "0000001001001110",
13517 => "0000001001001110",
13518 => "0000001001001110",
13519 => "0000001001001111",
13520 => "0000001001001111",
13521 => "0000001001001111",
13522 => "0000001001001111",
13523 => "0000001001001111",
13524 => "0000001001001111",
13525 => "0000001001001111",
13526 => "0000001001010000",
13527 => "0000001001010000",
13528 => "0000001001010000",
13529 => "0000001001010000",
13530 => "0000001001010000",
13531 => "0000001001010000",
13532 => "0000001001010000",
13533 => "0000001001010001",
13534 => "0000001001010001",
13535 => "0000001001010001",
13536 => "0000001001010001",
13537 => "0000001001010001",
13538 => "0000001001010001",
13539 => "0000001001010001",
13540 => "0000001001010010",
13541 => "0000001001010010",
13542 => "0000001001010010",
13543 => "0000001001010010",
13544 => "0000001001010010",
13545 => "0000001001010010",
13546 => "0000001001010010",
13547 => "0000001001010011",
13548 => "0000001001010011",
13549 => "0000001001010011",
13550 => "0000001001010011",
13551 => "0000001001010011",
13552 => "0000001001010011",
13553 => "0000001001010011",
13554 => "0000001001010100",
13555 => "0000001001010100",
13556 => "0000001001010100",
13557 => "0000001001010100",
13558 => "0000001001010100",
13559 => "0000001001010100",
13560 => "0000001001010100",
13561 => "0000001001010101",
13562 => "0000001001010101",
13563 => "0000001001010101",
13564 => "0000001001010101",
13565 => "0000001001010101",
13566 => "0000001001010101",
13567 => "0000001001010101",
13568 => "0000001001010110",
13569 => "0000001001010110",
13570 => "0000001001010110",
13571 => "0000001001010110",
13572 => "0000001001010110",
13573 => "0000001001010110",
13574 => "0000001001010110",
13575 => "0000001001010111",
13576 => "0000001001010111",
13577 => "0000001001010111",
13578 => "0000001001010111",
13579 => "0000001001010111",
13580 => "0000001001010111",
13581 => "0000001001010111",
13582 => "0000001001011000",
13583 => "0000001001011000",
13584 => "0000001001011000",
13585 => "0000001001011000",
13586 => "0000001001011000",
13587 => "0000001001011000",
13588 => "0000001001011000",
13589 => "0000001001011001",
13590 => "0000001001011001",
13591 => "0000001001011001",
13592 => "0000001001011001",
13593 => "0000001001011001",
13594 => "0000001001011001",
13595 => "0000001001011010",
13596 => "0000001001011010",
13597 => "0000001001011010",
13598 => "0000001001011010",
13599 => "0000001001011010",
13600 => "0000001001011010",
13601 => "0000001001011010",
13602 => "0000001001011011",
13603 => "0000001001011011",
13604 => "0000001001011011",
13605 => "0000001001011011",
13606 => "0000001001011011",
13607 => "0000001001011011",
13608 => "0000001001011011",
13609 => "0000001001011100",
13610 => "0000001001011100",
13611 => "0000001001011100",
13612 => "0000001001011100",
13613 => "0000001001011100",
13614 => "0000001001011100",
13615 => "0000001001011100",
13616 => "0000001001011101",
13617 => "0000001001011101",
13618 => "0000001001011101",
13619 => "0000001001011101",
13620 => "0000001001011101",
13621 => "0000001001011101",
13622 => "0000001001011101",
13623 => "0000001001011110",
13624 => "0000001001011110",
13625 => "0000001001011110",
13626 => "0000001001011110",
13627 => "0000001001011110",
13628 => "0000001001011110",
13629 => "0000001001011110",
13630 => "0000001001011111",
13631 => "0000001001011111",
13632 => "0000001001011111",
13633 => "0000001001011111",
13634 => "0000001001011111",
13635 => "0000001001011111",
13636 => "0000001001100000",
13637 => "0000001001100000",
13638 => "0000001001100000",
13639 => "0000001001100000",
13640 => "0000001001100000",
13641 => "0000001001100000",
13642 => "0000001001100000",
13643 => "0000001001100001",
13644 => "0000001001100001",
13645 => "0000001001100001",
13646 => "0000001001100001",
13647 => "0000001001100001",
13648 => "0000001001100001",
13649 => "0000001001100001",
13650 => "0000001001100010",
13651 => "0000001001100010",
13652 => "0000001001100010",
13653 => "0000001001100010",
13654 => "0000001001100010",
13655 => "0000001001100010",
13656 => "0000001001100010",
13657 => "0000001001100011",
13658 => "0000001001100011",
13659 => "0000001001100011",
13660 => "0000001001100011",
13661 => "0000001001100011",
13662 => "0000001001100011",
13663 => "0000001001100011",
13664 => "0000001001100100",
13665 => "0000001001100100",
13666 => "0000001001100100",
13667 => "0000001001100100",
13668 => "0000001001100100",
13669 => "0000001001100100",
13670 => "0000001001100101",
13671 => "0000001001100101",
13672 => "0000001001100101",
13673 => "0000001001100101",
13674 => "0000001001100101",
13675 => "0000001001100101",
13676 => "0000001001100101",
13677 => "0000001001100110",
13678 => "0000001001100110",
13679 => "0000001001100110",
13680 => "0000001001100110",
13681 => "0000001001100110",
13682 => "0000001001100110",
13683 => "0000001001100110",
13684 => "0000001001100111",
13685 => "0000001001100111",
13686 => "0000001001100111",
13687 => "0000001001100111",
13688 => "0000001001100111",
13689 => "0000001001100111",
13690 => "0000001001101000",
13691 => "0000001001101000",
13692 => "0000001001101000",
13693 => "0000001001101000",
13694 => "0000001001101000",
13695 => "0000001001101000",
13696 => "0000001001101000",
13697 => "0000001001101001",
13698 => "0000001001101001",
13699 => "0000001001101001",
13700 => "0000001001101001",
13701 => "0000001001101001",
13702 => "0000001001101001",
13703 => "0000001001101001",
13704 => "0000001001101010",
13705 => "0000001001101010",
13706 => "0000001001101010",
13707 => "0000001001101010",
13708 => "0000001001101010",
13709 => "0000001001101010",
13710 => "0000001001101010",
13711 => "0000001001101011",
13712 => "0000001001101011",
13713 => "0000001001101011",
13714 => "0000001001101011",
13715 => "0000001001101011",
13716 => "0000001001101011",
13717 => "0000001001101100",
13718 => "0000001001101100",
13719 => "0000001001101100",
13720 => "0000001001101100",
13721 => "0000001001101100",
13722 => "0000001001101100",
13723 => "0000001001101100",
13724 => "0000001001101101",
13725 => "0000001001101101",
13726 => "0000001001101101",
13727 => "0000001001101101",
13728 => "0000001001101101",
13729 => "0000001001101101",
13730 => "0000001001101101",
13731 => "0000001001101110",
13732 => "0000001001101110",
13733 => "0000001001101110",
13734 => "0000001001101110",
13735 => "0000001001101110",
13736 => "0000001001101110",
13737 => "0000001001101111",
13738 => "0000001001101111",
13739 => "0000001001101111",
13740 => "0000001001101111",
13741 => "0000001001101111",
13742 => "0000001001101111",
13743 => "0000001001101111",
13744 => "0000001001110000",
13745 => "0000001001110000",
13746 => "0000001001110000",
13747 => "0000001001110000",
13748 => "0000001001110000",
13749 => "0000001001110000",
13750 => "0000001001110001",
13751 => "0000001001110001",
13752 => "0000001001110001",
13753 => "0000001001110001",
13754 => "0000001001110001",
13755 => "0000001001110001",
13756 => "0000001001110001",
13757 => "0000001001110010",
13758 => "0000001001110010",
13759 => "0000001001110010",
13760 => "0000001001110010",
13761 => "0000001001110010",
13762 => "0000001001110010",
13763 => "0000001001110010",
13764 => "0000001001110011",
13765 => "0000001001110011",
13766 => "0000001001110011",
13767 => "0000001001110011",
13768 => "0000001001110011",
13769 => "0000001001110011",
13770 => "0000001001110100",
13771 => "0000001001110100",
13772 => "0000001001110100",
13773 => "0000001001110100",
13774 => "0000001001110100",
13775 => "0000001001110100",
13776 => "0000001001110100",
13777 => "0000001001110101",
13778 => "0000001001110101",
13779 => "0000001001110101",
13780 => "0000001001110101",
13781 => "0000001001110101",
13782 => "0000001001110101",
13783 => "0000001001110110",
13784 => "0000001001110110",
13785 => "0000001001110110",
13786 => "0000001001110110",
13787 => "0000001001110110",
13788 => "0000001001110110",
13789 => "0000001001110110",
13790 => "0000001001110111",
13791 => "0000001001110111",
13792 => "0000001001110111",
13793 => "0000001001110111",
13794 => "0000001001110111",
13795 => "0000001001110111",
13796 => "0000001001110111",
13797 => "0000001001111000",
13798 => "0000001001111000",
13799 => "0000001001111000",
13800 => "0000001001111000",
13801 => "0000001001111000",
13802 => "0000001001111000",
13803 => "0000001001111001",
13804 => "0000001001111001",
13805 => "0000001001111001",
13806 => "0000001001111001",
13807 => "0000001001111001",
13808 => "0000001001111001",
13809 => "0000001001111001",
13810 => "0000001001111010",
13811 => "0000001001111010",
13812 => "0000001001111010",
13813 => "0000001001111010",
13814 => "0000001001111010",
13815 => "0000001001111010",
13816 => "0000001001111011",
13817 => "0000001001111011",
13818 => "0000001001111011",
13819 => "0000001001111011",
13820 => "0000001001111011",
13821 => "0000001001111011",
13822 => "0000001001111011",
13823 => "0000001001111100",
13824 => "0000001001111100",
13825 => "0000001001111100",
13826 => "0000001001111100",
13827 => "0000001001111100",
13828 => "0000001001111100",
13829 => "0000001001111101",
13830 => "0000001001111101",
13831 => "0000001001111101",
13832 => "0000001001111101",
13833 => "0000001001111101",
13834 => "0000001001111101",
13835 => "0000001001111101",
13836 => "0000001001111110",
13837 => "0000001001111110",
13838 => "0000001001111110",
13839 => "0000001001111110",
13840 => "0000001001111110",
13841 => "0000001001111110",
13842 => "0000001001111111",
13843 => "0000001001111111",
13844 => "0000001001111111",
13845 => "0000001001111111",
13846 => "0000001001111111",
13847 => "0000001001111111",
13848 => "0000001001111111",
13849 => "0000001010000000",
13850 => "0000001010000000",
13851 => "0000001010000000",
13852 => "0000001010000000",
13853 => "0000001010000000",
13854 => "0000001010000000",
13855 => "0000001010000001",
13856 => "0000001010000001",
13857 => "0000001010000001",
13858 => "0000001010000001",
13859 => "0000001010000001",
13860 => "0000001010000001",
13861 => "0000001010000010",
13862 => "0000001010000010",
13863 => "0000001010000010",
13864 => "0000001010000010",
13865 => "0000001010000010",
13866 => "0000001010000010",
13867 => "0000001010000010",
13868 => "0000001010000011",
13869 => "0000001010000011",
13870 => "0000001010000011",
13871 => "0000001010000011",
13872 => "0000001010000011",
13873 => "0000001010000011",
13874 => "0000001010000100",
13875 => "0000001010000100",
13876 => "0000001010000100",
13877 => "0000001010000100",
13878 => "0000001010000100",
13879 => "0000001010000100",
13880 => "0000001010000100",
13881 => "0000001010000101",
13882 => "0000001010000101",
13883 => "0000001010000101",
13884 => "0000001010000101",
13885 => "0000001010000101",
13886 => "0000001010000101",
13887 => "0000001010000110",
13888 => "0000001010000110",
13889 => "0000001010000110",
13890 => "0000001010000110",
13891 => "0000001010000110",
13892 => "0000001010000110",
13893 => "0000001010000110",
13894 => "0000001010000111",
13895 => "0000001010000111",
13896 => "0000001010000111",
13897 => "0000001010000111",
13898 => "0000001010000111",
13899 => "0000001010000111",
13900 => "0000001010001000",
13901 => "0000001010001000",
13902 => "0000001010001000",
13903 => "0000001010001000",
13904 => "0000001010001000",
13905 => "0000001010001000",
13906 => "0000001010001001",
13907 => "0000001010001001",
13908 => "0000001010001001",
13909 => "0000001010001001",
13910 => "0000001010001001",
13911 => "0000001010001001",
13912 => "0000001010001001",
13913 => "0000001010001010",
13914 => "0000001010001010",
13915 => "0000001010001010",
13916 => "0000001010001010",
13917 => "0000001010001010",
13918 => "0000001010001010",
13919 => "0000001010001011",
13920 => "0000001010001011",
13921 => "0000001010001011",
13922 => "0000001010001011",
13923 => "0000001010001011",
13924 => "0000001010001011",
13925 => "0000001010001100",
13926 => "0000001010001100",
13927 => "0000001010001100",
13928 => "0000001010001100",
13929 => "0000001010001100",
13930 => "0000001010001100",
13931 => "0000001010001100",
13932 => "0000001010001101",
13933 => "0000001010001101",
13934 => "0000001010001101",
13935 => "0000001010001101",
13936 => "0000001010001101",
13937 => "0000001010001101",
13938 => "0000001010001110",
13939 => "0000001010001110",
13940 => "0000001010001110",
13941 => "0000001010001110",
13942 => "0000001010001110",
13943 => "0000001010001110",
13944 => "0000001010001111",
13945 => "0000001010001111",
13946 => "0000001010001111",
13947 => "0000001010001111",
13948 => "0000001010001111",
13949 => "0000001010001111",
13950 => "0000001010001111",
13951 => "0000001010010000",
13952 => "0000001010010000",
13953 => "0000001010010000",
13954 => "0000001010010000",
13955 => "0000001010010000",
13956 => "0000001010010000",
13957 => "0000001010010001",
13958 => "0000001010010001",
13959 => "0000001010010001",
13960 => "0000001010010001",
13961 => "0000001010010001",
13962 => "0000001010010001",
13963 => "0000001010010010",
13964 => "0000001010010010",
13965 => "0000001010010010",
13966 => "0000001010010010",
13967 => "0000001010010010",
13968 => "0000001010010010",
13969 => "0000001010010010",
13970 => "0000001010010011",
13971 => "0000001010010011",
13972 => "0000001010010011",
13973 => "0000001010010011",
13974 => "0000001010010011",
13975 => "0000001010010011",
13976 => "0000001010010100",
13977 => "0000001010010100",
13978 => "0000001010010100",
13979 => "0000001010010100",
13980 => "0000001010010100",
13981 => "0000001010010100",
13982 => "0000001010010101",
13983 => "0000001010010101",
13984 => "0000001010010101",
13985 => "0000001010010101",
13986 => "0000001010010101",
13987 => "0000001010010101",
13988 => "0000001010010110",
13989 => "0000001010010110",
13990 => "0000001010010110",
13991 => "0000001010010110",
13992 => "0000001010010110",
13993 => "0000001010010110",
13994 => "0000001010010110",
13995 => "0000001010010111",
13996 => "0000001010010111",
13997 => "0000001010010111",
13998 => "0000001010010111",
13999 => "0000001010010111",
14000 => "0000001010010111",
14001 => "0000001010011000",
14002 => "0000001010011000",
14003 => "0000001010011000",
14004 => "0000001010011000",
14005 => "0000001010011000",
14006 => "0000001010011000",
14007 => "0000001010011001",
14008 => "0000001010011001",
14009 => "0000001010011001",
14010 => "0000001010011001",
14011 => "0000001010011001",
14012 => "0000001010011001",
14013 => "0000001010011010",
14014 => "0000001010011010",
14015 => "0000001010011010",
14016 => "0000001010011010",
14017 => "0000001010011010",
14018 => "0000001010011010",
14019 => "0000001010011010",
14020 => "0000001010011011",
14021 => "0000001010011011",
14022 => "0000001010011011",
14023 => "0000001010011011",
14024 => "0000001010011011",
14025 => "0000001010011011",
14026 => "0000001010011100",
14027 => "0000001010011100",
14028 => "0000001010011100",
14029 => "0000001010011100",
14030 => "0000001010011100",
14031 => "0000001010011100",
14032 => "0000001010011101",
14033 => "0000001010011101",
14034 => "0000001010011101",
14035 => "0000001010011101",
14036 => "0000001010011101",
14037 => "0000001010011101",
14038 => "0000001010011110",
14039 => "0000001010011110",
14040 => "0000001010011110",
14041 => "0000001010011110",
14042 => "0000001010011110",
14043 => "0000001010011110",
14044 => "0000001010011111",
14045 => "0000001010011111",
14046 => "0000001010011111",
14047 => "0000001010011111",
14048 => "0000001010011111",
14049 => "0000001010011111",
14050 => "0000001010100000",
14051 => "0000001010100000",
14052 => "0000001010100000",
14053 => "0000001010100000",
14054 => "0000001010100000",
14055 => "0000001010100000",
14056 => "0000001010100000",
14057 => "0000001010100001",
14058 => "0000001010100001",
14059 => "0000001010100001",
14060 => "0000001010100001",
14061 => "0000001010100001",
14062 => "0000001010100001",
14063 => "0000001010100010",
14064 => "0000001010100010",
14065 => "0000001010100010",
14066 => "0000001010100010",
14067 => "0000001010100010",
14068 => "0000001010100010",
14069 => "0000001010100011",
14070 => "0000001010100011",
14071 => "0000001010100011",
14072 => "0000001010100011",
14073 => "0000001010100011",
14074 => "0000001010100011",
14075 => "0000001010100100",
14076 => "0000001010100100",
14077 => "0000001010100100",
14078 => "0000001010100100",
14079 => "0000001010100100",
14080 => "0000001010100100",
14081 => "0000001010100101",
14082 => "0000001010100101",
14083 => "0000001010100101",
14084 => "0000001010100101",
14085 => "0000001010100101",
14086 => "0000001010100101",
14087 => "0000001010100110",
14088 => "0000001010100110",
14089 => "0000001010100110",
14090 => "0000001010100110",
14091 => "0000001010100110",
14092 => "0000001010100110",
14093 => "0000001010100111",
14094 => "0000001010100111",
14095 => "0000001010100111",
14096 => "0000001010100111",
14097 => "0000001010100111",
14098 => "0000001010100111",
14099 => "0000001010101000",
14100 => "0000001010101000",
14101 => "0000001010101000",
14102 => "0000001010101000",
14103 => "0000001010101000",
14104 => "0000001010101000",
14105 => "0000001010101001",
14106 => "0000001010101001",
14107 => "0000001010101001",
14108 => "0000001010101001",
14109 => "0000001010101001",
14110 => "0000001010101001",
14111 => "0000001010101001",
14112 => "0000001010101010",
14113 => "0000001010101010",
14114 => "0000001010101010",
14115 => "0000001010101010",
14116 => "0000001010101010",
14117 => "0000001010101010",
14118 => "0000001010101011",
14119 => "0000001010101011",
14120 => "0000001010101011",
14121 => "0000001010101011",
14122 => "0000001010101011",
14123 => "0000001010101011",
14124 => "0000001010101100",
14125 => "0000001010101100",
14126 => "0000001010101100",
14127 => "0000001010101100",
14128 => "0000001010101100",
14129 => "0000001010101100",
14130 => "0000001010101101",
14131 => "0000001010101101",
14132 => "0000001010101101",
14133 => "0000001010101101",
14134 => "0000001010101101",
14135 => "0000001010101101",
14136 => "0000001010101110",
14137 => "0000001010101110",
14138 => "0000001010101110",
14139 => "0000001010101110",
14140 => "0000001010101110",
14141 => "0000001010101110",
14142 => "0000001010101111",
14143 => "0000001010101111",
14144 => "0000001010101111",
14145 => "0000001010101111",
14146 => "0000001010101111",
14147 => "0000001010101111",
14148 => "0000001010110000",
14149 => "0000001010110000",
14150 => "0000001010110000",
14151 => "0000001010110000",
14152 => "0000001010110000",
14153 => "0000001010110000",
14154 => "0000001010110001",
14155 => "0000001010110001",
14156 => "0000001010110001",
14157 => "0000001010110001",
14158 => "0000001010110001",
14159 => "0000001010110001",
14160 => "0000001010110010",
14161 => "0000001010110010",
14162 => "0000001010110010",
14163 => "0000001010110010",
14164 => "0000001010110010",
14165 => "0000001010110010",
14166 => "0000001010110011",
14167 => "0000001010110011",
14168 => "0000001010110011",
14169 => "0000001010110011",
14170 => "0000001010110011",
14171 => "0000001010110011",
14172 => "0000001010110100",
14173 => "0000001010110100",
14174 => "0000001010110100",
14175 => "0000001010110100",
14176 => "0000001010110100",
14177 => "0000001010110100",
14178 => "0000001010110101",
14179 => "0000001010110101",
14180 => "0000001010110101",
14181 => "0000001010110101",
14182 => "0000001010110101",
14183 => "0000001010110101",
14184 => "0000001010110110",
14185 => "0000001010110110",
14186 => "0000001010110110",
14187 => "0000001010110110",
14188 => "0000001010110110",
14189 => "0000001010110110",
14190 => "0000001010110111",
14191 => "0000001010110111",
14192 => "0000001010110111",
14193 => "0000001010110111",
14194 => "0000001010110111",
14195 => "0000001010110111",
14196 => "0000001010111000",
14197 => "0000001010111000",
14198 => "0000001010111000",
14199 => "0000001010111000",
14200 => "0000001010111000",
14201 => "0000001010111000",
14202 => "0000001010111001",
14203 => "0000001010111001",
14204 => "0000001010111001",
14205 => "0000001010111001",
14206 => "0000001010111001",
14207 => "0000001010111001",
14208 => "0000001010111010",
14209 => "0000001010111010",
14210 => "0000001010111010",
14211 => "0000001010111010",
14212 => "0000001010111010",
14213 => "0000001010111011",
14214 => "0000001010111011",
14215 => "0000001010111011",
14216 => "0000001010111011",
14217 => "0000001010111011",
14218 => "0000001010111011",
14219 => "0000001010111100",
14220 => "0000001010111100",
14221 => "0000001010111100",
14222 => "0000001010111100",
14223 => "0000001010111100",
14224 => "0000001010111100",
14225 => "0000001010111101",
14226 => "0000001010111101",
14227 => "0000001010111101",
14228 => "0000001010111101",
14229 => "0000001010111101",
14230 => "0000001010111101",
14231 => "0000001010111110",
14232 => "0000001010111110",
14233 => "0000001010111110",
14234 => "0000001010111110",
14235 => "0000001010111110",
14236 => "0000001010111110",
14237 => "0000001010111111",
14238 => "0000001010111111",
14239 => "0000001010111111",
14240 => "0000001010111111",
14241 => "0000001010111111",
14242 => "0000001010111111",
14243 => "0000001011000000",
14244 => "0000001011000000",
14245 => "0000001011000000",
14246 => "0000001011000000",
14247 => "0000001011000000",
14248 => "0000001011000000",
14249 => "0000001011000001",
14250 => "0000001011000001",
14251 => "0000001011000001",
14252 => "0000001011000001",
14253 => "0000001011000001",
14254 => "0000001011000001",
14255 => "0000001011000010",
14256 => "0000001011000010",
14257 => "0000001011000010",
14258 => "0000001011000010",
14259 => "0000001011000010",
14260 => "0000001011000010",
14261 => "0000001011000011",
14262 => "0000001011000011",
14263 => "0000001011000011",
14264 => "0000001011000011",
14265 => "0000001011000011",
14266 => "0000001011000100",
14267 => "0000001011000100",
14268 => "0000001011000100",
14269 => "0000001011000100",
14270 => "0000001011000100",
14271 => "0000001011000100",
14272 => "0000001011000101",
14273 => "0000001011000101",
14274 => "0000001011000101",
14275 => "0000001011000101",
14276 => "0000001011000101",
14277 => "0000001011000101",
14278 => "0000001011000110",
14279 => "0000001011000110",
14280 => "0000001011000110",
14281 => "0000001011000110",
14282 => "0000001011000110",
14283 => "0000001011000110",
14284 => "0000001011000111",
14285 => "0000001011000111",
14286 => "0000001011000111",
14287 => "0000001011000111",
14288 => "0000001011000111",
14289 => "0000001011000111",
14290 => "0000001011001000",
14291 => "0000001011001000",
14292 => "0000001011001000",
14293 => "0000001011001000",
14294 => "0000001011001000",
14295 => "0000001011001000",
14296 => "0000001011001001",
14297 => "0000001011001001",
14298 => "0000001011001001",
14299 => "0000001011001001",
14300 => "0000001011001001",
14301 => "0000001011001010",
14302 => "0000001011001010",
14303 => "0000001011001010",
14304 => "0000001011001010",
14305 => "0000001011001010",
14306 => "0000001011001010",
14307 => "0000001011001011",
14308 => "0000001011001011",
14309 => "0000001011001011",
14310 => "0000001011001011",
14311 => "0000001011001011",
14312 => "0000001011001011",
14313 => "0000001011001100",
14314 => "0000001011001100",
14315 => "0000001011001100",
14316 => "0000001011001100",
14317 => "0000001011001100",
14318 => "0000001011001100",
14319 => "0000001011001101",
14320 => "0000001011001101",
14321 => "0000001011001101",
14322 => "0000001011001101",
14323 => "0000001011001101",
14324 => "0000001011001101",
14325 => "0000001011001110",
14326 => "0000001011001110",
14327 => "0000001011001110",
14328 => "0000001011001110",
14329 => "0000001011001110",
14330 => "0000001011001111",
14331 => "0000001011001111",
14332 => "0000001011001111",
14333 => "0000001011001111",
14334 => "0000001011001111",
14335 => "0000001011001111",
14336 => "0000001011010000",
14337 => "0000001011010000",
14338 => "0000001011010000",
14339 => "0000001011010000",
14340 => "0000001011010000",
14341 => "0000001011010000",
14342 => "0000001011010001",
14343 => "0000001011010001",
14344 => "0000001011010001",
14345 => "0000001011010001",
14346 => "0000001011010001",
14347 => "0000001011010001",
14348 => "0000001011010010",
14349 => "0000001011010010",
14350 => "0000001011010010",
14351 => "0000001011010010",
14352 => "0000001011010010",
14353 => "0000001011010011",
14354 => "0000001011010011",
14355 => "0000001011010011",
14356 => "0000001011010011",
14357 => "0000001011010011",
14358 => "0000001011010011",
14359 => "0000001011010100",
14360 => "0000001011010100",
14361 => "0000001011010100",
14362 => "0000001011010100",
14363 => "0000001011010100",
14364 => "0000001011010100",
14365 => "0000001011010101",
14366 => "0000001011010101",
14367 => "0000001011010101",
14368 => "0000001011010101",
14369 => "0000001011010101",
14370 => "0000001011010110",
14371 => "0000001011010110",
14372 => "0000001011010110",
14373 => "0000001011010110",
14374 => "0000001011010110",
14375 => "0000001011010110",
14376 => "0000001011010111",
14377 => "0000001011010111",
14378 => "0000001011010111",
14379 => "0000001011010111",
14380 => "0000001011010111",
14381 => "0000001011010111",
14382 => "0000001011011000",
14383 => "0000001011011000",
14384 => "0000001011011000",
14385 => "0000001011011000",
14386 => "0000001011011000",
14387 => "0000001011011000",
14388 => "0000001011011001",
14389 => "0000001011011001",
14390 => "0000001011011001",
14391 => "0000001011011001",
14392 => "0000001011011001",
14393 => "0000001011011010",
14394 => "0000001011011010",
14395 => "0000001011011010",
14396 => "0000001011011010",
14397 => "0000001011011010",
14398 => "0000001011011010",
14399 => "0000001011011011",
14400 => "0000001011011011",
14401 => "0000001011011011",
14402 => "0000001011011011",
14403 => "0000001011011011",
14404 => "0000001011011011",
14405 => "0000001011011100",
14406 => "0000001011011100",
14407 => "0000001011011100",
14408 => "0000001011011100",
14409 => "0000001011011100",
14410 => "0000001011011101",
14411 => "0000001011011101",
14412 => "0000001011011101",
14413 => "0000001011011101",
14414 => "0000001011011101",
14415 => "0000001011011101",
14416 => "0000001011011110",
14417 => "0000001011011110",
14418 => "0000001011011110",
14419 => "0000001011011110",
14420 => "0000001011011110",
14421 => "0000001011011111",
14422 => "0000001011011111",
14423 => "0000001011011111",
14424 => "0000001011011111",
14425 => "0000001011011111",
14426 => "0000001011011111",
14427 => "0000001011100000",
14428 => "0000001011100000",
14429 => "0000001011100000",
14430 => "0000001011100000",
14431 => "0000001011100000",
14432 => "0000001011100000",
14433 => "0000001011100001",
14434 => "0000001011100001",
14435 => "0000001011100001",
14436 => "0000001011100001",
14437 => "0000001011100001",
14438 => "0000001011100010",
14439 => "0000001011100010",
14440 => "0000001011100010",
14441 => "0000001011100010",
14442 => "0000001011100010",
14443 => "0000001011100010",
14444 => "0000001011100011",
14445 => "0000001011100011",
14446 => "0000001011100011",
14447 => "0000001011100011",
14448 => "0000001011100011",
14449 => "0000001011100011",
14450 => "0000001011100100",
14451 => "0000001011100100",
14452 => "0000001011100100",
14453 => "0000001011100100",
14454 => "0000001011100100",
14455 => "0000001011100101",
14456 => "0000001011100101",
14457 => "0000001011100101",
14458 => "0000001011100101",
14459 => "0000001011100101",
14460 => "0000001011100101",
14461 => "0000001011100110",
14462 => "0000001011100110",
14463 => "0000001011100110",
14464 => "0000001011100110",
14465 => "0000001011100110",
14466 => "0000001011100111",
14467 => "0000001011100111",
14468 => "0000001011100111",
14469 => "0000001011100111",
14470 => "0000001011100111",
14471 => "0000001011100111",
14472 => "0000001011101000",
14473 => "0000001011101000",
14474 => "0000001011101000",
14475 => "0000001011101000",
14476 => "0000001011101000",
14477 => "0000001011101001",
14478 => "0000001011101001",
14479 => "0000001011101001",
14480 => "0000001011101001",
14481 => "0000001011101001",
14482 => "0000001011101001",
14483 => "0000001011101010",
14484 => "0000001011101010",
14485 => "0000001011101010",
14486 => "0000001011101010",
14487 => "0000001011101010",
14488 => "0000001011101010",
14489 => "0000001011101011",
14490 => "0000001011101011",
14491 => "0000001011101011",
14492 => "0000001011101011",
14493 => "0000001011101011",
14494 => "0000001011101100",
14495 => "0000001011101100",
14496 => "0000001011101100",
14497 => "0000001011101100",
14498 => "0000001011101100",
14499 => "0000001011101100",
14500 => "0000001011101101",
14501 => "0000001011101101",
14502 => "0000001011101101",
14503 => "0000001011101101",
14504 => "0000001011101101",
14505 => "0000001011101110",
14506 => "0000001011101110",
14507 => "0000001011101110",
14508 => "0000001011101110",
14509 => "0000001011101110",
14510 => "0000001011101110",
14511 => "0000001011101111",
14512 => "0000001011101111",
14513 => "0000001011101111",
14514 => "0000001011101111",
14515 => "0000001011101111",
14516 => "0000001011110000",
14517 => "0000001011110000",
14518 => "0000001011110000",
14519 => "0000001011110000",
14520 => "0000001011110000",
14521 => "0000001011110000",
14522 => "0000001011110001",
14523 => "0000001011110001",
14524 => "0000001011110001",
14525 => "0000001011110001",
14526 => "0000001011110001",
14527 => "0000001011110010",
14528 => "0000001011110010",
14529 => "0000001011110010",
14530 => "0000001011110010",
14531 => "0000001011110010",
14532 => "0000001011110010",
14533 => "0000001011110011",
14534 => "0000001011110011",
14535 => "0000001011110011",
14536 => "0000001011110011",
14537 => "0000001011110011",
14538 => "0000001011110100",
14539 => "0000001011110100",
14540 => "0000001011110100",
14541 => "0000001011110100",
14542 => "0000001011110100",
14543 => "0000001011110100",
14544 => "0000001011110101",
14545 => "0000001011110101",
14546 => "0000001011110101",
14547 => "0000001011110101",
14548 => "0000001011110101",
14549 => "0000001011110110",
14550 => "0000001011110110",
14551 => "0000001011110110",
14552 => "0000001011110110",
14553 => "0000001011110110",
14554 => "0000001011110110",
14555 => "0000001011110111",
14556 => "0000001011110111",
14557 => "0000001011110111",
14558 => "0000001011110111",
14559 => "0000001011110111",
14560 => "0000001011111000",
14561 => "0000001011111000",
14562 => "0000001011111000",
14563 => "0000001011111000",
14564 => "0000001011111000",
14565 => "0000001011111001",
14566 => "0000001011111001",
14567 => "0000001011111001",
14568 => "0000001011111001",
14569 => "0000001011111001",
14570 => "0000001011111001",
14571 => "0000001011111010",
14572 => "0000001011111010",
14573 => "0000001011111010",
14574 => "0000001011111010",
14575 => "0000001011111010",
14576 => "0000001011111011",
14577 => "0000001011111011",
14578 => "0000001011111011",
14579 => "0000001011111011",
14580 => "0000001011111011",
14581 => "0000001011111011",
14582 => "0000001011111100",
14583 => "0000001011111100",
14584 => "0000001011111100",
14585 => "0000001011111100",
14586 => "0000001011111100",
14587 => "0000001011111101",
14588 => "0000001011111101",
14589 => "0000001011111101",
14590 => "0000001011111101",
14591 => "0000001011111101",
14592 => "0000001011111101",
14593 => "0000001011111110",
14594 => "0000001011111110",
14595 => "0000001011111110",
14596 => "0000001011111110",
14597 => "0000001011111110",
14598 => "0000001011111111",
14599 => "0000001011111111",
14600 => "0000001011111111",
14601 => "0000001011111111",
14602 => "0000001011111111",
14603 => "0000001100000000",
14604 => "0000001100000000",
14605 => "0000001100000000",
14606 => "0000001100000000",
14607 => "0000001100000000",
14608 => "0000001100000000",
14609 => "0000001100000001",
14610 => "0000001100000001",
14611 => "0000001100000001",
14612 => "0000001100000001",
14613 => "0000001100000001",
14614 => "0000001100000010",
14615 => "0000001100000010",
14616 => "0000001100000010",
14617 => "0000001100000010",
14618 => "0000001100000010",
14619 => "0000001100000010",
14620 => "0000001100000011",
14621 => "0000001100000011",
14622 => "0000001100000011",
14623 => "0000001100000011",
14624 => "0000001100000011",
14625 => "0000001100000100",
14626 => "0000001100000100",
14627 => "0000001100000100",
14628 => "0000001100000100",
14629 => "0000001100000100",
14630 => "0000001100000101",
14631 => "0000001100000101",
14632 => "0000001100000101",
14633 => "0000001100000101",
14634 => "0000001100000101",
14635 => "0000001100000101",
14636 => "0000001100000110",
14637 => "0000001100000110",
14638 => "0000001100000110",
14639 => "0000001100000110",
14640 => "0000001100000110",
14641 => "0000001100000111",
14642 => "0000001100000111",
14643 => "0000001100000111",
14644 => "0000001100000111",
14645 => "0000001100000111",
14646 => "0000001100001000",
14647 => "0000001100001000",
14648 => "0000001100001000",
14649 => "0000001100001000",
14650 => "0000001100001000",
14651 => "0000001100001000",
14652 => "0000001100001001",
14653 => "0000001100001001",
14654 => "0000001100001001",
14655 => "0000001100001001",
14656 => "0000001100001001",
14657 => "0000001100001010",
14658 => "0000001100001010",
14659 => "0000001100001010",
14660 => "0000001100001010",
14661 => "0000001100001010",
14662 => "0000001100001011",
14663 => "0000001100001011",
14664 => "0000001100001011",
14665 => "0000001100001011",
14666 => "0000001100001011",
14667 => "0000001100001011",
14668 => "0000001100001100",
14669 => "0000001100001100",
14670 => "0000001100001100",
14671 => "0000001100001100",
14672 => "0000001100001100",
14673 => "0000001100001101",
14674 => "0000001100001101",
14675 => "0000001100001101",
14676 => "0000001100001101",
14677 => "0000001100001101",
14678 => "0000001100001110",
14679 => "0000001100001110",
14680 => "0000001100001110",
14681 => "0000001100001110",
14682 => "0000001100001110",
14683 => "0000001100001110",
14684 => "0000001100001111",
14685 => "0000001100001111",
14686 => "0000001100001111",
14687 => "0000001100001111",
14688 => "0000001100001111",
14689 => "0000001100010000",
14690 => "0000001100010000",
14691 => "0000001100010000",
14692 => "0000001100010000",
14693 => "0000001100010000",
14694 => "0000001100010001",
14695 => "0000001100010001",
14696 => "0000001100010001",
14697 => "0000001100010001",
14698 => "0000001100010001",
14699 => "0000001100010010",
14700 => "0000001100010010",
14701 => "0000001100010010",
14702 => "0000001100010010",
14703 => "0000001100010010",
14704 => "0000001100010010",
14705 => "0000001100010011",
14706 => "0000001100010011",
14707 => "0000001100010011",
14708 => "0000001100010011",
14709 => "0000001100010011",
14710 => "0000001100010100",
14711 => "0000001100010100",
14712 => "0000001100010100",
14713 => "0000001100010100",
14714 => "0000001100010100",
14715 => "0000001100010101",
14716 => "0000001100010101",
14717 => "0000001100010101",
14718 => "0000001100010101",
14719 => "0000001100010101",
14720 => "0000001100010101",
14721 => "0000001100010110",
14722 => "0000001100010110",
14723 => "0000001100010110",
14724 => "0000001100010110",
14725 => "0000001100010110",
14726 => "0000001100010111",
14727 => "0000001100010111",
14728 => "0000001100010111",
14729 => "0000001100010111",
14730 => "0000001100010111",
14731 => "0000001100011000",
14732 => "0000001100011000",
14733 => "0000001100011000",
14734 => "0000001100011000",
14735 => "0000001100011000",
14736 => "0000001100011001",
14737 => "0000001100011001",
14738 => "0000001100011001",
14739 => "0000001100011001",
14740 => "0000001100011001",
14741 => "0000001100011010",
14742 => "0000001100011010",
14743 => "0000001100011010",
14744 => "0000001100011010",
14745 => "0000001100011010",
14746 => "0000001100011010",
14747 => "0000001100011011",
14748 => "0000001100011011",
14749 => "0000001100011011",
14750 => "0000001100011011",
14751 => "0000001100011011",
14752 => "0000001100011100",
14753 => "0000001100011100",
14754 => "0000001100011100",
14755 => "0000001100011100",
14756 => "0000001100011100",
14757 => "0000001100011101",
14758 => "0000001100011101",
14759 => "0000001100011101",
14760 => "0000001100011101",
14761 => "0000001100011101",
14762 => "0000001100011110",
14763 => "0000001100011110",
14764 => "0000001100011110",
14765 => "0000001100011110",
14766 => "0000001100011110",
14767 => "0000001100011111",
14768 => "0000001100011111",
14769 => "0000001100011111",
14770 => "0000001100011111",
14771 => "0000001100011111",
14772 => "0000001100011111",
14773 => "0000001100100000",
14774 => "0000001100100000",
14775 => "0000001100100000",
14776 => "0000001100100000",
14777 => "0000001100100000",
14778 => "0000001100100001",
14779 => "0000001100100001",
14780 => "0000001100100001",
14781 => "0000001100100001",
14782 => "0000001100100001",
14783 => "0000001100100010",
14784 => "0000001100100010",
14785 => "0000001100100010",
14786 => "0000001100100010",
14787 => "0000001100100010",
14788 => "0000001100100011",
14789 => "0000001100100011",
14790 => "0000001100100011",
14791 => "0000001100100011",
14792 => "0000001100100011",
14793 => "0000001100100100",
14794 => "0000001100100100",
14795 => "0000001100100100",
14796 => "0000001100100100",
14797 => "0000001100100100",
14798 => "0000001100100101",
14799 => "0000001100100101",
14800 => "0000001100100101",
14801 => "0000001100100101",
14802 => "0000001100100101",
14803 => "0000001100100101",
14804 => "0000001100100110",
14805 => "0000001100100110",
14806 => "0000001100100110",
14807 => "0000001100100110",
14808 => "0000001100100110",
14809 => "0000001100100111",
14810 => "0000001100100111",
14811 => "0000001100100111",
14812 => "0000001100100111",
14813 => "0000001100100111",
14814 => "0000001100101000",
14815 => "0000001100101000",
14816 => "0000001100101000",
14817 => "0000001100101000",
14818 => "0000001100101000",
14819 => "0000001100101001",
14820 => "0000001100101001",
14821 => "0000001100101001",
14822 => "0000001100101001",
14823 => "0000001100101001",
14824 => "0000001100101010",
14825 => "0000001100101010",
14826 => "0000001100101010",
14827 => "0000001100101010",
14828 => "0000001100101010",
14829 => "0000001100101011",
14830 => "0000001100101011",
14831 => "0000001100101011",
14832 => "0000001100101011",
14833 => "0000001100101011",
14834 => "0000001100101100",
14835 => "0000001100101100",
14836 => "0000001100101100",
14837 => "0000001100101100",
14838 => "0000001100101100",
14839 => "0000001100101100",
14840 => "0000001100101101",
14841 => "0000001100101101",
14842 => "0000001100101101",
14843 => "0000001100101101",
14844 => "0000001100101101",
14845 => "0000001100101110",
14846 => "0000001100101110",
14847 => "0000001100101110",
14848 => "0000001100101110",
14849 => "0000001100101110",
14850 => "0000001100101111",
14851 => "0000001100101111",
14852 => "0000001100101111",
14853 => "0000001100101111",
14854 => "0000001100101111",
14855 => "0000001100110000",
14856 => "0000001100110000",
14857 => "0000001100110000",
14858 => "0000001100110000",
14859 => "0000001100110000",
14860 => "0000001100110001",
14861 => "0000001100110001",
14862 => "0000001100110001",
14863 => "0000001100110001",
14864 => "0000001100110001",
14865 => "0000001100110010",
14866 => "0000001100110010",
14867 => "0000001100110010",
14868 => "0000001100110010",
14869 => "0000001100110010",
14870 => "0000001100110011",
14871 => "0000001100110011",
14872 => "0000001100110011",
14873 => "0000001100110011",
14874 => "0000001100110011",
14875 => "0000001100110100",
14876 => "0000001100110100",
14877 => "0000001100110100",
14878 => "0000001100110100",
14879 => "0000001100110100",
14880 => "0000001100110101",
14881 => "0000001100110101",
14882 => "0000001100110101",
14883 => "0000001100110101",
14884 => "0000001100110101",
14885 => "0000001100110110",
14886 => "0000001100110110",
14887 => "0000001100110110",
14888 => "0000001100110110",
14889 => "0000001100110110",
14890 => "0000001100110111",
14891 => "0000001100110111",
14892 => "0000001100110111",
14893 => "0000001100110111",
14894 => "0000001100110111",
14895 => "0000001100111000",
14896 => "0000001100111000",
14897 => "0000001100111000",
14898 => "0000001100111000",
14899 => "0000001100111000",
14900 => "0000001100111001",
14901 => "0000001100111001",
14902 => "0000001100111001",
14903 => "0000001100111001",
14904 => "0000001100111001",
14905 => "0000001100111010",
14906 => "0000001100111010",
14907 => "0000001100111010",
14908 => "0000001100111010",
14909 => "0000001100111010",
14910 => "0000001100111011",
14911 => "0000001100111011",
14912 => "0000001100111011",
14913 => "0000001100111011",
14914 => "0000001100111011",
14915 => "0000001100111100",
14916 => "0000001100111100",
14917 => "0000001100111100",
14918 => "0000001100111100",
14919 => "0000001100111100",
14920 => "0000001100111101",
14921 => "0000001100111101",
14922 => "0000001100111101",
14923 => "0000001100111101",
14924 => "0000001100111101",
14925 => "0000001100111110",
14926 => "0000001100111110",
14927 => "0000001100111110",
14928 => "0000001100111110",
14929 => "0000001100111110",
14930 => "0000001100111111",
14931 => "0000001100111111",
14932 => "0000001100111111",
14933 => "0000001100111111",
14934 => "0000001100111111",
14935 => "0000001101000000",
14936 => "0000001101000000",
14937 => "0000001101000000",
14938 => "0000001101000000",
14939 => "0000001101000000",
14940 => "0000001101000001",
14941 => "0000001101000001",
14942 => "0000001101000001",
14943 => "0000001101000001",
14944 => "0000001101000001",
14945 => "0000001101000010",
14946 => "0000001101000010",
14947 => "0000001101000010",
14948 => "0000001101000010",
14949 => "0000001101000010",
14950 => "0000001101000011",
14951 => "0000001101000011",
14952 => "0000001101000011",
14953 => "0000001101000011",
14954 => "0000001101000011",
14955 => "0000001101000100",
14956 => "0000001101000100",
14957 => "0000001101000100",
14958 => "0000001101000100",
14959 => "0000001101000100",
14960 => "0000001101000101",
14961 => "0000001101000101",
14962 => "0000001101000101",
14963 => "0000001101000101",
14964 => "0000001101000101",
14965 => "0000001101000110",
14966 => "0000001101000110",
14967 => "0000001101000110",
14968 => "0000001101000110",
14969 => "0000001101000110",
14970 => "0000001101000111",
14971 => "0000001101000111",
14972 => "0000001101000111",
14973 => "0000001101000111",
14974 => "0000001101000111",
14975 => "0000001101001000",
14976 => "0000001101001000",
14977 => "0000001101001000",
14978 => "0000001101001000",
14979 => "0000001101001000",
14980 => "0000001101001001",
14981 => "0000001101001001",
14982 => "0000001101001001",
14983 => "0000001101001001",
14984 => "0000001101001001",
14985 => "0000001101001010",
14986 => "0000001101001010",
14987 => "0000001101001010",
14988 => "0000001101001010",
14989 => "0000001101001010",
14990 => "0000001101001011",
14991 => "0000001101001011",
14992 => "0000001101001011",
14993 => "0000001101001011",
14994 => "0000001101001011",
14995 => "0000001101001100",
14996 => "0000001101001100",
14997 => "0000001101001100",
14998 => "0000001101001100",
14999 => "0000001101001100",
15000 => "0000001101001101",
15001 => "0000001101001101",
15002 => "0000001101001101",
15003 => "0000001101001101",
15004 => "0000001101001101",
15005 => "0000001101001110",
15006 => "0000001101001110",
15007 => "0000001101001110",
15008 => "0000001101001110",
15009 => "0000001101001111",
15010 => "0000001101001111",
15011 => "0000001101001111",
15012 => "0000001101001111",
15013 => "0000001101001111",
15014 => "0000001101010000",
15015 => "0000001101010000",
15016 => "0000001101010000",
15017 => "0000001101010000",
15018 => "0000001101010000",
15019 => "0000001101010001",
15020 => "0000001101010001",
15021 => "0000001101010001",
15022 => "0000001101010001",
15023 => "0000001101010001",
15024 => "0000001101010010",
15025 => "0000001101010010",
15026 => "0000001101010010",
15027 => "0000001101010010",
15028 => "0000001101010010",
15029 => "0000001101010011",
15030 => "0000001101010011",
15031 => "0000001101010011",
15032 => "0000001101010011",
15033 => "0000001101010011",
15034 => "0000001101010100",
15035 => "0000001101010100",
15036 => "0000001101010100",
15037 => "0000001101010100",
15038 => "0000001101010100",
15039 => "0000001101010101",
15040 => "0000001101010101",
15041 => "0000001101010101",
15042 => "0000001101010101",
15043 => "0000001101010101",
15044 => "0000001101010110",
15045 => "0000001101010110",
15046 => "0000001101010110",
15047 => "0000001101010110",
15048 => "0000001101010111",
15049 => "0000001101010111",
15050 => "0000001101010111",
15051 => "0000001101010111",
15052 => "0000001101010111",
15053 => "0000001101011000",
15054 => "0000001101011000",
15055 => "0000001101011000",
15056 => "0000001101011000",
15057 => "0000001101011000",
15058 => "0000001101011001",
15059 => "0000001101011001",
15060 => "0000001101011001",
15061 => "0000001101011001",
15062 => "0000001101011001",
15063 => "0000001101011010",
15064 => "0000001101011010",
15065 => "0000001101011010",
15066 => "0000001101011010",
15067 => "0000001101011010",
15068 => "0000001101011011",
15069 => "0000001101011011",
15070 => "0000001101011011",
15071 => "0000001101011011",
15072 => "0000001101011011",
15073 => "0000001101011100",
15074 => "0000001101011100",
15075 => "0000001101011100",
15076 => "0000001101011100",
15077 => "0000001101011100",
15078 => "0000001101011101",
15079 => "0000001101011101",
15080 => "0000001101011101",
15081 => "0000001101011101",
15082 => "0000001101011110",
15083 => "0000001101011110",
15084 => "0000001101011110",
15085 => "0000001101011110",
15086 => "0000001101011110",
15087 => "0000001101011111",
15088 => "0000001101011111",
15089 => "0000001101011111",
15090 => "0000001101011111",
15091 => "0000001101011111",
15092 => "0000001101100000",
15093 => "0000001101100000",
15094 => "0000001101100000",
15095 => "0000001101100000",
15096 => "0000001101100000",
15097 => "0000001101100001",
15098 => "0000001101100001",
15099 => "0000001101100001",
15100 => "0000001101100001",
15101 => "0000001101100001",
15102 => "0000001101100010",
15103 => "0000001101100010",
15104 => "0000001101100010",
15105 => "0000001101100010",
15106 => "0000001101100011",
15107 => "0000001101100011",
15108 => "0000001101100011",
15109 => "0000001101100011",
15110 => "0000001101100011",
15111 => "0000001101100100",
15112 => "0000001101100100",
15113 => "0000001101100100",
15114 => "0000001101100100",
15115 => "0000001101100100",
15116 => "0000001101100101",
15117 => "0000001101100101",
15118 => "0000001101100101",
15119 => "0000001101100101",
15120 => "0000001101100101",
15121 => "0000001101100110",
15122 => "0000001101100110",
15123 => "0000001101100110",
15124 => "0000001101100110",
15125 => "0000001101100111",
15126 => "0000001101100111",
15127 => "0000001101100111",
15128 => "0000001101100111",
15129 => "0000001101100111",
15130 => "0000001101101000",
15131 => "0000001101101000",
15132 => "0000001101101000",
15133 => "0000001101101000",
15134 => "0000001101101000",
15135 => "0000001101101001",
15136 => "0000001101101001",
15137 => "0000001101101001",
15138 => "0000001101101001",
15139 => "0000001101101001",
15140 => "0000001101101010",
15141 => "0000001101101010",
15142 => "0000001101101010",
15143 => "0000001101101010",
15144 => "0000001101101011",
15145 => "0000001101101011",
15146 => "0000001101101011",
15147 => "0000001101101011",
15148 => "0000001101101011",
15149 => "0000001101101100",
15150 => "0000001101101100",
15151 => "0000001101101100",
15152 => "0000001101101100",
15153 => "0000001101101100",
15154 => "0000001101101101",
15155 => "0000001101101101",
15156 => "0000001101101101",
15157 => "0000001101101101",
15158 => "0000001101101101",
15159 => "0000001101101110",
15160 => "0000001101101110",
15161 => "0000001101101110",
15162 => "0000001101101110",
15163 => "0000001101101111",
15164 => "0000001101101111",
15165 => "0000001101101111",
15166 => "0000001101101111",
15167 => "0000001101101111",
15168 => "0000001101110000",
15169 => "0000001101110000",
15170 => "0000001101110000",
15171 => "0000001101110000",
15172 => "0000001101110000",
15173 => "0000001101110001",
15174 => "0000001101110001",
15175 => "0000001101110001",
15176 => "0000001101110001",
15177 => "0000001101110001",
15178 => "0000001101110010",
15179 => "0000001101110010",
15180 => "0000001101110010",
15181 => "0000001101110010",
15182 => "0000001101110011",
15183 => "0000001101110011",
15184 => "0000001101110011",
15185 => "0000001101110011",
15186 => "0000001101110011",
15187 => "0000001101110100",
15188 => "0000001101110100",
15189 => "0000001101110100",
15190 => "0000001101110100",
15191 => "0000001101110100",
15192 => "0000001101110101",
15193 => "0000001101110101",
15194 => "0000001101110101",
15195 => "0000001101110101",
15196 => "0000001101110110",
15197 => "0000001101110110",
15198 => "0000001101110110",
15199 => "0000001101110110",
15200 => "0000001101110110",
15201 => "0000001101110111",
15202 => "0000001101110111",
15203 => "0000001101110111",
15204 => "0000001101110111",
15205 => "0000001101110111",
15206 => "0000001101111000",
15207 => "0000001101111000",
15208 => "0000001101111000",
15209 => "0000001101111000",
15210 => "0000001101111001",
15211 => "0000001101111001",
15212 => "0000001101111001",
15213 => "0000001101111001",
15214 => "0000001101111001",
15215 => "0000001101111010",
15216 => "0000001101111010",
15217 => "0000001101111010",
15218 => "0000001101111010",
15219 => "0000001101111010",
15220 => "0000001101111011",
15221 => "0000001101111011",
15222 => "0000001101111011",
15223 => "0000001101111011",
15224 => "0000001101111100",
15225 => "0000001101111100",
15226 => "0000001101111100",
15227 => "0000001101111100",
15228 => "0000001101111100",
15229 => "0000001101111101",
15230 => "0000001101111101",
15231 => "0000001101111101",
15232 => "0000001101111101",
15233 => "0000001101111101",
15234 => "0000001101111110",
15235 => "0000001101111110",
15236 => "0000001101111110",
15237 => "0000001101111110",
15238 => "0000001101111111",
15239 => "0000001101111111",
15240 => "0000001101111111",
15241 => "0000001101111111",
15242 => "0000001101111111",
15243 => "0000001110000000",
15244 => "0000001110000000",
15245 => "0000001110000000",
15246 => "0000001110000000",
15247 => "0000001110000000",
15248 => "0000001110000001",
15249 => "0000001110000001",
15250 => "0000001110000001",
15251 => "0000001110000001",
15252 => "0000001110000010",
15253 => "0000001110000010",
15254 => "0000001110000010",
15255 => "0000001110000010",
15256 => "0000001110000010",
15257 => "0000001110000011",
15258 => "0000001110000011",
15259 => "0000001110000011",
15260 => "0000001110000011",
15261 => "0000001110000100",
15262 => "0000001110000100",
15263 => "0000001110000100",
15264 => "0000001110000100",
15265 => "0000001110000100",
15266 => "0000001110000101",
15267 => "0000001110000101",
15268 => "0000001110000101",
15269 => "0000001110000101",
15270 => "0000001110000101",
15271 => "0000001110000110",
15272 => "0000001110000110",
15273 => "0000001110000110",
15274 => "0000001110000110",
15275 => "0000001110000111",
15276 => "0000001110000111",
15277 => "0000001110000111",
15278 => "0000001110000111",
15279 => "0000001110000111",
15280 => "0000001110001000",
15281 => "0000001110001000",
15282 => "0000001110001000",
15283 => "0000001110001000",
15284 => "0000001110001001",
15285 => "0000001110001001",
15286 => "0000001110001001",
15287 => "0000001110001001",
15288 => "0000001110001001",
15289 => "0000001110001010",
15290 => "0000001110001010",
15291 => "0000001110001010",
15292 => "0000001110001010",
15293 => "0000001110001010",
15294 => "0000001110001011",
15295 => "0000001110001011",
15296 => "0000001110001011",
15297 => "0000001110001011",
15298 => "0000001110001100",
15299 => "0000001110001100",
15300 => "0000001110001100",
15301 => "0000001110001100",
15302 => "0000001110001100",
15303 => "0000001110001101",
15304 => "0000001110001101",
15305 => "0000001110001101",
15306 => "0000001110001101",
15307 => "0000001110001110",
15308 => "0000001110001110",
15309 => "0000001110001110",
15310 => "0000001110001110",
15311 => "0000001110001110",
15312 => "0000001110001111",
15313 => "0000001110001111",
15314 => "0000001110001111",
15315 => "0000001110001111",
15316 => "0000001110010000",
15317 => "0000001110010000",
15318 => "0000001110010000",
15319 => "0000001110010000",
15320 => "0000001110010000",
15321 => "0000001110010001",
15322 => "0000001110010001",
15323 => "0000001110010001",
15324 => "0000001110010001",
15325 => "0000001110010001",
15326 => "0000001110010010",
15327 => "0000001110010010",
15328 => "0000001110010010",
15329 => "0000001110010010",
15330 => "0000001110010011",
15331 => "0000001110010011",
15332 => "0000001110010011",
15333 => "0000001110010011",
15334 => "0000001110010011",
15335 => "0000001110010100",
15336 => "0000001110010100",
15337 => "0000001110010100",
15338 => "0000001110010100",
15339 => "0000001110010101",
15340 => "0000001110010101",
15341 => "0000001110010101",
15342 => "0000001110010101",
15343 => "0000001110010101",
15344 => "0000001110010110",
15345 => "0000001110010110",
15346 => "0000001110010110",
15347 => "0000001110010110",
15348 => "0000001110010111",
15349 => "0000001110010111",
15350 => "0000001110010111",
15351 => "0000001110010111",
15352 => "0000001110010111",
15353 => "0000001110011000",
15354 => "0000001110011000",
15355 => "0000001110011000",
15356 => "0000001110011000",
15357 => "0000001110011001",
15358 => "0000001110011001",
15359 => "0000001110011001",
15360 => "0000001110011001",
15361 => "0000001110011001",
15362 => "0000001110011010",
15363 => "0000001110011010",
15364 => "0000001110011010",
15365 => "0000001110011010",
15366 => "0000001110011011",
15367 => "0000001110011011",
15368 => "0000001110011011",
15369 => "0000001110011011",
15370 => "0000001110011011",
15371 => "0000001110011100",
15372 => "0000001110011100",
15373 => "0000001110011100",
15374 => "0000001110011100",
15375 => "0000001110011101",
15376 => "0000001110011101",
15377 => "0000001110011101",
15378 => "0000001110011101",
15379 => "0000001110011101",
15380 => "0000001110011110",
15381 => "0000001110011110",
15382 => "0000001110011110",
15383 => "0000001110011110",
15384 => "0000001110011111",
15385 => "0000001110011111",
15386 => "0000001110011111",
15387 => "0000001110011111",
15388 => "0000001110011111",
15389 => "0000001110100000",
15390 => "0000001110100000",
15391 => "0000001110100000",
15392 => "0000001110100000",
15393 => "0000001110100001",
15394 => "0000001110100001",
15395 => "0000001110100001",
15396 => "0000001110100001",
15397 => "0000001110100001",
15398 => "0000001110100010",
15399 => "0000001110100010",
15400 => "0000001110100010",
15401 => "0000001110100010",
15402 => "0000001110100011",
15403 => "0000001110100011",
15404 => "0000001110100011",
15405 => "0000001110100011",
15406 => "0000001110100011",
15407 => "0000001110100100",
15408 => "0000001110100100",
15409 => "0000001110100100",
15410 => "0000001110100100",
15411 => "0000001110100101",
15412 => "0000001110100101",
15413 => "0000001110100101",
15414 => "0000001110100101",
15415 => "0000001110100110",
15416 => "0000001110100110",
15417 => "0000001110100110",
15418 => "0000001110100110",
15419 => "0000001110100110",
15420 => "0000001110100111",
15421 => "0000001110100111",
15422 => "0000001110100111",
15423 => "0000001110100111",
15424 => "0000001110101000",
15425 => "0000001110101000",
15426 => "0000001110101000",
15427 => "0000001110101000",
15428 => "0000001110101000",
15429 => "0000001110101001",
15430 => "0000001110101001",
15431 => "0000001110101001",
15432 => "0000001110101001",
15433 => "0000001110101010",
15434 => "0000001110101010",
15435 => "0000001110101010",
15436 => "0000001110101010",
15437 => "0000001110101010",
15438 => "0000001110101011",
15439 => "0000001110101011",
15440 => "0000001110101011",
15441 => "0000001110101011",
15442 => "0000001110101100",
15443 => "0000001110101100",
15444 => "0000001110101100",
15445 => "0000001110101100",
15446 => "0000001110101101",
15447 => "0000001110101101",
15448 => "0000001110101101",
15449 => "0000001110101101",
15450 => "0000001110101101",
15451 => "0000001110101110",
15452 => "0000001110101110",
15453 => "0000001110101110",
15454 => "0000001110101110",
15455 => "0000001110101111",
15456 => "0000001110101111",
15457 => "0000001110101111",
15458 => "0000001110101111",
15459 => "0000001110101111",
15460 => "0000001110110000",
15461 => "0000001110110000",
15462 => "0000001110110000",
15463 => "0000001110110000",
15464 => "0000001110110001",
15465 => "0000001110110001",
15466 => "0000001110110001",
15467 => "0000001110110001",
15468 => "0000001110110001",
15469 => "0000001110110010",
15470 => "0000001110110010",
15471 => "0000001110110010",
15472 => "0000001110110010",
15473 => "0000001110110011",
15474 => "0000001110110011",
15475 => "0000001110110011",
15476 => "0000001110110011",
15477 => "0000001110110100",
15478 => "0000001110110100",
15479 => "0000001110110100",
15480 => "0000001110110100",
15481 => "0000001110110100",
15482 => "0000001110110101",
15483 => "0000001110110101",
15484 => "0000001110110101",
15485 => "0000001110110101",
15486 => "0000001110110110",
15487 => "0000001110110110",
15488 => "0000001110110110",
15489 => "0000001110110110",
15490 => "0000001110110111",
15491 => "0000001110110111",
15492 => "0000001110110111",
15493 => "0000001110110111",
15494 => "0000001110110111",
15495 => "0000001110111000",
15496 => "0000001110111000",
15497 => "0000001110111000",
15498 => "0000001110111000",
15499 => "0000001110111001",
15500 => "0000001110111001",
15501 => "0000001110111001",
15502 => "0000001110111001",
15503 => "0000001110111001",
15504 => "0000001110111010",
15505 => "0000001110111010",
15506 => "0000001110111010",
15507 => "0000001110111010",
15508 => "0000001110111011",
15509 => "0000001110111011",
15510 => "0000001110111011",
15511 => "0000001110111011",
15512 => "0000001110111100",
15513 => "0000001110111100",
15514 => "0000001110111100",
15515 => "0000001110111100",
15516 => "0000001110111100",
15517 => "0000001110111101",
15518 => "0000001110111101",
15519 => "0000001110111101",
15520 => "0000001110111101",
15521 => "0000001110111110",
15522 => "0000001110111110",
15523 => "0000001110111110",
15524 => "0000001110111110",
15525 => "0000001110111111",
15526 => "0000001110111111",
15527 => "0000001110111111",
15528 => "0000001110111111",
15529 => "0000001110111111",
15530 => "0000001111000000",
15531 => "0000001111000000",
15532 => "0000001111000000",
15533 => "0000001111000000",
15534 => "0000001111000001",
15535 => "0000001111000001",
15536 => "0000001111000001",
15537 => "0000001111000001",
15538 => "0000001111000010",
15539 => "0000001111000010",
15540 => "0000001111000010",
15541 => "0000001111000010",
15542 => "0000001111000010",
15543 => "0000001111000011",
15544 => "0000001111000011",
15545 => "0000001111000011",
15546 => "0000001111000011",
15547 => "0000001111000100",
15548 => "0000001111000100",
15549 => "0000001111000100",
15550 => "0000001111000100",
15551 => "0000001111000101",
15552 => "0000001111000101",
15553 => "0000001111000101",
15554 => "0000001111000101",
15555 => "0000001111000110",
15556 => "0000001111000110",
15557 => "0000001111000110",
15558 => "0000001111000110",
15559 => "0000001111000110",
15560 => "0000001111000111",
15561 => "0000001111000111",
15562 => "0000001111000111",
15563 => "0000001111000111",
15564 => "0000001111001000",
15565 => "0000001111001000",
15566 => "0000001111001000",
15567 => "0000001111001000",
15568 => "0000001111001001",
15569 => "0000001111001001",
15570 => "0000001111001001",
15571 => "0000001111001001",
15572 => "0000001111001001",
15573 => "0000001111001010",
15574 => "0000001111001010",
15575 => "0000001111001010",
15576 => "0000001111001010",
15577 => "0000001111001011",
15578 => "0000001111001011",
15579 => "0000001111001011",
15580 => "0000001111001011",
15581 => "0000001111001100",
15582 => "0000001111001100",
15583 => "0000001111001100",
15584 => "0000001111001100",
15585 => "0000001111001101",
15586 => "0000001111001101",
15587 => "0000001111001101",
15588 => "0000001111001101",
15589 => "0000001111001101",
15590 => "0000001111001110",
15591 => "0000001111001110",
15592 => "0000001111001110",
15593 => "0000001111001110",
15594 => "0000001111001111",
15595 => "0000001111001111",
15596 => "0000001111001111",
15597 => "0000001111001111",
15598 => "0000001111010000",
15599 => "0000001111010000",
15600 => "0000001111010000",
15601 => "0000001111010000",
15602 => "0000001111010000",
15603 => "0000001111010001",
15604 => "0000001111010001",
15605 => "0000001111010001",
15606 => "0000001111010001",
15607 => "0000001111010010",
15608 => "0000001111010010",
15609 => "0000001111010010",
15610 => "0000001111010010",
15611 => "0000001111010011",
15612 => "0000001111010011",
15613 => "0000001111010011",
15614 => "0000001111010011",
15615 => "0000001111010100",
15616 => "0000001111010100",
15617 => "0000001111010100",
15618 => "0000001111010100",
15619 => "0000001111010100",
15620 => "0000001111010101",
15621 => "0000001111010101",
15622 => "0000001111010101",
15623 => "0000001111010101",
15624 => "0000001111010110",
15625 => "0000001111010110",
15626 => "0000001111010110",
15627 => "0000001111010110",
15628 => "0000001111010111",
15629 => "0000001111010111",
15630 => "0000001111010111",
15631 => "0000001111010111",
15632 => "0000001111011000",
15633 => "0000001111011000",
15634 => "0000001111011000",
15635 => "0000001111011000",
15636 => "0000001111011001",
15637 => "0000001111011001",
15638 => "0000001111011001",
15639 => "0000001111011001",
15640 => "0000001111011001",
15641 => "0000001111011010",
15642 => "0000001111011010",
15643 => "0000001111011010",
15644 => "0000001111011010",
15645 => "0000001111011011",
15646 => "0000001111011011",
15647 => "0000001111011011",
15648 => "0000001111011011",
15649 => "0000001111011100",
15650 => "0000001111011100",
15651 => "0000001111011100",
15652 => "0000001111011100",
15653 => "0000001111011101",
15654 => "0000001111011101",
15655 => "0000001111011101",
15656 => "0000001111011101",
15657 => "0000001111011101",
15658 => "0000001111011110",
15659 => "0000001111011110",
15660 => "0000001111011110",
15661 => "0000001111011110",
15662 => "0000001111011111",
15663 => "0000001111011111",
15664 => "0000001111011111",
15665 => "0000001111011111",
15666 => "0000001111100000",
15667 => "0000001111100000",
15668 => "0000001111100000",
15669 => "0000001111100000",
15670 => "0000001111100001",
15671 => "0000001111100001",
15672 => "0000001111100001",
15673 => "0000001111100001",
15674 => "0000001111100010",
15675 => "0000001111100010",
15676 => "0000001111100010",
15677 => "0000001111100010",
15678 => "0000001111100011",
15679 => "0000001111100011",
15680 => "0000001111100011",
15681 => "0000001111100011",
15682 => "0000001111100011",
15683 => "0000001111100100",
15684 => "0000001111100100",
15685 => "0000001111100100",
15686 => "0000001111100100",
15687 => "0000001111100101",
15688 => "0000001111100101",
15689 => "0000001111100101",
15690 => "0000001111100101",
15691 => "0000001111100110",
15692 => "0000001111100110",
15693 => "0000001111100110",
15694 => "0000001111100110",
15695 => "0000001111100111",
15696 => "0000001111100111",
15697 => "0000001111100111",
15698 => "0000001111100111",
15699 => "0000001111101000",
15700 => "0000001111101000",
15701 => "0000001111101000",
15702 => "0000001111101000",
15703 => "0000001111101001",
15704 => "0000001111101001",
15705 => "0000001111101001",
15706 => "0000001111101001",
15707 => "0000001111101001",
15708 => "0000001111101010",
15709 => "0000001111101010",
15710 => "0000001111101010",
15711 => "0000001111101010",
15712 => "0000001111101011",
15713 => "0000001111101011",
15714 => "0000001111101011",
15715 => "0000001111101011",
15716 => "0000001111101100",
15717 => "0000001111101100",
15718 => "0000001111101100",
15719 => "0000001111101100",
15720 => "0000001111101101",
15721 => "0000001111101101",
15722 => "0000001111101101",
15723 => "0000001111101101",
15724 => "0000001111101110",
15725 => "0000001111101110",
15726 => "0000001111101110",
15727 => "0000001111101110",
15728 => "0000001111101111",
15729 => "0000001111101111",
15730 => "0000001111101111",
15731 => "0000001111101111",
15732 => "0000001111110000",
15733 => "0000001111110000",
15734 => "0000001111110000",
15735 => "0000001111110000",
15736 => "0000001111110000",
15737 => "0000001111110001",
15738 => "0000001111110001",
15739 => "0000001111110001",
15740 => "0000001111110001",
15741 => "0000001111110010",
15742 => "0000001111110010",
15743 => "0000001111110010",
15744 => "0000001111110010",
15745 => "0000001111110011",
15746 => "0000001111110011",
15747 => "0000001111110011",
15748 => "0000001111110011",
15749 => "0000001111110100",
15750 => "0000001111110100",
15751 => "0000001111110100",
15752 => "0000001111110100",
15753 => "0000001111110101",
15754 => "0000001111110101",
15755 => "0000001111110101",
15756 => "0000001111110101",
15757 => "0000001111110110",
15758 => "0000001111110110",
15759 => "0000001111110110",
15760 => "0000001111110110",
15761 => "0000001111110111",
15762 => "0000001111110111",
15763 => "0000001111110111",
15764 => "0000001111110111",
15765 => "0000001111111000",
15766 => "0000001111111000",
15767 => "0000001111111000",
15768 => "0000001111111000",
15769 => "0000001111111001",
15770 => "0000001111111001",
15771 => "0000001111111001",
15772 => "0000001111111001",
15773 => "0000001111111001",
15774 => "0000001111111010",
15775 => "0000001111111010",
15776 => "0000001111111010",
15777 => "0000001111111010",
15778 => "0000001111111011",
15779 => "0000001111111011",
15780 => "0000001111111011",
15781 => "0000001111111011",
15782 => "0000001111111100",
15783 => "0000001111111100",
15784 => "0000001111111100",
15785 => "0000001111111100",
15786 => "0000001111111101",
15787 => "0000001111111101",
15788 => "0000001111111101",
15789 => "0000001111111101",
15790 => "0000001111111110",
15791 => "0000001111111110",
15792 => "0000001111111110",
15793 => "0000001111111110",
15794 => "0000001111111111",
15795 => "0000001111111111",
15796 => "0000001111111111",
15797 => "0000001111111111",
15798 => "0000010000000000",
15799 => "0000010000000000",
15800 => "0000010000000000",
15801 => "0000010000000000",
15802 => "0000010000000001",
15803 => "0000010000000001",
15804 => "0000010000000001",
15805 => "0000010000000001",
15806 => "0000010000000010",
15807 => "0000010000000010",
15808 => "0000010000000010",
15809 => "0000010000000010",
15810 => "0000010000000011",
15811 => "0000010000000011",
15812 => "0000010000000011",
15813 => "0000010000000011",
15814 => "0000010000000100",
15815 => "0000010000000100",
15816 => "0000010000000100",
15817 => "0000010000000100",
15818 => "0000010000000101",
15819 => "0000010000000101",
15820 => "0000010000000101",
15821 => "0000010000000101",
15822 => "0000010000000110",
15823 => "0000010000000110",
15824 => "0000010000000110",
15825 => "0000010000000110",
15826 => "0000010000000111",
15827 => "0000010000000111",
15828 => "0000010000000111",
15829 => "0000010000000111",
15830 => "0000010000001000",
15831 => "0000010000001000",
15832 => "0000010000001000",
15833 => "0000010000001000",
15834 => "0000010000001001",
15835 => "0000010000001001",
15836 => "0000010000001001",
15837 => "0000010000001001",
15838 => "0000010000001010",
15839 => "0000010000001010",
15840 => "0000010000001010",
15841 => "0000010000001010",
15842 => "0000010000001011",
15843 => "0000010000001011",
15844 => "0000010000001011",
15845 => "0000010000001011",
15846 => "0000010000001100",
15847 => "0000010000001100",
15848 => "0000010000001100",
15849 => "0000010000001100",
15850 => "0000010000001101",
15851 => "0000010000001101",
15852 => "0000010000001101",
15853 => "0000010000001101",
15854 => "0000010000001110",
15855 => "0000010000001110",
15856 => "0000010000001110",
15857 => "0000010000001110",
15858 => "0000010000001111",
15859 => "0000010000001111",
15860 => "0000010000001111",
15861 => "0000010000001111",
15862 => "0000010000010000",
15863 => "0000010000010000",
15864 => "0000010000010000",
15865 => "0000010000010000",
15866 => "0000010000010001",
15867 => "0000010000010001",
15868 => "0000010000010001",
15869 => "0000010000010001",
15870 => "0000010000010010",
15871 => "0000010000010010",
15872 => "0000010000010010",
15873 => "0000010000010010",
15874 => "0000010000010011",
15875 => "0000010000010011",
15876 => "0000010000010011",
15877 => "0000010000010011",
15878 => "0000010000010100",
15879 => "0000010000010100",
15880 => "0000010000010100",
15881 => "0000010000010100",
15882 => "0000010000010101",
15883 => "0000010000010101",
15884 => "0000010000010101",
15885 => "0000010000010101",
15886 => "0000010000010110",
15887 => "0000010000010110",
15888 => "0000010000010110",
15889 => "0000010000010110",
15890 => "0000010000010111",
15891 => "0000010000010111",
15892 => "0000010000010111",
15893 => "0000010000010111",
15894 => "0000010000011000",
15895 => "0000010000011000",
15896 => "0000010000011000",
15897 => "0000010000011000",
15898 => "0000010000011001",
15899 => "0000010000011001",
15900 => "0000010000011001",
15901 => "0000010000011001",
15902 => "0000010000011010",
15903 => "0000010000011010",
15904 => "0000010000011010",
15905 => "0000010000011010",
15906 => "0000010000011011",
15907 => "0000010000011011",
15908 => "0000010000011011",
15909 => "0000010000011011",
15910 => "0000010000011100",
15911 => "0000010000011100",
15912 => "0000010000011100",
15913 => "0000010000011100",
15914 => "0000010000011101",
15915 => "0000010000011101",
15916 => "0000010000011101",
15917 => "0000010000011101",
15918 => "0000010000011110",
15919 => "0000010000011110",
15920 => "0000010000011110",
15921 => "0000010000011110",
15922 => "0000010000011111",
15923 => "0000010000011111",
15924 => "0000010000011111",
15925 => "0000010000011111",
15926 => "0000010000100000",
15927 => "0000010000100000",
15928 => "0000010000100000",
15929 => "0000010000100000",
15930 => "0000010000100001",
15931 => "0000010000100001",
15932 => "0000010000100001",
15933 => "0000010000100001",
15934 => "0000010000100010",
15935 => "0000010000100010",
15936 => "0000010000100010",
15937 => "0000010000100010",
15938 => "0000010000100011",
15939 => "0000010000100011",
15940 => "0000010000100011",
15941 => "0000010000100011",
15942 => "0000010000100100",
15943 => "0000010000100100",
15944 => "0000010000100100",
15945 => "0000010000100100",
15946 => "0000010000100101",
15947 => "0000010000100101",
15948 => "0000010000100101",
15949 => "0000010000100101",
15950 => "0000010000100110",
15951 => "0000010000100110",
15952 => "0000010000100110",
15953 => "0000010000100110",
15954 => "0000010000100111",
15955 => "0000010000100111",
15956 => "0000010000100111",
15957 => "0000010000101000",
15958 => "0000010000101000",
15959 => "0000010000101000",
15960 => "0000010000101000",
15961 => "0000010000101001",
15962 => "0000010000101001",
15963 => "0000010000101001",
15964 => "0000010000101001",
15965 => "0000010000101010",
15966 => "0000010000101010",
15967 => "0000010000101010",
15968 => "0000010000101010",
15969 => "0000010000101011",
15970 => "0000010000101011",
15971 => "0000010000101011",
15972 => "0000010000101011",
15973 => "0000010000101100",
15974 => "0000010000101100",
15975 => "0000010000101100",
15976 => "0000010000101100",
15977 => "0000010000101101",
15978 => "0000010000101101",
15979 => "0000010000101101",
15980 => "0000010000101101",
15981 => "0000010000101110",
15982 => "0000010000101110",
15983 => "0000010000101110",
15984 => "0000010000101110",
15985 => "0000010000101111",
15986 => "0000010000101111",
15987 => "0000010000101111",
15988 => "0000010000101111",
15989 => "0000010000110000",
15990 => "0000010000110000",
15991 => "0000010000110000",
15992 => "0000010000110000",
15993 => "0000010000110001",
15994 => "0000010000110001",
15995 => "0000010000110001",
15996 => "0000010000110010",
15997 => "0000010000110010",
15998 => "0000010000110010",
15999 => "0000010000110010",
16000 => "0000010000110011",
16001 => "0000010000110011",
16002 => "0000010000110011",
16003 => "0000010000110011",
16004 => "0000010000110100",
16005 => "0000010000110100",
16006 => "0000010000110100",
16007 => "0000010000110100",
16008 => "0000010000110101",
16009 => "0000010000110101",
16010 => "0000010000110101",
16011 => "0000010000110101",
16012 => "0000010000110110",
16013 => "0000010000110110",
16014 => "0000010000110110",
16015 => "0000010000110110",
16016 => "0000010000110111",
16017 => "0000010000110111",
16018 => "0000010000110111",
16019 => "0000010000110111",
16020 => "0000010000111000",
16021 => "0000010000111000",
16022 => "0000010000111000",
16023 => "0000010000111001",
16024 => "0000010000111001",
16025 => "0000010000111001",
16026 => "0000010000111001",
16027 => "0000010000111010",
16028 => "0000010000111010",
16029 => "0000010000111010",
16030 => "0000010000111010",
16031 => "0000010000111011",
16032 => "0000010000111011",
16033 => "0000010000111011",
16034 => "0000010000111011",
16035 => "0000010000111100",
16036 => "0000010000111100",
16037 => "0000010000111100",
16038 => "0000010000111100",
16039 => "0000010000111101",
16040 => "0000010000111101",
16041 => "0000010000111101",
16042 => "0000010000111101",
16043 => "0000010000111110",
16044 => "0000010000111110",
16045 => "0000010000111110",
16046 => "0000010000111110",
16047 => "0000010000111111",
16048 => "0000010000111111",
16049 => "0000010000111111",
16050 => "0000010001000000",
16051 => "0000010001000000",
16052 => "0000010001000000",
16053 => "0000010001000000",
16054 => "0000010001000001",
16055 => "0000010001000001",
16056 => "0000010001000001",
16057 => "0000010001000001",
16058 => "0000010001000010",
16059 => "0000010001000010",
16060 => "0000010001000010",
16061 => "0000010001000010",
16062 => "0000010001000011",
16063 => "0000010001000011",
16064 => "0000010001000011",
16065 => "0000010001000011",
16066 => "0000010001000100",
16067 => "0000010001000100",
16068 => "0000010001000100",
16069 => "0000010001000101",
16070 => "0000010001000101",
16071 => "0000010001000101",
16072 => "0000010001000101",
16073 => "0000010001000110",
16074 => "0000010001000110",
16075 => "0000010001000110",
16076 => "0000010001000110",
16077 => "0000010001000111",
16078 => "0000010001000111",
16079 => "0000010001000111",
16080 => "0000010001000111",
16081 => "0000010001001000",
16082 => "0000010001001000",
16083 => "0000010001001000",
16084 => "0000010001001000",
16085 => "0000010001001001",
16086 => "0000010001001001",
16087 => "0000010001001001",
16088 => "0000010001001010",
16089 => "0000010001001010",
16090 => "0000010001001010",
16091 => "0000010001001010",
16092 => "0000010001001011",
16093 => "0000010001001011",
16094 => "0000010001001011",
16095 => "0000010001001011",
16096 => "0000010001001100",
16097 => "0000010001001100",
16098 => "0000010001001100",
16099 => "0000010001001100",
16100 => "0000010001001101",
16101 => "0000010001001101",
16102 => "0000010001001101",
16103 => "0000010001001101",
16104 => "0000010001001110",
16105 => "0000010001001110",
16106 => "0000010001001110",
16107 => "0000010001001111",
16108 => "0000010001001111",
16109 => "0000010001001111",
16110 => "0000010001001111",
16111 => "0000010001010000",
16112 => "0000010001010000",
16113 => "0000010001010000",
16114 => "0000010001010000",
16115 => "0000010001010001",
16116 => "0000010001010001",
16117 => "0000010001010001",
16118 => "0000010001010001",
16119 => "0000010001010010",
16120 => "0000010001010010",
16121 => "0000010001010010",
16122 => "0000010001010011",
16123 => "0000010001010011",
16124 => "0000010001010011",
16125 => "0000010001010011",
16126 => "0000010001010100",
16127 => "0000010001010100",
16128 => "0000010001010100",
16129 => "0000010001010100",
16130 => "0000010001010101",
16131 => "0000010001010101",
16132 => "0000010001010101",
16133 => "0000010001010101",
16134 => "0000010001010110",
16135 => "0000010001010110",
16136 => "0000010001010110",
16137 => "0000010001010110",
16138 => "0000010001010111",
16139 => "0000010001010111",
16140 => "0000010001010111",
16141 => "0000010001011000",
16142 => "0000010001011000",
16143 => "0000010001011000",
16144 => "0000010001011000",
16145 => "0000010001011001",
16146 => "0000010001011001",
16147 => "0000010001011001",
16148 => "0000010001011001",
16149 => "0000010001011010",
16150 => "0000010001011010",
16151 => "0000010001011010",
16152 => "0000010001011011",
16153 => "0000010001011011",
16154 => "0000010001011011",
16155 => "0000010001011011",
16156 => "0000010001011100",
16157 => "0000010001011100",
16158 => "0000010001011100",
16159 => "0000010001011100",
16160 => "0000010001011101",
16161 => "0000010001011101",
16162 => "0000010001011101",
16163 => "0000010001011101",
16164 => "0000010001011110",
16165 => "0000010001011110",
16166 => "0000010001011110",
16167 => "0000010001011111",
16168 => "0000010001011111",
16169 => "0000010001011111",
16170 => "0000010001011111",
16171 => "0000010001100000",
16172 => "0000010001100000",
16173 => "0000010001100000",
16174 => "0000010001100000",
16175 => "0000010001100001",
16176 => "0000010001100001",
16177 => "0000010001100001",
16178 => "0000010001100001",
16179 => "0000010001100010",
16180 => "0000010001100010",
16181 => "0000010001100010",
16182 => "0000010001100011",
16183 => "0000010001100011",
16184 => "0000010001100011",
16185 => "0000010001100011",
16186 => "0000010001100100",
16187 => "0000010001100100",
16188 => "0000010001100100",
16189 => "0000010001100100",
16190 => "0000010001100101",
16191 => "0000010001100101",
16192 => "0000010001100101",
16193 => "0000010001100110",
16194 => "0000010001100110",
16195 => "0000010001100110",
16196 => "0000010001100110",
16197 => "0000010001100111",
16198 => "0000010001100111",
16199 => "0000010001100111",
16200 => "0000010001100111",
16201 => "0000010001101000",
16202 => "0000010001101000",
16203 => "0000010001101000",
16204 => "0000010001101001",
16205 => "0000010001101001",
16206 => "0000010001101001",
16207 => "0000010001101001",
16208 => "0000010001101010",
16209 => "0000010001101010",
16210 => "0000010001101010",
16211 => "0000010001101010",
16212 => "0000010001101011",
16213 => "0000010001101011",
16214 => "0000010001101011",
16215 => "0000010001101011",
16216 => "0000010001101100",
16217 => "0000010001101100",
16218 => "0000010001101100",
16219 => "0000010001101101",
16220 => "0000010001101101",
16221 => "0000010001101101",
16222 => "0000010001101101",
16223 => "0000010001101110",
16224 => "0000010001101110",
16225 => "0000010001101110",
16226 => "0000010001101110",
16227 => "0000010001101111",
16228 => "0000010001101111",
16229 => "0000010001101111",
16230 => "0000010001110000",
16231 => "0000010001110000",
16232 => "0000010001110000",
16233 => "0000010001110000",
16234 => "0000010001110001",
16235 => "0000010001110001",
16236 => "0000010001110001",
16237 => "0000010001110001",
16238 => "0000010001110010",
16239 => "0000010001110010",
16240 => "0000010001110010",
16241 => "0000010001110011",
16242 => "0000010001110011",
16243 => "0000010001110011",
16244 => "0000010001110011",
16245 => "0000010001110100",
16246 => "0000010001110100",
16247 => "0000010001110100",
16248 => "0000010001110100",
16249 => "0000010001110101",
16250 => "0000010001110101",
16251 => "0000010001110101",
16252 => "0000010001110110",
16253 => "0000010001110110",
16254 => "0000010001110110",
16255 => "0000010001110110",
16256 => "0000010001110111",
16257 => "0000010001110111",
16258 => "0000010001110111",
16259 => "0000010001111000",
16260 => "0000010001111000",
16261 => "0000010001111000",
16262 => "0000010001111000",
16263 => "0000010001111001",
16264 => "0000010001111001",
16265 => "0000010001111001",
16266 => "0000010001111001",
16267 => "0000010001111010",
16268 => "0000010001111010",
16269 => "0000010001111010",
16270 => "0000010001111011",
16271 => "0000010001111011",
16272 => "0000010001111011",
16273 => "0000010001111011",
16274 => "0000010001111100",
16275 => "0000010001111100",
16276 => "0000010001111100",
16277 => "0000010001111100",
16278 => "0000010001111101",
16279 => "0000010001111101",
16280 => "0000010001111101",
16281 => "0000010001111110",
16282 => "0000010001111110",
16283 => "0000010001111110",
16284 => "0000010001111110",
16285 => "0000010001111111",
16286 => "0000010001111111",
16287 => "0000010001111111",
16288 => "0000010001111111",
16289 => "0000010010000000",
16290 => "0000010010000000",
16291 => "0000010010000000",
16292 => "0000010010000001",
16293 => "0000010010000001",
16294 => "0000010010000001",
16295 => "0000010010000001",
16296 => "0000010010000010",
16297 => "0000010010000010",
16298 => "0000010010000010",
16299 => "0000010010000011",
16300 => "0000010010000011",
16301 => "0000010010000011",
16302 => "0000010010000011",
16303 => "0000010010000100",
16304 => "0000010010000100",
16305 => "0000010010000100",
16306 => "0000010010000100",
16307 => "0000010010000101",
16308 => "0000010010000101",
16309 => "0000010010000101",
16310 => "0000010010000110",
16311 => "0000010010000110",
16312 => "0000010010000110",
16313 => "0000010010000110",
16314 => "0000010010000111",
16315 => "0000010010000111",
16316 => "0000010010000111",
16317 => "0000010010001000",
16318 => "0000010010001000",
16319 => "0000010010001000",
16320 => "0000010010001000",
16321 => "0000010010001001",
16322 => "0000010010001001",
16323 => "0000010010001001",
16324 => "0000010010001001",
16325 => "0000010010001010",
16326 => "0000010010001010",
16327 => "0000010010001010",
16328 => "0000010010001011",
16329 => "0000010010001011",
16330 => "0000010010001011",
16331 => "0000010010001011",
16332 => "0000010010001100",
16333 => "0000010010001100",
16334 => "0000010010001100",
16335 => "0000010010001101",
16336 => "0000010010001101",
16337 => "0000010010001101",
16338 => "0000010010001101",
16339 => "0000010010001110",
16340 => "0000010010001110",
16341 => "0000010010001110",
16342 => "0000010010001111",
16343 => "0000010010001111",
16344 => "0000010010001111",
16345 => "0000010010001111",
16346 => "0000010010010000",
16347 => "0000010010010000",
16348 => "0000010010010000",
16349 => "0000010010010000",
16350 => "0000010010010001",
16351 => "0000010010010001",
16352 => "0000010010010001",
16353 => "0000010010010010",
16354 => "0000010010010010",
16355 => "0000010010010010",
16356 => "0000010010010010",
16357 => "0000010010010011",
16358 => "0000010010010011",
16359 => "0000010010010011",
16360 => "0000010010010100",
16361 => "0000010010010100",
16362 => "0000010010010100",
16363 => "0000010010010100",
16364 => "0000010010010101",
16365 => "0000010010010101",
16366 => "0000010010010101",
16367 => "0000010010010110",
16368 => "0000010010010110",
16369 => "0000010010010110",
16370 => "0000010010010110",
16371 => "0000010010010111",
16372 => "0000010010010111",
16373 => "0000010010010111",
16374 => "0000010010010111",
16375 => "0000010010011000",
16376 => "0000010010011000",
16377 => "0000010010011000",
16378 => "0000010010011001",
16379 => "0000010010011001",
16380 => "0000010010011001",
16381 => "0000010010011001",
16382 => "0000010010011010",
16383 => "0000010010011010",
16384 => "0000010010011010",
16385 => "0000010010011011",
16386 => "0000010010011011",
16387 => "0000010010011011",
16388 => "0000010010011011",
16389 => "0000010010011100",
16390 => "0000010010011100",
16391 => "0000010010011100",
16392 => "0000010010011101",
16393 => "0000010010011101",
16394 => "0000010010011101",
16395 => "0000010010011101",
16396 => "0000010010011110",
16397 => "0000010010011110",
16398 => "0000010010011110",
16399 => "0000010010011111",
16400 => "0000010010011111",
16401 => "0000010010011111",
16402 => "0000010010011111",
16403 => "0000010010100000",
16404 => "0000010010100000",
16405 => "0000010010100000",
16406 => "0000010010100001",
16407 => "0000010010100001",
16408 => "0000010010100001",
16409 => "0000010010100001",
16410 => "0000010010100010",
16411 => "0000010010100010",
16412 => "0000010010100010",
16413 => "0000010010100011",
16414 => "0000010010100011",
16415 => "0000010010100011",
16416 => "0000010010100011",
16417 => "0000010010100100",
16418 => "0000010010100100",
16419 => "0000010010100100",
16420 => "0000010010100101",
16421 => "0000010010100101",
16422 => "0000010010100101",
16423 => "0000010010100101",
16424 => "0000010010100110",
16425 => "0000010010100110",
16426 => "0000010010100110",
16427 => "0000010010100111",
16428 => "0000010010100111",
16429 => "0000010010100111",
16430 => "0000010010100111",
16431 => "0000010010101000",
16432 => "0000010010101000",
16433 => "0000010010101000",
16434 => "0000010010101001",
16435 => "0000010010101001",
16436 => "0000010010101001",
16437 => "0000010010101001",
16438 => "0000010010101010",
16439 => "0000010010101010",
16440 => "0000010010101010",
16441 => "0000010010101011",
16442 => "0000010010101011",
16443 => "0000010010101011",
16444 => "0000010010101011",
16445 => "0000010010101100",
16446 => "0000010010101100",
16447 => "0000010010101100",
16448 => "0000010010101101",
16449 => "0000010010101101",
16450 => "0000010010101101",
16451 => "0000010010101101",
16452 => "0000010010101110",
16453 => "0000010010101110",
16454 => "0000010010101110",
16455 => "0000010010101111",
16456 => "0000010010101111",
16457 => "0000010010101111",
16458 => "0000010010101111",
16459 => "0000010010110000",
16460 => "0000010010110000",
16461 => "0000010010110000",
16462 => "0000010010110001",
16463 => "0000010010110001",
16464 => "0000010010110001",
16465 => "0000010010110001",
16466 => "0000010010110010",
16467 => "0000010010110010",
16468 => "0000010010110010",
16469 => "0000010010110011",
16470 => "0000010010110011",
16471 => "0000010010110011",
16472 => "0000010010110011",
16473 => "0000010010110100",
16474 => "0000010010110100",
16475 => "0000010010110100",
16476 => "0000010010110101",
16477 => "0000010010110101",
16478 => "0000010010110101",
16479 => "0000010010110101",
16480 => "0000010010110110",
16481 => "0000010010110110",
16482 => "0000010010110110",
16483 => "0000010010110111",
16484 => "0000010010110111",
16485 => "0000010010110111",
16486 => "0000010010110111",
16487 => "0000010010111000",
16488 => "0000010010111000",
16489 => "0000010010111000",
16490 => "0000010010111001",
16491 => "0000010010111001",
16492 => "0000010010111001",
16493 => "0000010010111010",
16494 => "0000010010111010",
16495 => "0000010010111010",
16496 => "0000010010111010",
16497 => "0000010010111011",
16498 => "0000010010111011",
16499 => "0000010010111011",
16500 => "0000010010111100",
16501 => "0000010010111100",
16502 => "0000010010111100",
16503 => "0000010010111100",
16504 => "0000010010111101",
16505 => "0000010010111101",
16506 => "0000010010111101",
16507 => "0000010010111110",
16508 => "0000010010111110",
16509 => "0000010010111110",
16510 => "0000010010111110",
16511 => "0000010010111111",
16512 => "0000010010111111",
16513 => "0000010010111111",
16514 => "0000010011000000",
16515 => "0000010011000000",
16516 => "0000010011000000",
16517 => "0000010011000000",
16518 => "0000010011000001",
16519 => "0000010011000001",
16520 => "0000010011000001",
16521 => "0000010011000010",
16522 => "0000010011000010",
16523 => "0000010011000010",
16524 => "0000010011000011",
16525 => "0000010011000011",
16526 => "0000010011000011",
16527 => "0000010011000011",
16528 => "0000010011000100",
16529 => "0000010011000100",
16530 => "0000010011000100",
16531 => "0000010011000101",
16532 => "0000010011000101",
16533 => "0000010011000101",
16534 => "0000010011000101",
16535 => "0000010011000110",
16536 => "0000010011000110",
16537 => "0000010011000110",
16538 => "0000010011000111",
16539 => "0000010011000111",
16540 => "0000010011000111",
16541 => "0000010011001000",
16542 => "0000010011001000",
16543 => "0000010011001000",
16544 => "0000010011001000",
16545 => "0000010011001001",
16546 => "0000010011001001",
16547 => "0000010011001001",
16548 => "0000010011001010",
16549 => "0000010011001010",
16550 => "0000010011001010",
16551 => "0000010011001010",
16552 => "0000010011001011",
16553 => "0000010011001011",
16554 => "0000010011001011",
16555 => "0000010011001100",
16556 => "0000010011001100",
16557 => "0000010011001100",
16558 => "0000010011001101",
16559 => "0000010011001101",
16560 => "0000010011001101",
16561 => "0000010011001101",
16562 => "0000010011001110",
16563 => "0000010011001110",
16564 => "0000010011001110",
16565 => "0000010011001111",
16566 => "0000010011001111",
16567 => "0000010011001111",
16568 => "0000010011001111",
16569 => "0000010011010000",
16570 => "0000010011010000",
16571 => "0000010011010000",
16572 => "0000010011010001",
16573 => "0000010011010001",
16574 => "0000010011010001",
16575 => "0000010011010010",
16576 => "0000010011010010",
16577 => "0000010011010010",
16578 => "0000010011010010",
16579 => "0000010011010011",
16580 => "0000010011010011",
16581 => "0000010011010011",
16582 => "0000010011010100",
16583 => "0000010011010100",
16584 => "0000010011010100",
16585 => "0000010011010100",
16586 => "0000010011010101",
16587 => "0000010011010101",
16588 => "0000010011010101",
16589 => "0000010011010110",
16590 => "0000010011010110",
16591 => "0000010011010110",
16592 => "0000010011010111",
16593 => "0000010011010111",
16594 => "0000010011010111",
16595 => "0000010011010111",
16596 => "0000010011011000",
16597 => "0000010011011000",
16598 => "0000010011011000",
16599 => "0000010011011001",
16600 => "0000010011011001",
16601 => "0000010011011001",
16602 => "0000010011011010",
16603 => "0000010011011010",
16604 => "0000010011011010",
16605 => "0000010011011010",
16606 => "0000010011011011",
16607 => "0000010011011011",
16608 => "0000010011011011",
16609 => "0000010011011100",
16610 => "0000010011011100",
16611 => "0000010011011100",
16612 => "0000010011011101",
16613 => "0000010011011101",
16614 => "0000010011011101",
16615 => "0000010011011101",
16616 => "0000010011011110",
16617 => "0000010011011110",
16618 => "0000010011011110",
16619 => "0000010011011111",
16620 => "0000010011011111",
16621 => "0000010011011111",
16622 => "0000010011011111",
16623 => "0000010011100000",
16624 => "0000010011100000",
16625 => "0000010011100000",
16626 => "0000010011100001",
16627 => "0000010011100001",
16628 => "0000010011100001",
16629 => "0000010011100010",
16630 => "0000010011100010",
16631 => "0000010011100010",
16632 => "0000010011100010",
16633 => "0000010011100011",
16634 => "0000010011100011",
16635 => "0000010011100011",
16636 => "0000010011100100",
16637 => "0000010011100100",
16638 => "0000010011100100",
16639 => "0000010011100101",
16640 => "0000010011100101",
16641 => "0000010011100101",
16642 => "0000010011100101",
16643 => "0000010011100110",
16644 => "0000010011100110",
16645 => "0000010011100110",
16646 => "0000010011100111",
16647 => "0000010011100111",
16648 => "0000010011100111",
16649 => "0000010011101000",
16650 => "0000010011101000",
16651 => "0000010011101000",
16652 => "0000010011101000",
16653 => "0000010011101001",
16654 => "0000010011101001",
16655 => "0000010011101001",
16656 => "0000010011101010",
16657 => "0000010011101010",
16658 => "0000010011101010",
16659 => "0000010011101011",
16660 => "0000010011101011",
16661 => "0000010011101011",
16662 => "0000010011101100",
16663 => "0000010011101100",
16664 => "0000010011101100",
16665 => "0000010011101100",
16666 => "0000010011101101",
16667 => "0000010011101101",
16668 => "0000010011101101",
16669 => "0000010011101110",
16670 => "0000010011101110",
16671 => "0000010011101110",
16672 => "0000010011101111",
16673 => "0000010011101111",
16674 => "0000010011101111",
16675 => "0000010011101111",
16676 => "0000010011110000",
16677 => "0000010011110000",
16678 => "0000010011110000",
16679 => "0000010011110001",
16680 => "0000010011110001",
16681 => "0000010011110001",
16682 => "0000010011110010",
16683 => "0000010011110010",
16684 => "0000010011110010",
16685 => "0000010011110010",
16686 => "0000010011110011",
16687 => "0000010011110011",
16688 => "0000010011110011",
16689 => "0000010011110100",
16690 => "0000010011110100",
16691 => "0000010011110100",
16692 => "0000010011110101",
16693 => "0000010011110101",
16694 => "0000010011110101",
16695 => "0000010011110110",
16696 => "0000010011110110",
16697 => "0000010011110110",
16698 => "0000010011110110",
16699 => "0000010011110111",
16700 => "0000010011110111",
16701 => "0000010011110111",
16702 => "0000010011111000",
16703 => "0000010011111000",
16704 => "0000010011111000",
16705 => "0000010011111001",
16706 => "0000010011111001",
16707 => "0000010011111001",
16708 => "0000010011111001",
16709 => "0000010011111010",
16710 => "0000010011111010",
16711 => "0000010011111010",
16712 => "0000010011111011",
16713 => "0000010011111011",
16714 => "0000010011111011",
16715 => "0000010011111100",
16716 => "0000010011111100",
16717 => "0000010011111100",
16718 => "0000010011111101",
16719 => "0000010011111101",
16720 => "0000010011111101",
16721 => "0000010011111101",
16722 => "0000010011111110",
16723 => "0000010011111110",
16724 => "0000010011111110",
16725 => "0000010011111111",
16726 => "0000010011111111",
16727 => "0000010011111111",
16728 => "0000010100000000",
16729 => "0000010100000000",
16730 => "0000010100000000",
16731 => "0000010100000000",
16732 => "0000010100000001",
16733 => "0000010100000001",
16734 => "0000010100000001",
16735 => "0000010100000010",
16736 => "0000010100000010",
16737 => "0000010100000010",
16738 => "0000010100000011",
16739 => "0000010100000011",
16740 => "0000010100000011",
16741 => "0000010100000100",
16742 => "0000010100000100",
16743 => "0000010100000100",
16744 => "0000010100000100",
16745 => "0000010100000101",
16746 => "0000010100000101",
16747 => "0000010100000101",
16748 => "0000010100000110",
16749 => "0000010100000110",
16750 => "0000010100000110",
16751 => "0000010100000111",
16752 => "0000010100000111",
16753 => "0000010100000111",
16754 => "0000010100001000",
16755 => "0000010100001000",
16756 => "0000010100001000",
16757 => "0000010100001000",
16758 => "0000010100001001",
16759 => "0000010100001001",
16760 => "0000010100001001",
16761 => "0000010100001010",
16762 => "0000010100001010",
16763 => "0000010100001010",
16764 => "0000010100001011",
16765 => "0000010100001011",
16766 => "0000010100001011",
16767 => "0000010100001100",
16768 => "0000010100001100",
16769 => "0000010100001100",
16770 => "0000010100001101",
16771 => "0000010100001101",
16772 => "0000010100001101",
16773 => "0000010100001101",
16774 => "0000010100001110",
16775 => "0000010100001110",
16776 => "0000010100001110",
16777 => "0000010100001111",
16778 => "0000010100001111",
16779 => "0000010100001111",
16780 => "0000010100010000",
16781 => "0000010100010000",
16782 => "0000010100010000",
16783 => "0000010100010001",
16784 => "0000010100010001",
16785 => "0000010100010001",
16786 => "0000010100010001",
16787 => "0000010100010010",
16788 => "0000010100010010",
16789 => "0000010100010010",
16790 => "0000010100010011",
16791 => "0000010100010011",
16792 => "0000010100010011",
16793 => "0000010100010100",
16794 => "0000010100010100",
16795 => "0000010100010100",
16796 => "0000010100010101",
16797 => "0000010100010101",
16798 => "0000010100010101",
16799 => "0000010100010110",
16800 => "0000010100010110",
16801 => "0000010100010110",
16802 => "0000010100010110",
16803 => "0000010100010111",
16804 => "0000010100010111",
16805 => "0000010100010111",
16806 => "0000010100011000",
16807 => "0000010100011000",
16808 => "0000010100011000",
16809 => "0000010100011001",
16810 => "0000010100011001",
16811 => "0000010100011001",
16812 => "0000010100011010",
16813 => "0000010100011010",
16814 => "0000010100011010",
16815 => "0000010100011011",
16816 => "0000010100011011",
16817 => "0000010100011011",
16818 => "0000010100011011",
16819 => "0000010100011100",
16820 => "0000010100011100",
16821 => "0000010100011100",
16822 => "0000010100011101",
16823 => "0000010100011101",
16824 => "0000010100011101",
16825 => "0000010100011110",
16826 => "0000010100011110",
16827 => "0000010100011110",
16828 => "0000010100011111",
16829 => "0000010100011111",
16830 => "0000010100011111",
16831 => "0000010100100000",
16832 => "0000010100100000",
16833 => "0000010100100000",
16834 => "0000010100100000",
16835 => "0000010100100001",
16836 => "0000010100100001",
16837 => "0000010100100001",
16838 => "0000010100100010",
16839 => "0000010100100010",
16840 => "0000010100100010",
16841 => "0000010100100011",
16842 => "0000010100100011",
16843 => "0000010100100011",
16844 => "0000010100100100",
16845 => "0000010100100100",
16846 => "0000010100100100",
16847 => "0000010100100101",
16848 => "0000010100100101",
16849 => "0000010100100101",
16850 => "0000010100100110",
16851 => "0000010100100110",
16852 => "0000010100100110",
16853 => "0000010100100110",
16854 => "0000010100100111",
16855 => "0000010100100111",
16856 => "0000010100100111",
16857 => "0000010100101000",
16858 => "0000010100101000",
16859 => "0000010100101000",
16860 => "0000010100101001",
16861 => "0000010100101001",
16862 => "0000010100101001",
16863 => "0000010100101010",
16864 => "0000010100101010",
16865 => "0000010100101010",
16866 => "0000010100101011",
16867 => "0000010100101011",
16868 => "0000010100101011",
16869 => "0000010100101100",
16870 => "0000010100101100",
16871 => "0000010100101100",
16872 => "0000010100101100",
16873 => "0000010100101101",
16874 => "0000010100101101",
16875 => "0000010100101101",
16876 => "0000010100101110",
16877 => "0000010100101110",
16878 => "0000010100101110",
16879 => "0000010100101111",
16880 => "0000010100101111",
16881 => "0000010100101111",
16882 => "0000010100110000",
16883 => "0000010100110000",
16884 => "0000010100110000",
16885 => "0000010100110001",
16886 => "0000010100110001",
16887 => "0000010100110001",
16888 => "0000010100110010",
16889 => "0000010100110010",
16890 => "0000010100110010",
16891 => "0000010100110010",
16892 => "0000010100110011",
16893 => "0000010100110011",
16894 => "0000010100110011",
16895 => "0000010100110100",
16896 => "0000010100110100",
16897 => "0000010100110100",
16898 => "0000010100110101",
16899 => "0000010100110101",
16900 => "0000010100110101",
16901 => "0000010100110110",
16902 => "0000010100110110",
16903 => "0000010100110110",
16904 => "0000010100110111",
16905 => "0000010100110111",
16906 => "0000010100110111",
16907 => "0000010100111000",
16908 => "0000010100111000",
16909 => "0000010100111000",
16910 => "0000010100111001",
16911 => "0000010100111001",
16912 => "0000010100111001",
16913 => "0000010100111010",
16914 => "0000010100111010",
16915 => "0000010100111010",
16916 => "0000010100111010",
16917 => "0000010100111011",
16918 => "0000010100111011",
16919 => "0000010100111011",
16920 => "0000010100111100",
16921 => "0000010100111100",
16922 => "0000010100111100",
16923 => "0000010100111101",
16924 => "0000010100111101",
16925 => "0000010100111101",
16926 => "0000010100111110",
16927 => "0000010100111110",
16928 => "0000010100111110",
16929 => "0000010100111111",
16930 => "0000010100111111",
16931 => "0000010100111111",
16932 => "0000010101000000",
16933 => "0000010101000000",
16934 => "0000010101000000",
16935 => "0000010101000001",
16936 => "0000010101000001",
16937 => "0000010101000001",
16938 => "0000010101000010",
16939 => "0000010101000010",
16940 => "0000010101000010",
16941 => "0000010101000011",
16942 => "0000010101000011",
16943 => "0000010101000011",
16944 => "0000010101000011",
16945 => "0000010101000100",
16946 => "0000010101000100",
16947 => "0000010101000100",
16948 => "0000010101000101",
16949 => "0000010101000101",
16950 => "0000010101000101",
16951 => "0000010101000110",
16952 => "0000010101000110",
16953 => "0000010101000110",
16954 => "0000010101000111",
16955 => "0000010101000111",
16956 => "0000010101000111",
16957 => "0000010101001000",
16958 => "0000010101001000",
16959 => "0000010101001000",
16960 => "0000010101001001",
16961 => "0000010101001001",
16962 => "0000010101001001",
16963 => "0000010101001010",
16964 => "0000010101001010",
16965 => "0000010101001010",
16966 => "0000010101001011",
16967 => "0000010101001011",
16968 => "0000010101001011",
16969 => "0000010101001100",
16970 => "0000010101001100",
16971 => "0000010101001100",
16972 => "0000010101001101",
16973 => "0000010101001101",
16974 => "0000010101001101",
16975 => "0000010101001101",
16976 => "0000010101001110",
16977 => "0000010101001110",
16978 => "0000010101001110",
16979 => "0000010101001111",
16980 => "0000010101001111",
16981 => "0000010101001111",
16982 => "0000010101010000",
16983 => "0000010101010000",
16984 => "0000010101010000",
16985 => "0000010101010001",
16986 => "0000010101010001",
16987 => "0000010101010001",
16988 => "0000010101010010",
16989 => "0000010101010010",
16990 => "0000010101010010",
16991 => "0000010101010011",
16992 => "0000010101010011",
16993 => "0000010101010011",
16994 => "0000010101010100",
16995 => "0000010101010100",
16996 => "0000010101010100",
16997 => "0000010101010101",
16998 => "0000010101010101",
16999 => "0000010101010101",
17000 => "0000010101010110",
17001 => "0000010101010110",
17002 => "0000010101010110",
17003 => "0000010101010111",
17004 => "0000010101010111",
17005 => "0000010101010111",
17006 => "0000010101011000",
17007 => "0000010101011000",
17008 => "0000010101011000",
17009 => "0000010101011001",
17010 => "0000010101011001",
17011 => "0000010101011001",
17012 => "0000010101011010",
17013 => "0000010101011010",
17014 => "0000010101011010",
17015 => "0000010101011011",
17016 => "0000010101011011",
17017 => "0000010101011011",
17018 => "0000010101011100",
17019 => "0000010101011100",
17020 => "0000010101011100",
17021 => "0000010101011101",
17022 => "0000010101011101",
17023 => "0000010101011101",
17024 => "0000010101011101",
17025 => "0000010101011110",
17026 => "0000010101011110",
17027 => "0000010101011110",
17028 => "0000010101011111",
17029 => "0000010101011111",
17030 => "0000010101011111",
17031 => "0000010101100000",
17032 => "0000010101100000",
17033 => "0000010101100000",
17034 => "0000010101100001",
17035 => "0000010101100001",
17036 => "0000010101100001",
17037 => "0000010101100010",
17038 => "0000010101100010",
17039 => "0000010101100010",
17040 => "0000010101100011",
17041 => "0000010101100011",
17042 => "0000010101100011",
17043 => "0000010101100100",
17044 => "0000010101100100",
17045 => "0000010101100100",
17046 => "0000010101100101",
17047 => "0000010101100101",
17048 => "0000010101100101",
17049 => "0000010101100110",
17050 => "0000010101100110",
17051 => "0000010101100110",
17052 => "0000010101100111",
17053 => "0000010101100111",
17054 => "0000010101100111",
17055 => "0000010101101000",
17056 => "0000010101101000",
17057 => "0000010101101000",
17058 => "0000010101101001",
17059 => "0000010101101001",
17060 => "0000010101101001",
17061 => "0000010101101010",
17062 => "0000010101101010",
17063 => "0000010101101010",
17064 => "0000010101101011",
17065 => "0000010101101011",
17066 => "0000010101101011",
17067 => "0000010101101100",
17068 => "0000010101101100",
17069 => "0000010101101100",
17070 => "0000010101101101",
17071 => "0000010101101101",
17072 => "0000010101101101",
17073 => "0000010101101110",
17074 => "0000010101101110",
17075 => "0000010101101110",
17076 => "0000010101101111",
17077 => "0000010101101111",
17078 => "0000010101101111",
17079 => "0000010101110000",
17080 => "0000010101110000",
17081 => "0000010101110000",
17082 => "0000010101110001",
17083 => "0000010101110001",
17084 => "0000010101110001",
17085 => "0000010101110010",
17086 => "0000010101110010",
17087 => "0000010101110010",
17088 => "0000010101110011",
17089 => "0000010101110011",
17090 => "0000010101110011",
17091 => "0000010101110100",
17092 => "0000010101110100",
17093 => "0000010101110100",
17094 => "0000010101110101",
17095 => "0000010101110101",
17096 => "0000010101110101",
17097 => "0000010101110110",
17098 => "0000010101110110",
17099 => "0000010101110110",
17100 => "0000010101110111",
17101 => "0000010101110111",
17102 => "0000010101110111",
17103 => "0000010101111000",
17104 => "0000010101111000",
17105 => "0000010101111000",
17106 => "0000010101111001",
17107 => "0000010101111001",
17108 => "0000010101111001",
17109 => "0000010101111010",
17110 => "0000010101111010",
17111 => "0000010101111010",
17112 => "0000010101111011",
17113 => "0000010101111011",
17114 => "0000010101111011",
17115 => "0000010101111100",
17116 => "0000010101111100",
17117 => "0000010101111100",
17118 => "0000010101111101",
17119 => "0000010101111101",
17120 => "0000010101111101",
17121 => "0000010101111110",
17122 => "0000010101111110",
17123 => "0000010101111110",
17124 => "0000010101111111",
17125 => "0000010101111111",
17126 => "0000010101111111",
17127 => "0000010110000000",
17128 => "0000010110000000",
17129 => "0000010110000000",
17130 => "0000010110000001",
17131 => "0000010110000001",
17132 => "0000010110000001",
17133 => "0000010110000010",
17134 => "0000010110000010",
17135 => "0000010110000010",
17136 => "0000010110000011",
17137 => "0000010110000011",
17138 => "0000010110000011",
17139 => "0000010110000100",
17140 => "0000010110000100",
17141 => "0000010110000100",
17142 => "0000010110000101",
17143 => "0000010110000101",
17144 => "0000010110000101",
17145 => "0000010110000110",
17146 => "0000010110000110",
17147 => "0000010110000110",
17148 => "0000010110000111",
17149 => "0000010110000111",
17150 => "0000010110000111",
17151 => "0000010110001000",
17152 => "0000010110001000",
17153 => "0000010110001001",
17154 => "0000010110001001",
17155 => "0000010110001001",
17156 => "0000010110001010",
17157 => "0000010110001010",
17158 => "0000010110001010",
17159 => "0000010110001011",
17160 => "0000010110001011",
17161 => "0000010110001011",
17162 => "0000010110001100",
17163 => "0000010110001100",
17164 => "0000010110001100",
17165 => "0000010110001101",
17166 => "0000010110001101",
17167 => "0000010110001101",
17168 => "0000010110001110",
17169 => "0000010110001110",
17170 => "0000010110001110",
17171 => "0000010110001111",
17172 => "0000010110001111",
17173 => "0000010110001111",
17174 => "0000010110010000",
17175 => "0000010110010000",
17176 => "0000010110010000",
17177 => "0000010110010001",
17178 => "0000010110010001",
17179 => "0000010110010001",
17180 => "0000010110010010",
17181 => "0000010110010010",
17182 => "0000010110010010",
17183 => "0000010110010011",
17184 => "0000010110010011",
17185 => "0000010110010011",
17186 => "0000010110010100",
17187 => "0000010110010100",
17188 => "0000010110010100",
17189 => "0000010110010101",
17190 => "0000010110010101",
17191 => "0000010110010101",
17192 => "0000010110010110",
17193 => "0000010110010110",
17194 => "0000010110010110",
17195 => "0000010110010111",
17196 => "0000010110010111",
17197 => "0000010110010111",
17198 => "0000010110011000",
17199 => "0000010110011000",
17200 => "0000010110011001",
17201 => "0000010110011001",
17202 => "0000010110011001",
17203 => "0000010110011010",
17204 => "0000010110011010",
17205 => "0000010110011010",
17206 => "0000010110011011",
17207 => "0000010110011011",
17208 => "0000010110011011",
17209 => "0000010110011100",
17210 => "0000010110011100",
17211 => "0000010110011100",
17212 => "0000010110011101",
17213 => "0000010110011101",
17214 => "0000010110011101",
17215 => "0000010110011110",
17216 => "0000010110011110",
17217 => "0000010110011110",
17218 => "0000010110011111",
17219 => "0000010110011111",
17220 => "0000010110011111",
17221 => "0000010110100000",
17222 => "0000010110100000",
17223 => "0000010110100000",
17224 => "0000010110100001",
17225 => "0000010110100001",
17226 => "0000010110100001",
17227 => "0000010110100010",
17228 => "0000010110100010",
17229 => "0000010110100010",
17230 => "0000010110100011",
17231 => "0000010110100011",
17232 => "0000010110100011",
17233 => "0000010110100100",
17234 => "0000010110100100",
17235 => "0000010110100101",
17236 => "0000010110100101",
17237 => "0000010110100101",
17238 => "0000010110100110",
17239 => "0000010110100110",
17240 => "0000010110100110",
17241 => "0000010110100111",
17242 => "0000010110100111",
17243 => "0000010110100111",
17244 => "0000010110101000",
17245 => "0000010110101000",
17246 => "0000010110101000",
17247 => "0000010110101001",
17248 => "0000010110101001",
17249 => "0000010110101001",
17250 => "0000010110101010",
17251 => "0000010110101010",
17252 => "0000010110101010",
17253 => "0000010110101011",
17254 => "0000010110101011",
17255 => "0000010110101011",
17256 => "0000010110101100",
17257 => "0000010110101100",
17258 => "0000010110101100",
17259 => "0000010110101101",
17260 => "0000010110101101",
17261 => "0000010110101110",
17262 => "0000010110101110",
17263 => "0000010110101110",
17264 => "0000010110101111",
17265 => "0000010110101111",
17266 => "0000010110101111",
17267 => "0000010110110000",
17268 => "0000010110110000",
17269 => "0000010110110000",
17270 => "0000010110110001",
17271 => "0000010110110001",
17272 => "0000010110110001",
17273 => "0000010110110010",
17274 => "0000010110110010",
17275 => "0000010110110010",
17276 => "0000010110110011",
17277 => "0000010110110011",
17278 => "0000010110110011",
17279 => "0000010110110100",
17280 => "0000010110110100",
17281 => "0000010110110100",
17282 => "0000010110110101",
17283 => "0000010110110101",
17284 => "0000010110110110",
17285 => "0000010110110110",
17286 => "0000010110110110",
17287 => "0000010110110111",
17288 => "0000010110110111",
17289 => "0000010110110111",
17290 => "0000010110111000",
17291 => "0000010110111000",
17292 => "0000010110111000",
17293 => "0000010110111001",
17294 => "0000010110111001",
17295 => "0000010110111001",
17296 => "0000010110111010",
17297 => "0000010110111010",
17298 => "0000010110111010",
17299 => "0000010110111011",
17300 => "0000010110111011",
17301 => "0000010110111011",
17302 => "0000010110111100",
17303 => "0000010110111100",
17304 => "0000010110111101",
17305 => "0000010110111101",
17306 => "0000010110111101",
17307 => "0000010110111110",
17308 => "0000010110111110",
17309 => "0000010110111110",
17310 => "0000010110111111",
17311 => "0000010110111111",
17312 => "0000010110111111",
17313 => "0000010111000000",
17314 => "0000010111000000",
17315 => "0000010111000000",
17316 => "0000010111000001",
17317 => "0000010111000001",
17318 => "0000010111000001",
17319 => "0000010111000010",
17320 => "0000010111000010",
17321 => "0000010111000011",
17322 => "0000010111000011",
17323 => "0000010111000011",
17324 => "0000010111000100",
17325 => "0000010111000100",
17326 => "0000010111000100",
17327 => "0000010111000101",
17328 => "0000010111000101",
17329 => "0000010111000101",
17330 => "0000010111000110",
17331 => "0000010111000110",
17332 => "0000010111000110",
17333 => "0000010111000111",
17334 => "0000010111000111",
17335 => "0000010111000111",
17336 => "0000010111001000",
17337 => "0000010111001000",
17338 => "0000010111001000",
17339 => "0000010111001001",
17340 => "0000010111001001",
17341 => "0000010111001010",
17342 => "0000010111001010",
17343 => "0000010111001010",
17344 => "0000010111001011",
17345 => "0000010111001011",
17346 => "0000010111001011",
17347 => "0000010111001100",
17348 => "0000010111001100",
17349 => "0000010111001100",
17350 => "0000010111001101",
17351 => "0000010111001101",
17352 => "0000010111001101",
17353 => "0000010111001110",
17354 => "0000010111001110",
17355 => "0000010111001111",
17356 => "0000010111001111",
17357 => "0000010111001111",
17358 => "0000010111010000",
17359 => "0000010111010000",
17360 => "0000010111010000",
17361 => "0000010111010001",
17362 => "0000010111010001",
17363 => "0000010111010001",
17364 => "0000010111010010",
17365 => "0000010111010010",
17366 => "0000010111010010",
17367 => "0000010111010011",
17368 => "0000010111010011",
17369 => "0000010111010011",
17370 => "0000010111010100",
17371 => "0000010111010100",
17372 => "0000010111010101",
17373 => "0000010111010101",
17374 => "0000010111010101",
17375 => "0000010111010110",
17376 => "0000010111010110",
17377 => "0000010111010110",
17378 => "0000010111010111",
17379 => "0000010111010111",
17380 => "0000010111010111",
17381 => "0000010111011000",
17382 => "0000010111011000",
17383 => "0000010111011000",
17384 => "0000010111011001",
17385 => "0000010111011001",
17386 => "0000010111011010",
17387 => "0000010111011010",
17388 => "0000010111011010",
17389 => "0000010111011011",
17390 => "0000010111011011",
17391 => "0000010111011011",
17392 => "0000010111011100",
17393 => "0000010111011100",
17394 => "0000010111011100",
17395 => "0000010111011101",
17396 => "0000010111011101",
17397 => "0000010111011101",
17398 => "0000010111011110",
17399 => "0000010111011110",
17400 => "0000010111011111",
17401 => "0000010111011111",
17402 => "0000010111011111",
17403 => "0000010111100000",
17404 => "0000010111100000",
17405 => "0000010111100000",
17406 => "0000010111100001",
17407 => "0000010111100001",
17408 => "0000010111100001",
17409 => "0000010111100010",
17410 => "0000010111100010",
17411 => "0000010111100011",
17412 => "0000010111100011",
17413 => "0000010111100011",
17414 => "0000010111100100",
17415 => "0000010111100100",
17416 => "0000010111100100",
17417 => "0000010111100101",
17418 => "0000010111100101",
17419 => "0000010111100101",
17420 => "0000010111100110",
17421 => "0000010111100110",
17422 => "0000010111100110",
17423 => "0000010111100111",
17424 => "0000010111100111",
17425 => "0000010111101000",
17426 => "0000010111101000",
17427 => "0000010111101000",
17428 => "0000010111101001",
17429 => "0000010111101001",
17430 => "0000010111101001",
17431 => "0000010111101010",
17432 => "0000010111101010",
17433 => "0000010111101010",
17434 => "0000010111101011",
17435 => "0000010111101011",
17436 => "0000010111101100",
17437 => "0000010111101100",
17438 => "0000010111101100",
17439 => "0000010111101101",
17440 => "0000010111101101",
17441 => "0000010111101101",
17442 => "0000010111101110",
17443 => "0000010111101110",
17444 => "0000010111101110",
17445 => "0000010111101111",
17446 => "0000010111101111",
17447 => "0000010111110000",
17448 => "0000010111110000",
17449 => "0000010111110000",
17450 => "0000010111110001",
17451 => "0000010111110001",
17452 => "0000010111110001",
17453 => "0000010111110010",
17454 => "0000010111110010",
17455 => "0000010111110010",
17456 => "0000010111110011",
17457 => "0000010111110011",
17458 => "0000010111110100",
17459 => "0000010111110100",
17460 => "0000010111110100",
17461 => "0000010111110101",
17462 => "0000010111110101",
17463 => "0000010111110101",
17464 => "0000010111110110",
17465 => "0000010111110110",
17466 => "0000010111110110",
17467 => "0000010111110111",
17468 => "0000010111110111",
17469 => "0000010111111000",
17470 => "0000010111111000",
17471 => "0000010111111000",
17472 => "0000010111111001",
17473 => "0000010111111001",
17474 => "0000010111111001",
17475 => "0000010111111010",
17476 => "0000010111111010",
17477 => "0000010111111010",
17478 => "0000010111111011",
17479 => "0000010111111011",
17480 => "0000010111111100",
17481 => "0000010111111100",
17482 => "0000010111111100",
17483 => "0000010111111101",
17484 => "0000010111111101",
17485 => "0000010111111101",
17486 => "0000010111111110",
17487 => "0000010111111110",
17488 => "0000010111111110",
17489 => "0000010111111111",
17490 => "0000010111111111",
17491 => "0000011000000000",
17492 => "0000011000000000",
17493 => "0000011000000000",
17494 => "0000011000000001",
17495 => "0000011000000001",
17496 => "0000011000000001",
17497 => "0000011000000010",
17498 => "0000011000000010",
17499 => "0000011000000010",
17500 => "0000011000000011",
17501 => "0000011000000011",
17502 => "0000011000000100",
17503 => "0000011000000100",
17504 => "0000011000000100",
17505 => "0000011000000101",
17506 => "0000011000000101",
17507 => "0000011000000101",
17508 => "0000011000000110",
17509 => "0000011000000110",
17510 => "0000011000000111",
17511 => "0000011000000111",
17512 => "0000011000000111",
17513 => "0000011000001000",
17514 => "0000011000001000",
17515 => "0000011000001000",
17516 => "0000011000001001",
17517 => "0000011000001001",
17518 => "0000011000001001",
17519 => "0000011000001010",
17520 => "0000011000001010",
17521 => "0000011000001011",
17522 => "0000011000001011",
17523 => "0000011000001011",
17524 => "0000011000001100",
17525 => "0000011000001100",
17526 => "0000011000001100",
17527 => "0000011000001101",
17528 => "0000011000001101",
17529 => "0000011000001110",
17530 => "0000011000001110",
17531 => "0000011000001110",
17532 => "0000011000001111",
17533 => "0000011000001111",
17534 => "0000011000001111",
17535 => "0000011000010000",
17536 => "0000011000010000",
17537 => "0000011000010000",
17538 => "0000011000010001",
17539 => "0000011000010001",
17540 => "0000011000010010",
17541 => "0000011000010010",
17542 => "0000011000010010",
17543 => "0000011000010011",
17544 => "0000011000010011",
17545 => "0000011000010011",
17546 => "0000011000010100",
17547 => "0000011000010100",
17548 => "0000011000010101",
17549 => "0000011000010101",
17550 => "0000011000010101",
17551 => "0000011000010110",
17552 => "0000011000010110",
17553 => "0000011000010110",
17554 => "0000011000010111",
17555 => "0000011000010111",
17556 => "0000011000011000",
17557 => "0000011000011000",
17558 => "0000011000011000",
17559 => "0000011000011001",
17560 => "0000011000011001",
17561 => "0000011000011001",
17562 => "0000011000011010",
17563 => "0000011000011010",
17564 => "0000011000011011",
17565 => "0000011000011011",
17566 => "0000011000011011",
17567 => "0000011000011100",
17568 => "0000011000011100",
17569 => "0000011000011100",
17570 => "0000011000011101",
17571 => "0000011000011101",
17572 => "0000011000011101",
17573 => "0000011000011110",
17574 => "0000011000011110",
17575 => "0000011000011111",
17576 => "0000011000011111",
17577 => "0000011000011111",
17578 => "0000011000100000",
17579 => "0000011000100000",
17580 => "0000011000100000",
17581 => "0000011000100001",
17582 => "0000011000100001",
17583 => "0000011000100010",
17584 => "0000011000100010",
17585 => "0000011000100010",
17586 => "0000011000100011",
17587 => "0000011000100011",
17588 => "0000011000100011",
17589 => "0000011000100100",
17590 => "0000011000100100",
17591 => "0000011000100101",
17592 => "0000011000100101",
17593 => "0000011000100101",
17594 => "0000011000100110",
17595 => "0000011000100110",
17596 => "0000011000100110",
17597 => "0000011000100111",
17598 => "0000011000100111",
17599 => "0000011000101000",
17600 => "0000011000101000",
17601 => "0000011000101000",
17602 => "0000011000101001",
17603 => "0000011000101001",
17604 => "0000011000101001",
17605 => "0000011000101010",
17606 => "0000011000101010",
17607 => "0000011000101011",
17608 => "0000011000101011",
17609 => "0000011000101011",
17610 => "0000011000101100",
17611 => "0000011000101100",
17612 => "0000011000101100",
17613 => "0000011000101101",
17614 => "0000011000101101",
17615 => "0000011000101110",
17616 => "0000011000101110",
17617 => "0000011000101110",
17618 => "0000011000101111",
17619 => "0000011000101111",
17620 => "0000011000110000",
17621 => "0000011000110000",
17622 => "0000011000110000",
17623 => "0000011000110001",
17624 => "0000011000110001",
17625 => "0000011000110001",
17626 => "0000011000110010",
17627 => "0000011000110010",
17628 => "0000011000110011",
17629 => "0000011000110011",
17630 => "0000011000110011",
17631 => "0000011000110100",
17632 => "0000011000110100",
17633 => "0000011000110100",
17634 => "0000011000110101",
17635 => "0000011000110101",
17636 => "0000011000110110",
17637 => "0000011000110110",
17638 => "0000011000110110",
17639 => "0000011000110111",
17640 => "0000011000110111",
17641 => "0000011000110111",
17642 => "0000011000111000",
17643 => "0000011000111000",
17644 => "0000011000111001",
17645 => "0000011000111001",
17646 => "0000011000111001",
17647 => "0000011000111010",
17648 => "0000011000111010",
17649 => "0000011000111010",
17650 => "0000011000111011",
17651 => "0000011000111011",
17652 => "0000011000111100",
17653 => "0000011000111100",
17654 => "0000011000111100",
17655 => "0000011000111101",
17656 => "0000011000111101",
17657 => "0000011000111110",
17658 => "0000011000111110",
17659 => "0000011000111110",
17660 => "0000011000111111",
17661 => "0000011000111111",
17662 => "0000011000111111",
17663 => "0000011001000000",
17664 => "0000011001000000",
17665 => "0000011001000001",
17666 => "0000011001000001",
17667 => "0000011001000001",
17668 => "0000011001000010",
17669 => "0000011001000010",
17670 => "0000011001000010",
17671 => "0000011001000011",
17672 => "0000011001000011",
17673 => "0000011001000100",
17674 => "0000011001000100",
17675 => "0000011001000100",
17676 => "0000011001000101",
17677 => "0000011001000101",
17678 => "0000011001000110",
17679 => "0000011001000110",
17680 => "0000011001000110",
17681 => "0000011001000111",
17682 => "0000011001000111",
17683 => "0000011001000111",
17684 => "0000011001001000",
17685 => "0000011001001000",
17686 => "0000011001001001",
17687 => "0000011001001001",
17688 => "0000011001001001",
17689 => "0000011001001010",
17690 => "0000011001001010",
17691 => "0000011001001011",
17692 => "0000011001001011",
17693 => "0000011001001011",
17694 => "0000011001001100",
17695 => "0000011001001100",
17696 => "0000011001001100",
17697 => "0000011001001101",
17698 => "0000011001001101",
17699 => "0000011001001110",
17700 => "0000011001001110",
17701 => "0000011001001110",
17702 => "0000011001001111",
17703 => "0000011001001111",
17704 => "0000011001010000",
17705 => "0000011001010000",
17706 => "0000011001010000",
17707 => "0000011001010001",
17708 => "0000011001010001",
17709 => "0000011001010001",
17710 => "0000011001010010",
17711 => "0000011001010010",
17712 => "0000011001010011",
17713 => "0000011001010011",
17714 => "0000011001010011",
17715 => "0000011001010100",
17716 => "0000011001010100",
17717 => "0000011001010101",
17718 => "0000011001010101",
17719 => "0000011001010101",
17720 => "0000011001010110",
17721 => "0000011001010110",
17722 => "0000011001010110",
17723 => "0000011001010111",
17724 => "0000011001010111",
17725 => "0000011001011000",
17726 => "0000011001011000",
17727 => "0000011001011000",
17728 => "0000011001011001",
17729 => "0000011001011001",
17730 => "0000011001011010",
17731 => "0000011001011010",
17732 => "0000011001011010",
17733 => "0000011001011011",
17734 => "0000011001011011",
17735 => "0000011001011011",
17736 => "0000011001011100",
17737 => "0000011001011100",
17738 => "0000011001011101",
17739 => "0000011001011101",
17740 => "0000011001011101",
17741 => "0000011001011110",
17742 => "0000011001011110",
17743 => "0000011001011111",
17744 => "0000011001011111",
17745 => "0000011001011111",
17746 => "0000011001100000",
17747 => "0000011001100000",
17748 => "0000011001100001",
17749 => "0000011001100001",
17750 => "0000011001100001",
17751 => "0000011001100010",
17752 => "0000011001100010",
17753 => "0000011001100010",
17754 => "0000011001100011",
17755 => "0000011001100011",
17756 => "0000011001100100",
17757 => "0000011001100100",
17758 => "0000011001100100",
17759 => "0000011001100101",
17760 => "0000011001100101",
17761 => "0000011001100110",
17762 => "0000011001100110",
17763 => "0000011001100110",
17764 => "0000011001100111",
17765 => "0000011001100111",
17766 => "0000011001101000",
17767 => "0000011001101000",
17768 => "0000011001101000",
17769 => "0000011001101001",
17770 => "0000011001101001",
17771 => "0000011001101001",
17772 => "0000011001101010",
17773 => "0000011001101010",
17774 => "0000011001101011",
17775 => "0000011001101011",
17776 => "0000011001101011",
17777 => "0000011001101100",
17778 => "0000011001101100",
17779 => "0000011001101101",
17780 => "0000011001101101",
17781 => "0000011001101101",
17782 => "0000011001101110",
17783 => "0000011001101110",
17784 => "0000011001101111",
17785 => "0000011001101111",
17786 => "0000011001101111",
17787 => "0000011001110000",
17788 => "0000011001110000",
17789 => "0000011001110001",
17790 => "0000011001110001",
17791 => "0000011001110001",
17792 => "0000011001110010",
17793 => "0000011001110010",
17794 => "0000011001110011",
17795 => "0000011001110011",
17796 => "0000011001110011",
17797 => "0000011001110100",
17798 => "0000011001110100",
17799 => "0000011001110100",
17800 => "0000011001110101",
17801 => "0000011001110101",
17802 => "0000011001110110",
17803 => "0000011001110110",
17804 => "0000011001110110",
17805 => "0000011001110111",
17806 => "0000011001110111",
17807 => "0000011001111000",
17808 => "0000011001111000",
17809 => "0000011001111000",
17810 => "0000011001111001",
17811 => "0000011001111001",
17812 => "0000011001111010",
17813 => "0000011001111010",
17814 => "0000011001111010",
17815 => "0000011001111011",
17816 => "0000011001111011",
17817 => "0000011001111100",
17818 => "0000011001111100",
17819 => "0000011001111100",
17820 => "0000011001111101",
17821 => "0000011001111101",
17822 => "0000011001111110",
17823 => "0000011001111110",
17824 => "0000011001111110",
17825 => "0000011001111111",
17826 => "0000011001111111",
17827 => "0000011010000000",
17828 => "0000011010000000",
17829 => "0000011010000000",
17830 => "0000011010000001",
17831 => "0000011010000001",
17832 => "0000011010000010",
17833 => "0000011010000010",
17834 => "0000011010000010",
17835 => "0000011010000011",
17836 => "0000011010000011",
17837 => "0000011010000011",
17838 => "0000011010000100",
17839 => "0000011010000100",
17840 => "0000011010000101",
17841 => "0000011010000101",
17842 => "0000011010000101",
17843 => "0000011010000110",
17844 => "0000011010000110",
17845 => "0000011010000111",
17846 => "0000011010000111",
17847 => "0000011010000111",
17848 => "0000011010001000",
17849 => "0000011010001000",
17850 => "0000011010001001",
17851 => "0000011010001001",
17852 => "0000011010001001",
17853 => "0000011010001010",
17854 => "0000011010001010",
17855 => "0000011010001011",
17856 => "0000011010001011",
17857 => "0000011010001011",
17858 => "0000011010001100",
17859 => "0000011010001100",
17860 => "0000011010001101",
17861 => "0000011010001101",
17862 => "0000011010001101",
17863 => "0000011010001110",
17864 => "0000011010001110",
17865 => "0000011010001111",
17866 => "0000011010001111",
17867 => "0000011010001111",
17868 => "0000011010010000",
17869 => "0000011010010000",
17870 => "0000011010010001",
17871 => "0000011010010001",
17872 => "0000011010010001",
17873 => "0000011010010010",
17874 => "0000011010010010",
17875 => "0000011010010011",
17876 => "0000011010010011",
17877 => "0000011010010011",
17878 => "0000011010010100",
17879 => "0000011010010100",
17880 => "0000011010010101",
17881 => "0000011010010101",
17882 => "0000011010010101",
17883 => "0000011010010110",
17884 => "0000011010010110",
17885 => "0000011010010111",
17886 => "0000011010010111",
17887 => "0000011010010111",
17888 => "0000011010011000",
17889 => "0000011010011000",
17890 => "0000011010011001",
17891 => "0000011010011001",
17892 => "0000011010011001",
17893 => "0000011010011010",
17894 => "0000011010011010",
17895 => "0000011010011011",
17896 => "0000011010011011",
17897 => "0000011010011011",
17898 => "0000011010011100",
17899 => "0000011010011100",
17900 => "0000011010011101",
17901 => "0000011010011101",
17902 => "0000011010011101",
17903 => "0000011010011110",
17904 => "0000011010011110",
17905 => "0000011010011111",
17906 => "0000011010011111",
17907 => "0000011010100000",
17908 => "0000011010100000",
17909 => "0000011010100000",
17910 => "0000011010100001",
17911 => "0000011010100001",
17912 => "0000011010100010",
17913 => "0000011010100010",
17914 => "0000011010100010",
17915 => "0000011010100011",
17916 => "0000011010100011",
17917 => "0000011010100100",
17918 => "0000011010100100",
17919 => "0000011010100100",
17920 => "0000011010100101",
17921 => "0000011010100101",
17922 => "0000011010100110",
17923 => "0000011010100110",
17924 => "0000011010100110",
17925 => "0000011010100111",
17926 => "0000011010100111",
17927 => "0000011010101000",
17928 => "0000011010101000",
17929 => "0000011010101000",
17930 => "0000011010101001",
17931 => "0000011010101001",
17932 => "0000011010101010",
17933 => "0000011010101010",
17934 => "0000011010101010",
17935 => "0000011010101011",
17936 => "0000011010101011",
17937 => "0000011010101100",
17938 => "0000011010101100",
17939 => "0000011010101100",
17940 => "0000011010101101",
17941 => "0000011010101101",
17942 => "0000011010101110",
17943 => "0000011010101110",
17944 => "0000011010101110",
17945 => "0000011010101111",
17946 => "0000011010101111",
17947 => "0000011010110000",
17948 => "0000011010110000",
17949 => "0000011010110001",
17950 => "0000011010110001",
17951 => "0000011010110001",
17952 => "0000011010110010",
17953 => "0000011010110010",
17954 => "0000011010110011",
17955 => "0000011010110011",
17956 => "0000011010110011",
17957 => "0000011010110100",
17958 => "0000011010110100",
17959 => "0000011010110101",
17960 => "0000011010110101",
17961 => "0000011010110101",
17962 => "0000011010110110",
17963 => "0000011010110110",
17964 => "0000011010110111",
17965 => "0000011010110111",
17966 => "0000011010110111",
17967 => "0000011010111000",
17968 => "0000011010111000",
17969 => "0000011010111001",
17970 => "0000011010111001",
17971 => "0000011010111010",
17972 => "0000011010111010",
17973 => "0000011010111010",
17974 => "0000011010111011",
17975 => "0000011010111011",
17976 => "0000011010111100",
17977 => "0000011010111100",
17978 => "0000011010111100",
17979 => "0000011010111101",
17980 => "0000011010111101",
17981 => "0000011010111110",
17982 => "0000011010111110",
17983 => "0000011010111110",
17984 => "0000011010111111",
17985 => "0000011010111111",
17986 => "0000011011000000",
17987 => "0000011011000000",
17988 => "0000011011000000",
17989 => "0000011011000001",
17990 => "0000011011000001",
17991 => "0000011011000010",
17992 => "0000011011000010",
17993 => "0000011011000011",
17994 => "0000011011000011",
17995 => "0000011011000011",
17996 => "0000011011000100",
17997 => "0000011011000100",
17998 => "0000011011000101",
17999 => "0000011011000101",
18000 => "0000011011000101",
18001 => "0000011011000110",
18002 => "0000011011000110",
18003 => "0000011011000111",
18004 => "0000011011000111",
18005 => "0000011011000111",
18006 => "0000011011001000",
18007 => "0000011011001000",
18008 => "0000011011001001",
18009 => "0000011011001001",
18010 => "0000011011001010",
18011 => "0000011011001010",
18012 => "0000011011001010",
18013 => "0000011011001011",
18014 => "0000011011001011",
18015 => "0000011011001100",
18016 => "0000011011001100",
18017 => "0000011011001100",
18018 => "0000011011001101",
18019 => "0000011011001101",
18020 => "0000011011001110",
18021 => "0000011011001110",
18022 => "0000011011001111",
18023 => "0000011011001111",
18024 => "0000011011001111",
18025 => "0000011011010000",
18026 => "0000011011010000",
18027 => "0000011011010001",
18028 => "0000011011010001",
18029 => "0000011011010001",
18030 => "0000011011010010",
18031 => "0000011011010010",
18032 => "0000011011010011",
18033 => "0000011011010011",
18034 => "0000011011010011",
18035 => "0000011011010100",
18036 => "0000011011010100",
18037 => "0000011011010101",
18038 => "0000011011010101",
18039 => "0000011011010110",
18040 => "0000011011010110",
18041 => "0000011011010110",
18042 => "0000011011010111",
18043 => "0000011011010111",
18044 => "0000011011011000",
18045 => "0000011011011000",
18046 => "0000011011011000",
18047 => "0000011011011001",
18048 => "0000011011011001",
18049 => "0000011011011010",
18050 => "0000011011011010",
18051 => "0000011011011011",
18052 => "0000011011011011",
18053 => "0000011011011011",
18054 => "0000011011011100",
18055 => "0000011011011100",
18056 => "0000011011011101",
18057 => "0000011011011101",
18058 => "0000011011011101",
18059 => "0000011011011110",
18060 => "0000011011011110",
18061 => "0000011011011111",
18062 => "0000011011011111",
18063 => "0000011011100000",
18064 => "0000011011100000",
18065 => "0000011011100000",
18066 => "0000011011100001",
18067 => "0000011011100001",
18068 => "0000011011100010",
18069 => "0000011011100010",
18070 => "0000011011100011",
18071 => "0000011011100011",
18072 => "0000011011100011",
18073 => "0000011011100100",
18074 => "0000011011100100",
18075 => "0000011011100101",
18076 => "0000011011100101",
18077 => "0000011011100101",
18078 => "0000011011100110",
18079 => "0000011011100110",
18080 => "0000011011100111",
18081 => "0000011011100111",
18082 => "0000011011101000",
18083 => "0000011011101000",
18084 => "0000011011101000",
18085 => "0000011011101001",
18086 => "0000011011101001",
18087 => "0000011011101010",
18088 => "0000011011101010",
18089 => "0000011011101010",
18090 => "0000011011101011",
18091 => "0000011011101011",
18092 => "0000011011101100",
18093 => "0000011011101100",
18094 => "0000011011101101",
18095 => "0000011011101101",
18096 => "0000011011101101",
18097 => "0000011011101110",
18098 => "0000011011101110",
18099 => "0000011011101111",
18100 => "0000011011101111",
18101 => "0000011011110000",
18102 => "0000011011110000",
18103 => "0000011011110000",
18104 => "0000011011110001",
18105 => "0000011011110001",
18106 => "0000011011110010",
18107 => "0000011011110010",
18108 => "0000011011110010",
18109 => "0000011011110011",
18110 => "0000011011110011",
18111 => "0000011011110100",
18112 => "0000011011110100",
18113 => "0000011011110101",
18114 => "0000011011110101",
18115 => "0000011011110101",
18116 => "0000011011110110",
18117 => "0000011011110110",
18118 => "0000011011110111",
18119 => "0000011011110111",
18120 => "0000011011111000",
18121 => "0000011011111000",
18122 => "0000011011111000",
18123 => "0000011011111001",
18124 => "0000011011111001",
18125 => "0000011011111010",
18126 => "0000011011111010",
18127 => "0000011011111011",
18128 => "0000011011111011",
18129 => "0000011011111011",
18130 => "0000011011111100",
18131 => "0000011011111100",
18132 => "0000011011111101",
18133 => "0000011011111101",
18134 => "0000011011111110",
18135 => "0000011011111110",
18136 => "0000011011111110",
18137 => "0000011011111111",
18138 => "0000011011111111",
18139 => "0000011100000000",
18140 => "0000011100000000",
18141 => "0000011100000000",
18142 => "0000011100000001",
18143 => "0000011100000001",
18144 => "0000011100000010",
18145 => "0000011100000010",
18146 => "0000011100000011",
18147 => "0000011100000011",
18148 => "0000011100000011",
18149 => "0000011100000100",
18150 => "0000011100000100",
18151 => "0000011100000101",
18152 => "0000011100000101",
18153 => "0000011100000110",
18154 => "0000011100000110",
18155 => "0000011100000110",
18156 => "0000011100000111",
18157 => "0000011100000111",
18158 => "0000011100001000",
18159 => "0000011100001000",
18160 => "0000011100001001",
18161 => "0000011100001001",
18162 => "0000011100001001",
18163 => "0000011100001010",
18164 => "0000011100001010",
18165 => "0000011100001011",
18166 => "0000011100001011",
18167 => "0000011100001100",
18168 => "0000011100001100",
18169 => "0000011100001100",
18170 => "0000011100001101",
18171 => "0000011100001101",
18172 => "0000011100001110",
18173 => "0000011100001110",
18174 => "0000011100001111",
18175 => "0000011100001111",
18176 => "0000011100001111",
18177 => "0000011100010000",
18178 => "0000011100010000",
18179 => "0000011100010001",
18180 => "0000011100010001",
18181 => "0000011100010010",
18182 => "0000011100010010",
18183 => "0000011100010010",
18184 => "0000011100010011",
18185 => "0000011100010011",
18186 => "0000011100010100",
18187 => "0000011100010100",
18188 => "0000011100010101",
18189 => "0000011100010101",
18190 => "0000011100010101",
18191 => "0000011100010110",
18192 => "0000011100010110",
18193 => "0000011100010111",
18194 => "0000011100010111",
18195 => "0000011100011000",
18196 => "0000011100011000",
18197 => "0000011100011000",
18198 => "0000011100011001",
18199 => "0000011100011001",
18200 => "0000011100011010",
18201 => "0000011100011010",
18202 => "0000011100011011",
18203 => "0000011100011011",
18204 => "0000011100011100",
18205 => "0000011100011100",
18206 => "0000011100011100",
18207 => "0000011100011101",
18208 => "0000011100011101",
18209 => "0000011100011110",
18210 => "0000011100011110",
18211 => "0000011100011111",
18212 => "0000011100011111",
18213 => "0000011100011111",
18214 => "0000011100100000",
18215 => "0000011100100000",
18216 => "0000011100100001",
18217 => "0000011100100001",
18218 => "0000011100100010",
18219 => "0000011100100010",
18220 => "0000011100100010",
18221 => "0000011100100011",
18222 => "0000011100100011",
18223 => "0000011100100100",
18224 => "0000011100100100",
18225 => "0000011100100101",
18226 => "0000011100100101",
18227 => "0000011100100101",
18228 => "0000011100100110",
18229 => "0000011100100110",
18230 => "0000011100100111",
18231 => "0000011100100111",
18232 => "0000011100101000",
18233 => "0000011100101000",
18234 => "0000011100101001",
18235 => "0000011100101001",
18236 => "0000011100101001",
18237 => "0000011100101010",
18238 => "0000011100101010",
18239 => "0000011100101011",
18240 => "0000011100101011",
18241 => "0000011100101100",
18242 => "0000011100101100",
18243 => "0000011100101100",
18244 => "0000011100101101",
18245 => "0000011100101101",
18246 => "0000011100101110",
18247 => "0000011100101110",
18248 => "0000011100101111",
18249 => "0000011100101111",
18250 => "0000011100101111",
18251 => "0000011100110000",
18252 => "0000011100110000",
18253 => "0000011100110001",
18254 => "0000011100110001",
18255 => "0000011100110010",
18256 => "0000011100110010",
18257 => "0000011100110011",
18258 => "0000011100110011",
18259 => "0000011100110011",
18260 => "0000011100110100",
18261 => "0000011100110100",
18262 => "0000011100110101",
18263 => "0000011100110101",
18264 => "0000011100110110",
18265 => "0000011100110110",
18266 => "0000011100110110",
18267 => "0000011100110111",
18268 => "0000011100110111",
18269 => "0000011100111000",
18270 => "0000011100111000",
18271 => "0000011100111001",
18272 => "0000011100111001",
18273 => "0000011100111010",
18274 => "0000011100111010",
18275 => "0000011100111010",
18276 => "0000011100111011",
18277 => "0000011100111011",
18278 => "0000011100111100",
18279 => "0000011100111100",
18280 => "0000011100111101",
18281 => "0000011100111101",
18282 => "0000011100111110",
18283 => "0000011100111110",
18284 => "0000011100111110",
18285 => "0000011100111111",
18286 => "0000011100111111",
18287 => "0000011101000000",
18288 => "0000011101000000",
18289 => "0000011101000001",
18290 => "0000011101000001",
18291 => "0000011101000001",
18292 => "0000011101000010",
18293 => "0000011101000010",
18294 => "0000011101000011",
18295 => "0000011101000011",
18296 => "0000011101000100",
18297 => "0000011101000100",
18298 => "0000011101000101",
18299 => "0000011101000101",
18300 => "0000011101000101",
18301 => "0000011101000110",
18302 => "0000011101000110",
18303 => "0000011101000111",
18304 => "0000011101000111",
18305 => "0000011101001000",
18306 => "0000011101001000",
18307 => "0000011101001001",
18308 => "0000011101001001",
18309 => "0000011101001001",
18310 => "0000011101001010",
18311 => "0000011101001010",
18312 => "0000011101001011",
18313 => "0000011101001011",
18314 => "0000011101001100",
18315 => "0000011101001100",
18316 => "0000011101001101",
18317 => "0000011101001101",
18318 => "0000011101001101",
18319 => "0000011101001110",
18320 => "0000011101001110",
18321 => "0000011101001111",
18322 => "0000011101001111",
18323 => "0000011101010000",
18324 => "0000011101010000",
18325 => "0000011101010001",
18326 => "0000011101010001",
18327 => "0000011101010001",
18328 => "0000011101010010",
18329 => "0000011101010010",
18330 => "0000011101010011",
18331 => "0000011101010011",
18332 => "0000011101010100",
18333 => "0000011101010100",
18334 => "0000011101010101",
18335 => "0000011101010101",
18336 => "0000011101010101",
18337 => "0000011101010110",
18338 => "0000011101010110",
18339 => "0000011101010111",
18340 => "0000011101010111",
18341 => "0000011101011000",
18342 => "0000011101011000",
18343 => "0000011101011001",
18344 => "0000011101011001",
18345 => "0000011101011001",
18346 => "0000011101011010",
18347 => "0000011101011010",
18348 => "0000011101011011",
18349 => "0000011101011011",
18350 => "0000011101011100",
18351 => "0000011101011100",
18352 => "0000011101011101",
18353 => "0000011101011101",
18354 => "0000011101011101",
18355 => "0000011101011110",
18356 => "0000011101011110",
18357 => "0000011101011111",
18358 => "0000011101011111",
18359 => "0000011101100000",
18360 => "0000011101100000",
18361 => "0000011101100001",
18362 => "0000011101100001",
18363 => "0000011101100001",
18364 => "0000011101100010",
18365 => "0000011101100010",
18366 => "0000011101100011",
18367 => "0000011101100011",
18368 => "0000011101100100",
18369 => "0000011101100100",
18370 => "0000011101100101",
18371 => "0000011101100101",
18372 => "0000011101100110",
18373 => "0000011101100110",
18374 => "0000011101100110",
18375 => "0000011101100111",
18376 => "0000011101100111",
18377 => "0000011101101000",
18378 => "0000011101101000",
18379 => "0000011101101001",
18380 => "0000011101101001",
18381 => "0000011101101010",
18382 => "0000011101101010",
18383 => "0000011101101010",
18384 => "0000011101101011",
18385 => "0000011101101011",
18386 => "0000011101101100",
18387 => "0000011101101100",
18388 => "0000011101101101",
18389 => "0000011101101101",
18390 => "0000011101101110",
18391 => "0000011101101110",
18392 => "0000011101101111",
18393 => "0000011101101111",
18394 => "0000011101101111",
18395 => "0000011101110000",
18396 => "0000011101110000",
18397 => "0000011101110001",
18398 => "0000011101110001",
18399 => "0000011101110010",
18400 => "0000011101110010",
18401 => "0000011101110011",
18402 => "0000011101110011",
18403 => "0000011101110011",
18404 => "0000011101110100",
18405 => "0000011101110100",
18406 => "0000011101110101",
18407 => "0000011101110101",
18408 => "0000011101110110",
18409 => "0000011101110110",
18410 => "0000011101110111",
18411 => "0000011101110111",
18412 => "0000011101111000",
18413 => "0000011101111000",
18414 => "0000011101111000",
18415 => "0000011101111001",
18416 => "0000011101111001",
18417 => "0000011101111010",
18418 => "0000011101111010",
18419 => "0000011101111011",
18420 => "0000011101111011",
18421 => "0000011101111100",
18422 => "0000011101111100",
18423 => "0000011101111101",
18424 => "0000011101111101",
18425 => "0000011101111101",
18426 => "0000011101111110",
18427 => "0000011101111110",
18428 => "0000011101111111",
18429 => "0000011101111111",
18430 => "0000011110000000",
18431 => "0000011110000000",
18432 => "0000011110000001",
18433 => "0000011110000001",
18434 => "0000011110000010",
18435 => "0000011110000010",
18436 => "0000011110000010",
18437 => "0000011110000011",
18438 => "0000011110000011",
18439 => "0000011110000100",
18440 => "0000011110000100",
18441 => "0000011110000101",
18442 => "0000011110000101",
18443 => "0000011110000110",
18444 => "0000011110000110",
18445 => "0000011110000111",
18446 => "0000011110000111",
18447 => "0000011110000111",
18448 => "0000011110001000",
18449 => "0000011110001000",
18450 => "0000011110001001",
18451 => "0000011110001001",
18452 => "0000011110001010",
18453 => "0000011110001010",
18454 => "0000011110001011",
18455 => "0000011110001011",
18456 => "0000011110001100",
18457 => "0000011110001100",
18458 => "0000011110001101",
18459 => "0000011110001101",
18460 => "0000011110001101",
18461 => "0000011110001110",
18462 => "0000011110001110",
18463 => "0000011110001111",
18464 => "0000011110001111",
18465 => "0000011110010000",
18466 => "0000011110010000",
18467 => "0000011110010001",
18468 => "0000011110010001",
18469 => "0000011110010010",
18470 => "0000011110010010",
18471 => "0000011110010010",
18472 => "0000011110010011",
18473 => "0000011110010011",
18474 => "0000011110010100",
18475 => "0000011110010100",
18476 => "0000011110010101",
18477 => "0000011110010101",
18478 => "0000011110010110",
18479 => "0000011110010110",
18480 => "0000011110010111",
18481 => "0000011110010111",
18482 => "0000011110011000",
18483 => "0000011110011000",
18484 => "0000011110011000",
18485 => "0000011110011001",
18486 => "0000011110011001",
18487 => "0000011110011010",
18488 => "0000011110011010",
18489 => "0000011110011011",
18490 => "0000011110011011",
18491 => "0000011110011100",
18492 => "0000011110011100",
18493 => "0000011110011101",
18494 => "0000011110011101",
18495 => "0000011110011110",
18496 => "0000011110011110",
18497 => "0000011110011110",
18498 => "0000011110011111",
18499 => "0000011110011111",
18500 => "0000011110100000",
18501 => "0000011110100000",
18502 => "0000011110100001",
18503 => "0000011110100001",
18504 => "0000011110100010",
18505 => "0000011110100010",
18506 => "0000011110100011",
18507 => "0000011110100011",
18508 => "0000011110100100",
18509 => "0000011110100100",
18510 => "0000011110100100",
18511 => "0000011110100101",
18512 => "0000011110100101",
18513 => "0000011110100110",
18514 => "0000011110100110",
18515 => "0000011110100111",
18516 => "0000011110100111",
18517 => "0000011110101000",
18518 => "0000011110101000",
18519 => "0000011110101001",
18520 => "0000011110101001",
18521 => "0000011110101010",
18522 => "0000011110101010",
18523 => "0000011110101011",
18524 => "0000011110101011",
18525 => "0000011110101011",
18526 => "0000011110101100",
18527 => "0000011110101100",
18528 => "0000011110101101",
18529 => "0000011110101101",
18530 => "0000011110101110",
18531 => "0000011110101110",
18532 => "0000011110101111",
18533 => "0000011110101111",
18534 => "0000011110110000",
18535 => "0000011110110000",
18536 => "0000011110110001",
18537 => "0000011110110001",
18538 => "0000011110110001",
18539 => "0000011110110010",
18540 => "0000011110110010",
18541 => "0000011110110011",
18542 => "0000011110110011",
18543 => "0000011110110100",
18544 => "0000011110110100",
18545 => "0000011110110101",
18546 => "0000011110110101",
18547 => "0000011110110110",
18548 => "0000011110110110",
18549 => "0000011110110111",
18550 => "0000011110110111",
18551 => "0000011110111000",
18552 => "0000011110111000",
18553 => "0000011110111000",
18554 => "0000011110111001",
18555 => "0000011110111001",
18556 => "0000011110111010",
18557 => "0000011110111010",
18558 => "0000011110111011",
18559 => "0000011110111011",
18560 => "0000011110111100",
18561 => "0000011110111100",
18562 => "0000011110111101",
18563 => "0000011110111101",
18564 => "0000011110111110",
18565 => "0000011110111110",
18566 => "0000011110111111",
18567 => "0000011110111111",
18568 => "0000011111000000",
18569 => "0000011111000000",
18570 => "0000011111000000",
18571 => "0000011111000001",
18572 => "0000011111000001",
18573 => "0000011111000010",
18574 => "0000011111000010",
18575 => "0000011111000011",
18576 => "0000011111000011",
18577 => "0000011111000100",
18578 => "0000011111000100",
18579 => "0000011111000101",
18580 => "0000011111000101",
18581 => "0000011111000110",
18582 => "0000011111000110",
18583 => "0000011111000111",
18584 => "0000011111000111",
18585 => "0000011111001000",
18586 => "0000011111001000",
18587 => "0000011111001000",
18588 => "0000011111001001",
18589 => "0000011111001001",
18590 => "0000011111001010",
18591 => "0000011111001010",
18592 => "0000011111001011",
18593 => "0000011111001011",
18594 => "0000011111001100",
18595 => "0000011111001100",
18596 => "0000011111001101",
18597 => "0000011111001101",
18598 => "0000011111001110",
18599 => "0000011111001110",
18600 => "0000011111001111",
18601 => "0000011111001111",
18602 => "0000011111010000",
18603 => "0000011111010000",
18604 => "0000011111010001",
18605 => "0000011111010001",
18606 => "0000011111010001",
18607 => "0000011111010010",
18608 => "0000011111010010",
18609 => "0000011111010011",
18610 => "0000011111010011",
18611 => "0000011111010100",
18612 => "0000011111010100",
18613 => "0000011111010101",
18614 => "0000011111010101",
18615 => "0000011111010110",
18616 => "0000011111010110",
18617 => "0000011111010111",
18618 => "0000011111010111",
18619 => "0000011111011000",
18620 => "0000011111011000",
18621 => "0000011111011001",
18622 => "0000011111011001",
18623 => "0000011111011010",
18624 => "0000011111011010",
18625 => "0000011111011010",
18626 => "0000011111011011",
18627 => "0000011111011011",
18628 => "0000011111011100",
18629 => "0000011111011100",
18630 => "0000011111011101",
18631 => "0000011111011101",
18632 => "0000011111011110",
18633 => "0000011111011110",
18634 => "0000011111011111",
18635 => "0000011111011111",
18636 => "0000011111100000",
18637 => "0000011111100000",
18638 => "0000011111100001",
18639 => "0000011111100001",
18640 => "0000011111100010",
18641 => "0000011111100010",
18642 => "0000011111100011",
18643 => "0000011111100011",
18644 => "0000011111100100",
18645 => "0000011111100100",
18646 => "0000011111100100",
18647 => "0000011111100101",
18648 => "0000011111100101",
18649 => "0000011111100110",
18650 => "0000011111100110",
18651 => "0000011111100111",
18652 => "0000011111100111",
18653 => "0000011111101000",
18654 => "0000011111101000",
18655 => "0000011111101001",
18656 => "0000011111101001",
18657 => "0000011111101010",
18658 => "0000011111101010",
18659 => "0000011111101011",
18660 => "0000011111101011",
18661 => "0000011111101100",
18662 => "0000011111101100",
18663 => "0000011111101101",
18664 => "0000011111101101",
18665 => "0000011111101110",
18666 => "0000011111101110",
18667 => "0000011111101111",
18668 => "0000011111101111",
18669 => "0000011111110000",
18670 => "0000011111110000",
18671 => "0000011111110000",
18672 => "0000011111110001",
18673 => "0000011111110001",
18674 => "0000011111110010",
18675 => "0000011111110010",
18676 => "0000011111110011",
18677 => "0000011111110011",
18678 => "0000011111110100",
18679 => "0000011111110100",
18680 => "0000011111110101",
18681 => "0000011111110101",
18682 => "0000011111110110",
18683 => "0000011111110110",
18684 => "0000011111110111",
18685 => "0000011111110111",
18686 => "0000011111111000",
18687 => "0000011111111000",
18688 => "0000011111111001",
18689 => "0000011111111001",
18690 => "0000011111111010",
18691 => "0000011111111010",
18692 => "0000011111111011",
18693 => "0000011111111011",
18694 => "0000011111111100",
18695 => "0000011111111100",
18696 => "0000011111111101",
18697 => "0000011111111101",
18698 => "0000011111111110",
18699 => "0000011111111110",
18700 => "0000011111111110",
18701 => "0000011111111111",
18702 => "0000011111111111",
18703 => "0000100000000000",
18704 => "0000100000000000",
18705 => "0000100000000001",
18706 => "0000100000000001",
18707 => "0000100000000010",
18708 => "0000100000000010",
18709 => "0000100000000011",
18710 => "0000100000000011",
18711 => "0000100000000100",
18712 => "0000100000000100",
18713 => "0000100000000101",
18714 => "0000100000000101",
18715 => "0000100000000110",
18716 => "0000100000000110",
18717 => "0000100000000111",
18718 => "0000100000000111",
18719 => "0000100000001000",
18720 => "0000100000001000",
18721 => "0000100000001001",
18722 => "0000100000001001",
18723 => "0000100000001010",
18724 => "0000100000001010",
18725 => "0000100000001011",
18726 => "0000100000001011",
18727 => "0000100000001100",
18728 => "0000100000001100",
18729 => "0000100000001101",
18730 => "0000100000001101",
18731 => "0000100000001110",
18732 => "0000100000001110",
18733 => "0000100000001111",
18734 => "0000100000001111",
18735 => "0000100000001111",
18736 => "0000100000010000",
18737 => "0000100000010000",
18738 => "0000100000010001",
18739 => "0000100000010001",
18740 => "0000100000010010",
18741 => "0000100000010010",
18742 => "0000100000010011",
18743 => "0000100000010011",
18744 => "0000100000010100",
18745 => "0000100000010100",
18746 => "0000100000010101",
18747 => "0000100000010101",
18748 => "0000100000010110",
18749 => "0000100000010110",
18750 => "0000100000010111",
18751 => "0000100000010111",
18752 => "0000100000011000",
18753 => "0000100000011000",
18754 => "0000100000011001",
18755 => "0000100000011001",
18756 => "0000100000011010",
18757 => "0000100000011010",
18758 => "0000100000011011",
18759 => "0000100000011011",
18760 => "0000100000011100",
18761 => "0000100000011100",
18762 => "0000100000011101",
18763 => "0000100000011101",
18764 => "0000100000011110",
18765 => "0000100000011110",
18766 => "0000100000011111",
18767 => "0000100000011111",
18768 => "0000100000100000",
18769 => "0000100000100000",
18770 => "0000100000100001",
18771 => "0000100000100001",
18772 => "0000100000100010",
18773 => "0000100000100010",
18774 => "0000100000100011",
18775 => "0000100000100011",
18776 => "0000100000100100",
18777 => "0000100000100100",
18778 => "0000100000100101",
18779 => "0000100000100101",
18780 => "0000100000100110",
18781 => "0000100000100110",
18782 => "0000100000100111",
18783 => "0000100000100111",
18784 => "0000100000101000",
18785 => "0000100000101000",
18786 => "0000100000101001",
18787 => "0000100000101001",
18788 => "0000100000101010",
18789 => "0000100000101010",
18790 => "0000100000101011",
18791 => "0000100000101011",
18792 => "0000100000101011",
18793 => "0000100000101100",
18794 => "0000100000101100",
18795 => "0000100000101101",
18796 => "0000100000101101",
18797 => "0000100000101110",
18798 => "0000100000101110",
18799 => "0000100000101111",
18800 => "0000100000101111",
18801 => "0000100000110000",
18802 => "0000100000110000",
18803 => "0000100000110001",
18804 => "0000100000110001",
18805 => "0000100000110010",
18806 => "0000100000110010",
18807 => "0000100000110011",
18808 => "0000100000110011",
18809 => "0000100000110100",
18810 => "0000100000110100",
18811 => "0000100000110101",
18812 => "0000100000110101",
18813 => "0000100000110110",
18814 => "0000100000110110",
18815 => "0000100000110111",
18816 => "0000100000110111",
18817 => "0000100000111000",
18818 => "0000100000111000",
18819 => "0000100000111001",
18820 => "0000100000111001",
18821 => "0000100000111010",
18822 => "0000100000111010",
18823 => "0000100000111011",
18824 => "0000100000111011",
18825 => "0000100000111100",
18826 => "0000100000111100",
18827 => "0000100000111101",
18828 => "0000100000111101",
18829 => "0000100000111110",
18830 => "0000100000111110",
18831 => "0000100000111111",
18832 => "0000100000111111",
18833 => "0000100001000000",
18834 => "0000100001000000",
18835 => "0000100001000001",
18836 => "0000100001000001",
18837 => "0000100001000010",
18838 => "0000100001000010",
18839 => "0000100001000011",
18840 => "0000100001000011",
18841 => "0000100001000100",
18842 => "0000100001000100",
18843 => "0000100001000101",
18844 => "0000100001000101",
18845 => "0000100001000110",
18846 => "0000100001000110",
18847 => "0000100001000111",
18848 => "0000100001000111",
18849 => "0000100001001000",
18850 => "0000100001001000",
18851 => "0000100001001001",
18852 => "0000100001001001",
18853 => "0000100001001010",
18854 => "0000100001001010",
18855 => "0000100001001011",
18856 => "0000100001001011",
18857 => "0000100001001100",
18858 => "0000100001001100",
18859 => "0000100001001101",
18860 => "0000100001001101",
18861 => "0000100001001110",
18862 => "0000100001001110",
18863 => "0000100001001111",
18864 => "0000100001001111",
18865 => "0000100001010000",
18866 => "0000100001010000",
18867 => "0000100001010001",
18868 => "0000100001010001",
18869 => "0000100001010010",
18870 => "0000100001010010",
18871 => "0000100001010011",
18872 => "0000100001010011",
18873 => "0000100001010100",
18874 => "0000100001010100",
18875 => "0000100001010101",
18876 => "0000100001010101",
18877 => "0000100001010110",
18878 => "0000100001010110",
18879 => "0000100001010111",
18880 => "0000100001010111",
18881 => "0000100001011000",
18882 => "0000100001011000",
18883 => "0000100001011001",
18884 => "0000100001011001",
18885 => "0000100001011010",
18886 => "0000100001011010",
18887 => "0000100001011011",
18888 => "0000100001011011",
18889 => "0000100001011100",
18890 => "0000100001011100",
18891 => "0000100001011101",
18892 => "0000100001011110",
18893 => "0000100001011110",
18894 => "0000100001011111",
18895 => "0000100001011111",
18896 => "0000100001100000",
18897 => "0000100001100000",
18898 => "0000100001100001",
18899 => "0000100001100001",
18900 => "0000100001100010",
18901 => "0000100001100010",
18902 => "0000100001100011",
18903 => "0000100001100011",
18904 => "0000100001100100",
18905 => "0000100001100100",
18906 => "0000100001100101",
18907 => "0000100001100101",
18908 => "0000100001100110",
18909 => "0000100001100110",
18910 => "0000100001100111",
18911 => "0000100001100111",
18912 => "0000100001101000",
18913 => "0000100001101000",
18914 => "0000100001101001",
18915 => "0000100001101001",
18916 => "0000100001101010",
18917 => "0000100001101010",
18918 => "0000100001101011",
18919 => "0000100001101011",
18920 => "0000100001101100",
18921 => "0000100001101100",
18922 => "0000100001101101",
18923 => "0000100001101101",
18924 => "0000100001101110",
18925 => "0000100001101110",
18926 => "0000100001101111",
18927 => "0000100001101111",
18928 => "0000100001110000",
18929 => "0000100001110000",
18930 => "0000100001110001",
18931 => "0000100001110001",
18932 => "0000100001110010",
18933 => "0000100001110010",
18934 => "0000100001110011",
18935 => "0000100001110011",
18936 => "0000100001110100",
18937 => "0000100001110100",
18938 => "0000100001110101",
18939 => "0000100001110101",
18940 => "0000100001110110",
18941 => "0000100001110110",
18942 => "0000100001110111",
18943 => "0000100001110111",
18944 => "0000100001111000",
18945 => "0000100001111000",
18946 => "0000100001111001",
18947 => "0000100001111010",
18948 => "0000100001111010",
18949 => "0000100001111011",
18950 => "0000100001111011",
18951 => "0000100001111100",
18952 => "0000100001111100",
18953 => "0000100001111101",
18954 => "0000100001111101",
18955 => "0000100001111110",
18956 => "0000100001111110",
18957 => "0000100001111111",
18958 => "0000100001111111",
18959 => "0000100010000000",
18960 => "0000100010000000",
18961 => "0000100010000001",
18962 => "0000100010000001",
18963 => "0000100010000010",
18964 => "0000100010000010",
18965 => "0000100010000011",
18966 => "0000100010000011",
18967 => "0000100010000100",
18968 => "0000100010000100",
18969 => "0000100010000101",
18970 => "0000100010000101",
18971 => "0000100010000110",
18972 => "0000100010000110",
18973 => "0000100010000111",
18974 => "0000100010000111",
18975 => "0000100010001000",
18976 => "0000100010001000",
18977 => "0000100010001001",
18978 => "0000100010001001",
18979 => "0000100010001010",
18980 => "0000100010001010",
18981 => "0000100010001011",
18982 => "0000100010001100",
18983 => "0000100010001100",
18984 => "0000100010001101",
18985 => "0000100010001101",
18986 => "0000100010001110",
18987 => "0000100010001110",
18988 => "0000100010001111",
18989 => "0000100010001111",
18990 => "0000100010010000",
18991 => "0000100010010000",
18992 => "0000100010010001",
18993 => "0000100010010001",
18994 => "0000100010010010",
18995 => "0000100010010010",
18996 => "0000100010010011",
18997 => "0000100010010011",
18998 => "0000100010010100",
18999 => "0000100010010100",
19000 => "0000100010010101",
19001 => "0000100010010101",
19002 => "0000100010010110",
19003 => "0000100010010110",
19004 => "0000100010010111",
19005 => "0000100010010111",
19006 => "0000100010011000",
19007 => "0000100010011000",
19008 => "0000100010011001",
19009 => "0000100010011001",
19010 => "0000100010011010",
19011 => "0000100010011011",
19012 => "0000100010011011",
19013 => "0000100010011100",
19014 => "0000100010011100",
19015 => "0000100010011101",
19016 => "0000100010011101",
19017 => "0000100010011110",
19018 => "0000100010011110",
19019 => "0000100010011111",
19020 => "0000100010011111",
19021 => "0000100010100000",
19022 => "0000100010100000",
19023 => "0000100010100001",
19024 => "0000100010100001",
19025 => "0000100010100010",
19026 => "0000100010100010",
19027 => "0000100010100011",
19028 => "0000100010100011",
19029 => "0000100010100100",
19030 => "0000100010100100",
19031 => "0000100010100101",
19032 => "0000100010100101",
19033 => "0000100010100110",
19034 => "0000100010100111",
19035 => "0000100010100111",
19036 => "0000100010101000",
19037 => "0000100010101000",
19038 => "0000100010101001",
19039 => "0000100010101001",
19040 => "0000100010101010",
19041 => "0000100010101010",
19042 => "0000100010101011",
19043 => "0000100010101011",
19044 => "0000100010101100",
19045 => "0000100010101100",
19046 => "0000100010101101",
19047 => "0000100010101101",
19048 => "0000100010101110",
19049 => "0000100010101110",
19050 => "0000100010101111",
19051 => "0000100010101111",
19052 => "0000100010110000",
19053 => "0000100010110000",
19054 => "0000100010110001",
19055 => "0000100010110010",
19056 => "0000100010110010",
19057 => "0000100010110011",
19058 => "0000100010110011",
19059 => "0000100010110100",
19060 => "0000100010110100",
19061 => "0000100010110101",
19062 => "0000100010110101",
19063 => "0000100010110110",
19064 => "0000100010110110",
19065 => "0000100010110111",
19066 => "0000100010110111",
19067 => "0000100010111000",
19068 => "0000100010111000",
19069 => "0000100010111001",
19070 => "0000100010111001",
19071 => "0000100010111010",
19072 => "0000100010111010",
19073 => "0000100010111011",
19074 => "0000100010111100",
19075 => "0000100010111100",
19076 => "0000100010111101",
19077 => "0000100010111101",
19078 => "0000100010111110",
19079 => "0000100010111110",
19080 => "0000100010111111",
19081 => "0000100010111111",
19082 => "0000100011000000",
19083 => "0000100011000000",
19084 => "0000100011000001",
19085 => "0000100011000001",
19086 => "0000100011000010",
19087 => "0000100011000010",
19088 => "0000100011000011",
19089 => "0000100011000011",
19090 => "0000100011000100",
19091 => "0000100011000100",
19092 => "0000100011000101",
19093 => "0000100011000110",
19094 => "0000100011000110",
19095 => "0000100011000111",
19096 => "0000100011000111",
19097 => "0000100011001000",
19098 => "0000100011001000",
19099 => "0000100011001001",
19100 => "0000100011001001",
19101 => "0000100011001010",
19102 => "0000100011001010",
19103 => "0000100011001011",
19104 => "0000100011001011",
19105 => "0000100011001100",
19106 => "0000100011001100",
19107 => "0000100011001101",
19108 => "0000100011001110",
19109 => "0000100011001110",
19110 => "0000100011001111",
19111 => "0000100011001111",
19112 => "0000100011010000",
19113 => "0000100011010000",
19114 => "0000100011010001",
19115 => "0000100011010001",
19116 => "0000100011010010",
19117 => "0000100011010010",
19118 => "0000100011010011",
19119 => "0000100011010011",
19120 => "0000100011010100",
19121 => "0000100011010100",
19122 => "0000100011010101",
19123 => "0000100011010101",
19124 => "0000100011010110",
19125 => "0000100011010111",
19126 => "0000100011010111",
19127 => "0000100011011000",
19128 => "0000100011011000",
19129 => "0000100011011001",
19130 => "0000100011011001",
19131 => "0000100011011010",
19132 => "0000100011011010",
19133 => "0000100011011011",
19134 => "0000100011011011",
19135 => "0000100011011100",
19136 => "0000100011011100",
19137 => "0000100011011101",
19138 => "0000100011011110",
19139 => "0000100011011110",
19140 => "0000100011011111",
19141 => "0000100011011111",
19142 => "0000100011100000",
19143 => "0000100011100000",
19144 => "0000100011100001",
19145 => "0000100011100001",
19146 => "0000100011100010",
19147 => "0000100011100010",
19148 => "0000100011100011",
19149 => "0000100011100011",
19150 => "0000100011100100",
19151 => "0000100011100100",
19152 => "0000100011100101",
19153 => "0000100011100110",
19154 => "0000100011100110",
19155 => "0000100011100111",
19156 => "0000100011100111",
19157 => "0000100011101000",
19158 => "0000100011101000",
19159 => "0000100011101001",
19160 => "0000100011101001",
19161 => "0000100011101010",
19162 => "0000100011101010",
19163 => "0000100011101011",
19164 => "0000100011101011",
19165 => "0000100011101100",
19166 => "0000100011101101",
19167 => "0000100011101101",
19168 => "0000100011101110",
19169 => "0000100011101110",
19170 => "0000100011101111",
19171 => "0000100011101111",
19172 => "0000100011110000",
19173 => "0000100011110000",
19174 => "0000100011110001",
19175 => "0000100011110001",
19176 => "0000100011110010",
19177 => "0000100011110010",
19178 => "0000100011110011",
19179 => "0000100011110100",
19180 => "0000100011110100",
19181 => "0000100011110101",
19182 => "0000100011110101",
19183 => "0000100011110110",
19184 => "0000100011110110",
19185 => "0000100011110111",
19186 => "0000100011110111",
19187 => "0000100011111000",
19188 => "0000100011111000",
19189 => "0000100011111001",
19190 => "0000100011111001",
19191 => "0000100011111010",
19192 => "0000100011111011",
19193 => "0000100011111011",
19194 => "0000100011111100",
19195 => "0000100011111100",
19196 => "0000100011111101",
19197 => "0000100011111101",
19198 => "0000100011111110",
19199 => "0000100011111110",
19200 => "0000100011111111",
19201 => "0000100011111111",
19202 => "0000100100000000",
19203 => "0000100100000001",
19204 => "0000100100000001",
19205 => "0000100100000010",
19206 => "0000100100000010",
19207 => "0000100100000011",
19208 => "0000100100000011",
19209 => "0000100100000100",
19210 => "0000100100000100",
19211 => "0000100100000101",
19212 => "0000100100000101",
19213 => "0000100100000110",
19214 => "0000100100000111",
19215 => "0000100100000111",
19216 => "0000100100001000",
19217 => "0000100100001000",
19218 => "0000100100001001",
19219 => "0000100100001001",
19220 => "0000100100001010",
19221 => "0000100100001010",
19222 => "0000100100001011",
19223 => "0000100100001011",
19224 => "0000100100001100",
19225 => "0000100100001101",
19226 => "0000100100001101",
19227 => "0000100100001110",
19228 => "0000100100001110",
19229 => "0000100100001111",
19230 => "0000100100001111",
19231 => "0000100100010000",
19232 => "0000100100010000",
19233 => "0000100100010001",
19234 => "0000100100010001",
19235 => "0000100100010010",
19236 => "0000100100010011",
19237 => "0000100100010011",
19238 => "0000100100010100",
19239 => "0000100100010100",
19240 => "0000100100010101",
19241 => "0000100100010101",
19242 => "0000100100010110",
19243 => "0000100100010110",
19244 => "0000100100010111",
19245 => "0000100100010111",
19246 => "0000100100011000",
19247 => "0000100100011001",
19248 => "0000100100011001",
19249 => "0000100100011010",
19250 => "0000100100011010",
19251 => "0000100100011011",
19252 => "0000100100011011",
19253 => "0000100100011100",
19254 => "0000100100011100",
19255 => "0000100100011101",
19256 => "0000100100011101",
19257 => "0000100100011110",
19258 => "0000100100011111",
19259 => "0000100100011111",
19260 => "0000100100100000",
19261 => "0000100100100000",
19262 => "0000100100100001",
19263 => "0000100100100001",
19264 => "0000100100100010",
19265 => "0000100100100010",
19266 => "0000100100100011",
19267 => "0000100100100100",
19268 => "0000100100100100",
19269 => "0000100100100101",
19270 => "0000100100100101",
19271 => "0000100100100110",
19272 => "0000100100100110",
19273 => "0000100100100111",
19274 => "0000100100100111",
19275 => "0000100100101000",
19276 => "0000100100101001",
19277 => "0000100100101001",
19278 => "0000100100101010",
19279 => "0000100100101010",
19280 => "0000100100101011",
19281 => "0000100100101011",
19282 => "0000100100101100",
19283 => "0000100100101100",
19284 => "0000100100101101",
19285 => "0000100100101101",
19286 => "0000100100101110",
19287 => "0000100100101111",
19288 => "0000100100101111",
19289 => "0000100100110000",
19290 => "0000100100110000",
19291 => "0000100100110001",
19292 => "0000100100110001",
19293 => "0000100100110010",
19294 => "0000100100110010",
19295 => "0000100100110011",
19296 => "0000100100110100",
19297 => "0000100100110100",
19298 => "0000100100110101",
19299 => "0000100100110101",
19300 => "0000100100110110",
19301 => "0000100100110110",
19302 => "0000100100110111",
19303 => "0000100100110111",
19304 => "0000100100111000",
19305 => "0000100100111001",
19306 => "0000100100111001",
19307 => "0000100100111010",
19308 => "0000100100111010",
19309 => "0000100100111011",
19310 => "0000100100111011",
19311 => "0000100100111100",
19312 => "0000100100111100",
19313 => "0000100100111101",
19314 => "0000100100111110",
19315 => "0000100100111110",
19316 => "0000100100111111",
19317 => "0000100100111111",
19318 => "0000100101000000",
19319 => "0000100101000000",
19320 => "0000100101000001",
19321 => "0000100101000001",
19322 => "0000100101000010",
19323 => "0000100101000011",
19324 => "0000100101000011",
19325 => "0000100101000100",
19326 => "0000100101000100",
19327 => "0000100101000101",
19328 => "0000100101000101",
19329 => "0000100101000110",
19330 => "0000100101000110",
19331 => "0000100101000111",
19332 => "0000100101001000",
19333 => "0000100101001000",
19334 => "0000100101001001",
19335 => "0000100101001001",
19336 => "0000100101001010",
19337 => "0000100101001010",
19338 => "0000100101001011",
19339 => "0000100101001100",
19340 => "0000100101001100",
19341 => "0000100101001101",
19342 => "0000100101001101",
19343 => "0000100101001110",
19344 => "0000100101001110",
19345 => "0000100101001111",
19346 => "0000100101001111",
19347 => "0000100101010000",
19348 => "0000100101010001",
19349 => "0000100101010001",
19350 => "0000100101010010",
19351 => "0000100101010010",
19352 => "0000100101010011",
19353 => "0000100101010011",
19354 => "0000100101010100",
19355 => "0000100101010101",
19356 => "0000100101010101",
19357 => "0000100101010110",
19358 => "0000100101010110",
19359 => "0000100101010111",
19360 => "0000100101010111",
19361 => "0000100101011000",
19362 => "0000100101011000",
19363 => "0000100101011001",
19364 => "0000100101011010",
19365 => "0000100101011010",
19366 => "0000100101011011",
19367 => "0000100101011011",
19368 => "0000100101011100",
19369 => "0000100101011100",
19370 => "0000100101011101",
19371 => "0000100101011110",
19372 => "0000100101011110",
19373 => "0000100101011111",
19374 => "0000100101011111",
19375 => "0000100101100000",
19376 => "0000100101100000",
19377 => "0000100101100001",
19378 => "0000100101100001",
19379 => "0000100101100010",
19380 => "0000100101100011",
19381 => "0000100101100011",
19382 => "0000100101100100",
19383 => "0000100101100100",
19384 => "0000100101100101",
19385 => "0000100101100101",
19386 => "0000100101100110",
19387 => "0000100101100111",
19388 => "0000100101100111",
19389 => "0000100101101000",
19390 => "0000100101101000",
19391 => "0000100101101001",
19392 => "0000100101101001",
19393 => "0000100101101010",
19394 => "0000100101101011",
19395 => "0000100101101011",
19396 => "0000100101101100",
19397 => "0000100101101100",
19398 => "0000100101101101",
19399 => "0000100101101101",
19400 => "0000100101101110",
19401 => "0000100101101110",
19402 => "0000100101101111",
19403 => "0000100101110000",
19404 => "0000100101110000",
19405 => "0000100101110001",
19406 => "0000100101110001",
19407 => "0000100101110010",
19408 => "0000100101110010",
19409 => "0000100101110011",
19410 => "0000100101110100",
19411 => "0000100101110100",
19412 => "0000100101110101",
19413 => "0000100101110101",
19414 => "0000100101110110",
19415 => "0000100101110110",
19416 => "0000100101110111",
19417 => "0000100101111000",
19418 => "0000100101111000",
19419 => "0000100101111001",
19420 => "0000100101111001",
19421 => "0000100101111010",
19422 => "0000100101111010",
19423 => "0000100101111011",
19424 => "0000100101111100",
19425 => "0000100101111100",
19426 => "0000100101111101",
19427 => "0000100101111101",
19428 => "0000100101111110",
19429 => "0000100101111110",
19430 => "0000100101111111",
19431 => "0000100110000000",
19432 => "0000100110000000",
19433 => "0000100110000001",
19434 => "0000100110000001",
19435 => "0000100110000010",
19436 => "0000100110000010",
19437 => "0000100110000011",
19438 => "0000100110000100",
19439 => "0000100110000100",
19440 => "0000100110000101",
19441 => "0000100110000101",
19442 => "0000100110000110",
19443 => "0000100110000110",
19444 => "0000100110000111",
19445 => "0000100110001000",
19446 => "0000100110001000",
19447 => "0000100110001001",
19448 => "0000100110001001",
19449 => "0000100110001010",
19450 => "0000100110001010",
19451 => "0000100110001011",
19452 => "0000100110001100",
19453 => "0000100110001100",
19454 => "0000100110001101",
19455 => "0000100110001101",
19456 => "0000100110001110",
19457 => "0000100110001111",
19458 => "0000100110001111",
19459 => "0000100110010000",
19460 => "0000100110010000",
19461 => "0000100110010001",
19462 => "0000100110010001",
19463 => "0000100110010010",
19464 => "0000100110010011",
19465 => "0000100110010011",
19466 => "0000100110010100",
19467 => "0000100110010100",
19468 => "0000100110010101",
19469 => "0000100110010101",
19470 => "0000100110010110",
19471 => "0000100110010111",
19472 => "0000100110010111",
19473 => "0000100110011000",
19474 => "0000100110011000",
19475 => "0000100110011001",
19476 => "0000100110011001",
19477 => "0000100110011010",
19478 => "0000100110011011",
19479 => "0000100110011011",
19480 => "0000100110011100",
19481 => "0000100110011100",
19482 => "0000100110011101",
19483 => "0000100110011101",
19484 => "0000100110011110",
19485 => "0000100110011111",
19486 => "0000100110011111",
19487 => "0000100110100000",
19488 => "0000100110100000",
19489 => "0000100110100001",
19490 => "0000100110100010",
19491 => "0000100110100010",
19492 => "0000100110100011",
19493 => "0000100110100011",
19494 => "0000100110100100",
19495 => "0000100110100100",
19496 => "0000100110100101",
19497 => "0000100110100110",
19498 => "0000100110100110",
19499 => "0000100110100111",
19500 => "0000100110100111",
19501 => "0000100110101000",
19502 => "0000100110101001",
19503 => "0000100110101001",
19504 => "0000100110101010",
19505 => "0000100110101010",
19506 => "0000100110101011",
19507 => "0000100110101011",
19508 => "0000100110101100",
19509 => "0000100110101101",
19510 => "0000100110101101",
19511 => "0000100110101110",
19512 => "0000100110101110",
19513 => "0000100110101111",
19514 => "0000100110101111",
19515 => "0000100110110000",
19516 => "0000100110110001",
19517 => "0000100110110001",
19518 => "0000100110110010",
19519 => "0000100110110010",
19520 => "0000100110110011",
19521 => "0000100110110100",
19522 => "0000100110110100",
19523 => "0000100110110101",
19524 => "0000100110110101",
19525 => "0000100110110110",
19526 => "0000100110110110",
19527 => "0000100110110111",
19528 => "0000100110111000",
19529 => "0000100110111000",
19530 => "0000100110111001",
19531 => "0000100110111001",
19532 => "0000100110111010",
19533 => "0000100110111011",
19534 => "0000100110111011",
19535 => "0000100110111100",
19536 => "0000100110111100",
19537 => "0000100110111101",
19538 => "0000100110111110",
19539 => "0000100110111110",
19540 => "0000100110111111",
19541 => "0000100110111111",
19542 => "0000100111000000",
19543 => "0000100111000000",
19544 => "0000100111000001",
19545 => "0000100111000010",
19546 => "0000100111000010",
19547 => "0000100111000011",
19548 => "0000100111000011",
19549 => "0000100111000100",
19550 => "0000100111000101",
19551 => "0000100111000101",
19552 => "0000100111000110",
19553 => "0000100111000110",
19554 => "0000100111000111",
19555 => "0000100111000111",
19556 => "0000100111001000",
19557 => "0000100111001001",
19558 => "0000100111001001",
19559 => "0000100111001010",
19560 => "0000100111001010",
19561 => "0000100111001011",
19562 => "0000100111001100",
19563 => "0000100111001100",
19564 => "0000100111001101",
19565 => "0000100111001101",
19566 => "0000100111001110",
19567 => "0000100111001111",
19568 => "0000100111001111",
19569 => "0000100111010000",
19570 => "0000100111010000",
19571 => "0000100111010001",
19572 => "0000100111010010",
19573 => "0000100111010010",
19574 => "0000100111010011",
19575 => "0000100111010011",
19576 => "0000100111010100",
19577 => "0000100111010100",
19578 => "0000100111010101",
19579 => "0000100111010110",
19580 => "0000100111010110",
19581 => "0000100111010111",
19582 => "0000100111010111",
19583 => "0000100111011000",
19584 => "0000100111011001",
19585 => "0000100111011001",
19586 => "0000100111011010",
19587 => "0000100111011010",
19588 => "0000100111011011",
19589 => "0000100111011100",
19590 => "0000100111011100",
19591 => "0000100111011101",
19592 => "0000100111011101",
19593 => "0000100111011110",
19594 => "0000100111011111",
19595 => "0000100111011111",
19596 => "0000100111100000",
19597 => "0000100111100000",
19598 => "0000100111100001",
19599 => "0000100111100001",
19600 => "0000100111100010",
19601 => "0000100111100011",
19602 => "0000100111100011",
19603 => "0000100111100100",
19604 => "0000100111100100",
19605 => "0000100111100101",
19606 => "0000100111100110",
19607 => "0000100111100110",
19608 => "0000100111100111",
19609 => "0000100111100111",
19610 => "0000100111101000",
19611 => "0000100111101001",
19612 => "0000100111101001",
19613 => "0000100111101010",
19614 => "0000100111101010",
19615 => "0000100111101011",
19616 => "0000100111101100",
19617 => "0000100111101100",
19618 => "0000100111101101",
19619 => "0000100111101101",
19620 => "0000100111101110",
19621 => "0000100111101111",
19622 => "0000100111101111",
19623 => "0000100111110000",
19624 => "0000100111110000",
19625 => "0000100111110001",
19626 => "0000100111110010",
19627 => "0000100111110010",
19628 => "0000100111110011",
19629 => "0000100111110011",
19630 => "0000100111110100",
19631 => "0000100111110101",
19632 => "0000100111110101",
19633 => "0000100111110110",
19634 => "0000100111110110",
19635 => "0000100111110111",
19636 => "0000100111111000",
19637 => "0000100111111000",
19638 => "0000100111111001",
19639 => "0000100111111001",
19640 => "0000100111111010",
19641 => "0000100111111011",
19642 => "0000100111111011",
19643 => "0000100111111100",
19644 => "0000100111111100",
19645 => "0000100111111101",
19646 => "0000100111111110",
19647 => "0000100111111110",
19648 => "0000100111111111",
19649 => "0000100111111111",
19650 => "0000101000000000",
19651 => "0000101000000001",
19652 => "0000101000000001",
19653 => "0000101000000010",
19654 => "0000101000000010",
19655 => "0000101000000011",
19656 => "0000101000000100",
19657 => "0000101000000100",
19658 => "0000101000000101",
19659 => "0000101000000101",
19660 => "0000101000000110",
19661 => "0000101000000111",
19662 => "0000101000000111",
19663 => "0000101000001000",
19664 => "0000101000001000",
19665 => "0000101000001001",
19666 => "0000101000001010",
19667 => "0000101000001010",
19668 => "0000101000001011",
19669 => "0000101000001011",
19670 => "0000101000001100",
19671 => "0000101000001101",
19672 => "0000101000001101",
19673 => "0000101000001110",
19674 => "0000101000001110",
19675 => "0000101000001111",
19676 => "0000101000010000",
19677 => "0000101000010000",
19678 => "0000101000010001",
19679 => "0000101000010001",
19680 => "0000101000010010",
19681 => "0000101000010011",
19682 => "0000101000010011",
19683 => "0000101000010100",
19684 => "0000101000010100",
19685 => "0000101000010101",
19686 => "0000101000010110",
19687 => "0000101000010110",
19688 => "0000101000010111",
19689 => "0000101000010111",
19690 => "0000101000011000",
19691 => "0000101000011001",
19692 => "0000101000011001",
19693 => "0000101000011010",
19694 => "0000101000011011",
19695 => "0000101000011011",
19696 => "0000101000011100",
19697 => "0000101000011100",
19698 => "0000101000011101",
19699 => "0000101000011110",
19700 => "0000101000011110",
19701 => "0000101000011111",
19702 => "0000101000011111",
19703 => "0000101000100000",
19704 => "0000101000100001",
19705 => "0000101000100001",
19706 => "0000101000100010",
19707 => "0000101000100010",
19708 => "0000101000100011",
19709 => "0000101000100100",
19710 => "0000101000100100",
19711 => "0000101000100101",
19712 => "0000101000100101",
19713 => "0000101000100110",
19714 => "0000101000100111",
19715 => "0000101000100111",
19716 => "0000101000101000",
19717 => "0000101000101001",
19718 => "0000101000101001",
19719 => "0000101000101010",
19720 => "0000101000101010",
19721 => "0000101000101011",
19722 => "0000101000101100",
19723 => "0000101000101100",
19724 => "0000101000101101",
19725 => "0000101000101101",
19726 => "0000101000101110",
19727 => "0000101000101111",
19728 => "0000101000101111",
19729 => "0000101000110000",
19730 => "0000101000110000",
19731 => "0000101000110001",
19732 => "0000101000110010",
19733 => "0000101000110010",
19734 => "0000101000110011",
19735 => "0000101000110100",
19736 => "0000101000110100",
19737 => "0000101000110101",
19738 => "0000101000110101",
19739 => "0000101000110110",
19740 => "0000101000110111",
19741 => "0000101000110111",
19742 => "0000101000111000",
19743 => "0000101000111000",
19744 => "0000101000111001",
19745 => "0000101000111010",
19746 => "0000101000111010",
19747 => "0000101000111011",
19748 => "0000101000111011",
19749 => "0000101000111100",
19750 => "0000101000111101",
19751 => "0000101000111101",
19752 => "0000101000111110",
19753 => "0000101000111111",
19754 => "0000101000111111",
19755 => "0000101001000000",
19756 => "0000101001000000",
19757 => "0000101001000001",
19758 => "0000101001000010",
19759 => "0000101001000010",
19760 => "0000101001000011",
19761 => "0000101001000011",
19762 => "0000101001000100",
19763 => "0000101001000101",
19764 => "0000101001000101",
19765 => "0000101001000110",
19766 => "0000101001000111",
19767 => "0000101001000111",
19768 => "0000101001001000",
19769 => "0000101001001000",
19770 => "0000101001001001",
19771 => "0000101001001010",
19772 => "0000101001001010",
19773 => "0000101001001011",
19774 => "0000101001001011",
19775 => "0000101001001100",
19776 => "0000101001001101",
19777 => "0000101001001101",
19778 => "0000101001001110",
19779 => "0000101001001111",
19780 => "0000101001001111",
19781 => "0000101001010000",
19782 => "0000101001010000",
19783 => "0000101001010001",
19784 => "0000101001010010",
19785 => "0000101001010010",
19786 => "0000101001010011",
19787 => "0000101001010100",
19788 => "0000101001010100",
19789 => "0000101001010101",
19790 => "0000101001010101",
19791 => "0000101001010110",
19792 => "0000101001010111",
19793 => "0000101001010111",
19794 => "0000101001011000",
19795 => "0000101001011000",
19796 => "0000101001011001",
19797 => "0000101001011010",
19798 => "0000101001011010",
19799 => "0000101001011011",
19800 => "0000101001011100",
19801 => "0000101001011100",
19802 => "0000101001011101",
19803 => "0000101001011101",
19804 => "0000101001011110",
19805 => "0000101001011111",
19806 => "0000101001011111",
19807 => "0000101001100000",
19808 => "0000101001100001",
19809 => "0000101001100001",
19810 => "0000101001100010",
19811 => "0000101001100010",
19812 => "0000101001100011",
19813 => "0000101001100100",
19814 => "0000101001100100",
19815 => "0000101001100101",
19816 => "0000101001100110",
19817 => "0000101001100110",
19818 => "0000101001100111",
19819 => "0000101001100111",
19820 => "0000101001101000",
19821 => "0000101001101001",
19822 => "0000101001101001",
19823 => "0000101001101010",
19824 => "0000101001101011",
19825 => "0000101001101011",
19826 => "0000101001101100",
19827 => "0000101001101100",
19828 => "0000101001101101",
19829 => "0000101001101110",
19830 => "0000101001101110",
19831 => "0000101001101111",
19832 => "0000101001110000",
19833 => "0000101001110000",
19834 => "0000101001110001",
19835 => "0000101001110001",
19836 => "0000101001110010",
19837 => "0000101001110011",
19838 => "0000101001110011",
19839 => "0000101001110100",
19840 => "0000101001110101",
19841 => "0000101001110101",
19842 => "0000101001110110",
19843 => "0000101001110110",
19844 => "0000101001110111",
19845 => "0000101001111000",
19846 => "0000101001111000",
19847 => "0000101001111001",
19848 => "0000101001111010",
19849 => "0000101001111010",
19850 => "0000101001111011",
19851 => "0000101001111011",
19852 => "0000101001111100",
19853 => "0000101001111101",
19854 => "0000101001111101",
19855 => "0000101001111110",
19856 => "0000101001111111",
19857 => "0000101001111111",
19858 => "0000101010000000",
19859 => "0000101010000000",
19860 => "0000101010000001",
19861 => "0000101010000010",
19862 => "0000101010000010",
19863 => "0000101010000011",
19864 => "0000101010000100",
19865 => "0000101010000100",
19866 => "0000101010000101",
19867 => "0000101010000110",
19868 => "0000101010000110",
19869 => "0000101010000111",
19870 => "0000101010000111",
19871 => "0000101010001000",
19872 => "0000101010001001",
19873 => "0000101010001001",
19874 => "0000101010001010",
19875 => "0000101010001011",
19876 => "0000101010001011",
19877 => "0000101010001100",
19878 => "0000101010001100",
19879 => "0000101010001101",
19880 => "0000101010001110",
19881 => "0000101010001110",
19882 => "0000101010001111",
19883 => "0000101010010000",
19884 => "0000101010010000",
19885 => "0000101010010001",
19886 => "0000101010010010",
19887 => "0000101010010010",
19888 => "0000101010010011",
19889 => "0000101010010011",
19890 => "0000101010010100",
19891 => "0000101010010101",
19892 => "0000101010010101",
19893 => "0000101010010110",
19894 => "0000101010010111",
19895 => "0000101010010111",
19896 => "0000101010011000",
19897 => "0000101010011001",
19898 => "0000101010011001",
19899 => "0000101010011010",
19900 => "0000101010011010",
19901 => "0000101010011011",
19902 => "0000101010011100",
19903 => "0000101010011100",
19904 => "0000101010011101",
19905 => "0000101010011110",
19906 => "0000101010011110",
19907 => "0000101010011111",
19908 => "0000101010100000",
19909 => "0000101010100000",
19910 => "0000101010100001",
19911 => "0000101010100001",
19912 => "0000101010100010",
19913 => "0000101010100011",
19914 => "0000101010100011",
19915 => "0000101010100100",
19916 => "0000101010100101",
19917 => "0000101010100101",
19918 => "0000101010100110",
19919 => "0000101010100111",
19920 => "0000101010100111",
19921 => "0000101010101000",
19922 => "0000101010101000",
19923 => "0000101010101001",
19924 => "0000101010101010",
19925 => "0000101010101010",
19926 => "0000101010101011",
19927 => "0000101010101100",
19928 => "0000101010101100",
19929 => "0000101010101101",
19930 => "0000101010101110",
19931 => "0000101010101110",
19932 => "0000101010101111",
19933 => "0000101010101111",
19934 => "0000101010110000",
19935 => "0000101010110001",
19936 => "0000101010110001",
19937 => "0000101010110010",
19938 => "0000101010110011",
19939 => "0000101010110011",
19940 => "0000101010110100",
19941 => "0000101010110101",
19942 => "0000101010110101",
19943 => "0000101010110110",
19944 => "0000101010110111",
19945 => "0000101010110111",
19946 => "0000101010111000",
19947 => "0000101010111000",
19948 => "0000101010111001",
19949 => "0000101010111010",
19950 => "0000101010111010",
19951 => "0000101010111011",
19952 => "0000101010111100",
19953 => "0000101010111100",
19954 => "0000101010111101",
19955 => "0000101010111110",
19956 => "0000101010111110",
19957 => "0000101010111111",
19958 => "0000101011000000",
19959 => "0000101011000000",
19960 => "0000101011000001",
19961 => "0000101011000001",
19962 => "0000101011000010",
19963 => "0000101011000011",
19964 => "0000101011000011",
19965 => "0000101011000100",
19966 => "0000101011000101",
19967 => "0000101011000101",
19968 => "0000101011000110",
19969 => "0000101011000111",
19970 => "0000101011000111",
19971 => "0000101011001000",
19972 => "0000101011001001",
19973 => "0000101011001001",
19974 => "0000101011001010",
19975 => "0000101011001010",
19976 => "0000101011001011",
19977 => "0000101011001100",
19978 => "0000101011001100",
19979 => "0000101011001101",
19980 => "0000101011001110",
19981 => "0000101011001110",
19982 => "0000101011001111",
19983 => "0000101011010000",
19984 => "0000101011010000",
19985 => "0000101011010001",
19986 => "0000101011010010",
19987 => "0000101011010010",
19988 => "0000101011010011",
19989 => "0000101011010100",
19990 => "0000101011010100",
19991 => "0000101011010101",
19992 => "0000101011010101",
19993 => "0000101011010110",
19994 => "0000101011010111",
19995 => "0000101011010111",
19996 => "0000101011011000",
19997 => "0000101011011001",
19998 => "0000101011011001",
19999 => "0000101011011010",
20000 => "0000101011011011",
20001 => "0000101011011011",
20002 => "0000101011011100",
20003 => "0000101011011101",
20004 => "0000101011011101",
20005 => "0000101011011110",
20006 => "0000101011011111",
20007 => "0000101011011111",
20008 => "0000101011100000",
20009 => "0000101011100001",
20010 => "0000101011100001",
20011 => "0000101011100010",
20012 => "0000101011100010",
20013 => "0000101011100011",
20014 => "0000101011100100",
20015 => "0000101011100100",
20016 => "0000101011100101",
20017 => "0000101011100110",
20018 => "0000101011100110",
20019 => "0000101011100111",
20020 => "0000101011101000",
20021 => "0000101011101000",
20022 => "0000101011101001",
20023 => "0000101011101010",
20024 => "0000101011101010",
20025 => "0000101011101011",
20026 => "0000101011101100",
20027 => "0000101011101100",
20028 => "0000101011101101",
20029 => "0000101011101110",
20030 => "0000101011101110",
20031 => "0000101011101111",
20032 => "0000101011110000",
20033 => "0000101011110000",
20034 => "0000101011110001",
20035 => "0000101011110010",
20036 => "0000101011110010",
20037 => "0000101011110011",
20038 => "0000101011110011",
20039 => "0000101011110100",
20040 => "0000101011110101",
20041 => "0000101011110101",
20042 => "0000101011110110",
20043 => "0000101011110111",
20044 => "0000101011110111",
20045 => "0000101011111000",
20046 => "0000101011111001",
20047 => "0000101011111001",
20048 => "0000101011111010",
20049 => "0000101011111011",
20050 => "0000101011111011",
20051 => "0000101011111100",
20052 => "0000101011111101",
20053 => "0000101011111101",
20054 => "0000101011111110",
20055 => "0000101011111111",
20056 => "0000101011111111",
20057 => "0000101100000000",
20058 => "0000101100000001",
20059 => "0000101100000001",
20060 => "0000101100000010",
20061 => "0000101100000011",
20062 => "0000101100000011",
20063 => "0000101100000100",
20064 => "0000101100000101",
20065 => "0000101100000101",
20066 => "0000101100000110",
20067 => "0000101100000111",
20068 => "0000101100000111",
20069 => "0000101100001000",
20070 => "0000101100001001",
20071 => "0000101100001001",
20072 => "0000101100001010",
20073 => "0000101100001010",
20074 => "0000101100001011",
20075 => "0000101100001100",
20076 => "0000101100001100",
20077 => "0000101100001101",
20078 => "0000101100001110",
20079 => "0000101100001110",
20080 => "0000101100001111",
20081 => "0000101100010000",
20082 => "0000101100010000",
20083 => "0000101100010001",
20084 => "0000101100010010",
20085 => "0000101100010010",
20086 => "0000101100010011",
20087 => "0000101100010100",
20088 => "0000101100010100",
20089 => "0000101100010101",
20090 => "0000101100010110",
20091 => "0000101100010110",
20092 => "0000101100010111",
20093 => "0000101100011000",
20094 => "0000101100011000",
20095 => "0000101100011001",
20096 => "0000101100011010",
20097 => "0000101100011010",
20098 => "0000101100011011",
20099 => "0000101100011100",
20100 => "0000101100011100",
20101 => "0000101100011101",
20102 => "0000101100011110",
20103 => "0000101100011110",
20104 => "0000101100011111",
20105 => "0000101100100000",
20106 => "0000101100100000",
20107 => "0000101100100001",
20108 => "0000101100100010",
20109 => "0000101100100010",
20110 => "0000101100100011",
20111 => "0000101100100100",
20112 => "0000101100100100",
20113 => "0000101100100101",
20114 => "0000101100100110",
20115 => "0000101100100110",
20116 => "0000101100100111",
20117 => "0000101100101000",
20118 => "0000101100101000",
20119 => "0000101100101001",
20120 => "0000101100101010",
20121 => "0000101100101010",
20122 => "0000101100101011",
20123 => "0000101100101100",
20124 => "0000101100101100",
20125 => "0000101100101101",
20126 => "0000101100101110",
20127 => "0000101100101110",
20128 => "0000101100101111",
20129 => "0000101100110000",
20130 => "0000101100110000",
20131 => "0000101100110001",
20132 => "0000101100110010",
20133 => "0000101100110010",
20134 => "0000101100110011",
20135 => "0000101100110100",
20136 => "0000101100110100",
20137 => "0000101100110101",
20138 => "0000101100110110",
20139 => "0000101100110110",
20140 => "0000101100110111",
20141 => "0000101100111000",
20142 => "0000101100111000",
20143 => "0000101100111001",
20144 => "0000101100111010",
20145 => "0000101100111010",
20146 => "0000101100111011",
20147 => "0000101100111100",
20148 => "0000101100111100",
20149 => "0000101100111101",
20150 => "0000101100111110",
20151 => "0000101100111110",
20152 => "0000101100111111",
20153 => "0000101101000000",
20154 => "0000101101000000",
20155 => "0000101101000001",
20156 => "0000101101000010",
20157 => "0000101101000010",
20158 => "0000101101000011",
20159 => "0000101101000100",
20160 => "0000101101000101",
20161 => "0000101101000101",
20162 => "0000101101000110",
20163 => "0000101101000111",
20164 => "0000101101000111",
20165 => "0000101101001000",
20166 => "0000101101001001",
20167 => "0000101101001001",
20168 => "0000101101001010",
20169 => "0000101101001011",
20170 => "0000101101001011",
20171 => "0000101101001100",
20172 => "0000101101001101",
20173 => "0000101101001101",
20174 => "0000101101001110",
20175 => "0000101101001111",
20176 => "0000101101001111",
20177 => "0000101101010000",
20178 => "0000101101010001",
20179 => "0000101101010001",
20180 => "0000101101010010",
20181 => "0000101101010011",
20182 => "0000101101010011",
20183 => "0000101101010100",
20184 => "0000101101010101",
20185 => "0000101101010101",
20186 => "0000101101010110",
20187 => "0000101101010111",
20188 => "0000101101010111",
20189 => "0000101101011000",
20190 => "0000101101011001",
20191 => "0000101101011001",
20192 => "0000101101011010",
20193 => "0000101101011011",
20194 => "0000101101011011",
20195 => "0000101101011100",
20196 => "0000101101011101",
20197 => "0000101101011110",
20198 => "0000101101011110",
20199 => "0000101101011111",
20200 => "0000101101100000",
20201 => "0000101101100000",
20202 => "0000101101100001",
20203 => "0000101101100010",
20204 => "0000101101100010",
20205 => "0000101101100011",
20206 => "0000101101100100",
20207 => "0000101101100100",
20208 => "0000101101100101",
20209 => "0000101101100110",
20210 => "0000101101100110",
20211 => "0000101101100111",
20212 => "0000101101101000",
20213 => "0000101101101000",
20214 => "0000101101101001",
20215 => "0000101101101010",
20216 => "0000101101101010",
20217 => "0000101101101011",
20218 => "0000101101101100",
20219 => "0000101101101101",
20220 => "0000101101101101",
20221 => "0000101101101110",
20222 => "0000101101101111",
20223 => "0000101101101111",
20224 => "0000101101110000",
20225 => "0000101101110001",
20226 => "0000101101110001",
20227 => "0000101101110010",
20228 => "0000101101110011",
20229 => "0000101101110011",
20230 => "0000101101110100",
20231 => "0000101101110101",
20232 => "0000101101110101",
20233 => "0000101101110110",
20234 => "0000101101110111",
20235 => "0000101101110111",
20236 => "0000101101111000",
20237 => "0000101101111001",
20238 => "0000101101111001",
20239 => "0000101101111010",
20240 => "0000101101111011",
20241 => "0000101101111100",
20242 => "0000101101111100",
20243 => "0000101101111101",
20244 => "0000101101111110",
20245 => "0000101101111110",
20246 => "0000101101111111",
20247 => "0000101110000000",
20248 => "0000101110000000",
20249 => "0000101110000001",
20250 => "0000101110000010",
20251 => "0000101110000010",
20252 => "0000101110000011",
20253 => "0000101110000100",
20254 => "0000101110000100",
20255 => "0000101110000101",
20256 => "0000101110000110",
20257 => "0000101110000111",
20258 => "0000101110000111",
20259 => "0000101110001000",
20260 => "0000101110001001",
20261 => "0000101110001001",
20262 => "0000101110001010",
20263 => "0000101110001011",
20264 => "0000101110001011",
20265 => "0000101110001100",
20266 => "0000101110001101",
20267 => "0000101110001101",
20268 => "0000101110001110",
20269 => "0000101110001111",
20270 => "0000101110001111",
20271 => "0000101110010000",
20272 => "0000101110010001",
20273 => "0000101110010010",
20274 => "0000101110010010",
20275 => "0000101110010011",
20276 => "0000101110010100",
20277 => "0000101110010100",
20278 => "0000101110010101",
20279 => "0000101110010110",
20280 => "0000101110010110",
20281 => "0000101110010111",
20282 => "0000101110011000",
20283 => "0000101110011000",
20284 => "0000101110011001",
20285 => "0000101110011010",
20286 => "0000101110011011",
20287 => "0000101110011011",
20288 => "0000101110011100",
20289 => "0000101110011101",
20290 => "0000101110011101",
20291 => "0000101110011110",
20292 => "0000101110011111",
20293 => "0000101110011111",
20294 => "0000101110100000",
20295 => "0000101110100001",
20296 => "0000101110100001",
20297 => "0000101110100010",
20298 => "0000101110100011",
20299 => "0000101110100100",
20300 => "0000101110100100",
20301 => "0000101110100101",
20302 => "0000101110100110",
20303 => "0000101110100110",
20304 => "0000101110100111",
20305 => "0000101110101000",
20306 => "0000101110101000",
20307 => "0000101110101001",
20308 => "0000101110101010",
20309 => "0000101110101011",
20310 => "0000101110101011",
20311 => "0000101110101100",
20312 => "0000101110101101",
20313 => "0000101110101101",
20314 => "0000101110101110",
20315 => "0000101110101111",
20316 => "0000101110101111",
20317 => "0000101110110000",
20318 => "0000101110110001",
20319 => "0000101110110001",
20320 => "0000101110110010",
20321 => "0000101110110011",
20322 => "0000101110110100",
20323 => "0000101110110100",
20324 => "0000101110110101",
20325 => "0000101110110110",
20326 => "0000101110110110",
20327 => "0000101110110111",
20328 => "0000101110111000",
20329 => "0000101110111000",
20330 => "0000101110111001",
20331 => "0000101110111010",
20332 => "0000101110111011",
20333 => "0000101110111011",
20334 => "0000101110111100",
20335 => "0000101110111101",
20336 => "0000101110111101",
20337 => "0000101110111110",
20338 => "0000101110111111",
20339 => "0000101110111111",
20340 => "0000101111000000",
20341 => "0000101111000001",
20342 => "0000101111000010",
20343 => "0000101111000010",
20344 => "0000101111000011",
20345 => "0000101111000100",
20346 => "0000101111000100",
20347 => "0000101111000101",
20348 => "0000101111000110",
20349 => "0000101111000110",
20350 => "0000101111000111",
20351 => "0000101111001000",
20352 => "0000101111001001",
20353 => "0000101111001001",
20354 => "0000101111001010",
20355 => "0000101111001011",
20356 => "0000101111001011",
20357 => "0000101111001100",
20358 => "0000101111001101",
20359 => "0000101111001110",
20360 => "0000101111001110",
20361 => "0000101111001111",
20362 => "0000101111010000",
20363 => "0000101111010000",
20364 => "0000101111010001",
20365 => "0000101111010010",
20366 => "0000101111010010",
20367 => "0000101111010011",
20368 => "0000101111010100",
20369 => "0000101111010101",
20370 => "0000101111010101",
20371 => "0000101111010110",
20372 => "0000101111010111",
20373 => "0000101111010111",
20374 => "0000101111011000",
20375 => "0000101111011001",
20376 => "0000101111011010",
20377 => "0000101111011010",
20378 => "0000101111011011",
20379 => "0000101111011100",
20380 => "0000101111011100",
20381 => "0000101111011101",
20382 => "0000101111011110",
20383 => "0000101111011110",
20384 => "0000101111011111",
20385 => "0000101111100000",
20386 => "0000101111100001",
20387 => "0000101111100001",
20388 => "0000101111100010",
20389 => "0000101111100011",
20390 => "0000101111100011",
20391 => "0000101111100100",
20392 => "0000101111100101",
20393 => "0000101111100110",
20394 => "0000101111100110",
20395 => "0000101111100111",
20396 => "0000101111101000",
20397 => "0000101111101000",
20398 => "0000101111101001",
20399 => "0000101111101010",
20400 => "0000101111101011",
20401 => "0000101111101011",
20402 => "0000101111101100",
20403 => "0000101111101101",
20404 => "0000101111101101",
20405 => "0000101111101110",
20406 => "0000101111101111",
20407 => "0000101111101111",
20408 => "0000101111110000",
20409 => "0000101111110001",
20410 => "0000101111110010",
20411 => "0000101111110010",
20412 => "0000101111110011",
20413 => "0000101111110100",
20414 => "0000101111110100",
20415 => "0000101111110101",
20416 => "0000101111110110",
20417 => "0000101111110111",
20418 => "0000101111110111",
20419 => "0000101111111000",
20420 => "0000101111111001",
20421 => "0000101111111001",
20422 => "0000101111111010",
20423 => "0000101111111011",
20424 => "0000101111111100",
20425 => "0000101111111100",
20426 => "0000101111111101",
20427 => "0000101111111110",
20428 => "0000101111111110",
20429 => "0000101111111111",
20430 => "0000110000000000",
20431 => "0000110000000001",
20432 => "0000110000000001",
20433 => "0000110000000010",
20434 => "0000110000000011",
20435 => "0000110000000011",
20436 => "0000110000000100",
20437 => "0000110000000101",
20438 => "0000110000000110",
20439 => "0000110000000110",
20440 => "0000110000000111",
20441 => "0000110000001000",
20442 => "0000110000001000",
20443 => "0000110000001001",
20444 => "0000110000001010",
20445 => "0000110000001011",
20446 => "0000110000001011",
20447 => "0000110000001100",
20448 => "0000110000001101",
20449 => "0000110000001101",
20450 => "0000110000001110",
20451 => "0000110000001111",
20452 => "0000110000010000",
20453 => "0000110000010000",
20454 => "0000110000010001",
20455 => "0000110000010010",
20456 => "0000110000010011",
20457 => "0000110000010011",
20458 => "0000110000010100",
20459 => "0000110000010101",
20460 => "0000110000010101",
20461 => "0000110000010110",
20462 => "0000110000010111",
20463 => "0000110000011000",
20464 => "0000110000011000",
20465 => "0000110000011001",
20466 => "0000110000011010",
20467 => "0000110000011010",
20468 => "0000110000011011",
20469 => "0000110000011100",
20470 => "0000110000011101",
20471 => "0000110000011101",
20472 => "0000110000011110",
20473 => "0000110000011111",
20474 => "0000110000011111",
20475 => "0000110000100000",
20476 => "0000110000100001",
20477 => "0000110000100010",
20478 => "0000110000100010",
20479 => "0000110000100011",
20480 => "0000110000100100",
20481 => "0000110000100101",
20482 => "0000110000100101",
20483 => "0000110000100110",
20484 => "0000110000100111",
20485 => "0000110000100111",
20486 => "0000110000101000",
20487 => "0000110000101001",
20488 => "0000110000101010",
20489 => "0000110000101010",
20490 => "0000110000101011",
20491 => "0000110000101100",
20492 => "0000110000101101",
20493 => "0000110000101101",
20494 => "0000110000101110",
20495 => "0000110000101111",
20496 => "0000110000101111",
20497 => "0000110000110000",
20498 => "0000110000110001",
20499 => "0000110000110010",
20500 => "0000110000110010",
20501 => "0000110000110011",
20502 => "0000110000110100",
20503 => "0000110000110100",
20504 => "0000110000110101",
20505 => "0000110000110110",
20506 => "0000110000110111",
20507 => "0000110000110111",
20508 => "0000110000111000",
20509 => "0000110000111001",
20510 => "0000110000111010",
20511 => "0000110000111010",
20512 => "0000110000111011",
20513 => "0000110000111100",
20514 => "0000110000111100",
20515 => "0000110000111101",
20516 => "0000110000111110",
20517 => "0000110000111111",
20518 => "0000110000111111",
20519 => "0000110001000000",
20520 => "0000110001000001",
20521 => "0000110001000010",
20522 => "0000110001000010",
20523 => "0000110001000011",
20524 => "0000110001000100",
20525 => "0000110001000101",
20526 => "0000110001000101",
20527 => "0000110001000110",
20528 => "0000110001000111",
20529 => "0000110001000111",
20530 => "0000110001001000",
20531 => "0000110001001001",
20532 => "0000110001001010",
20533 => "0000110001001010",
20534 => "0000110001001011",
20535 => "0000110001001100",
20536 => "0000110001001101",
20537 => "0000110001001101",
20538 => "0000110001001110",
20539 => "0000110001001111",
20540 => "0000110001001111",
20541 => "0000110001010000",
20542 => "0000110001010001",
20543 => "0000110001010010",
20544 => "0000110001010010",
20545 => "0000110001010011",
20546 => "0000110001010100",
20547 => "0000110001010101",
20548 => "0000110001010101",
20549 => "0000110001010110",
20550 => "0000110001010111",
20551 => "0000110001011000",
20552 => "0000110001011000",
20553 => "0000110001011001",
20554 => "0000110001011010",
20555 => "0000110001011010",
20556 => "0000110001011011",
20557 => "0000110001011100",
20558 => "0000110001011101",
20559 => "0000110001011101",
20560 => "0000110001011110",
20561 => "0000110001011111",
20562 => "0000110001100000",
20563 => "0000110001100000",
20564 => "0000110001100001",
20565 => "0000110001100010",
20566 => "0000110001100011",
20567 => "0000110001100011",
20568 => "0000110001100100",
20569 => "0000110001100101",
20570 => "0000110001100110",
20571 => "0000110001100110",
20572 => "0000110001100111",
20573 => "0000110001101000",
20574 => "0000110001101000",
20575 => "0000110001101001",
20576 => "0000110001101010",
20577 => "0000110001101011",
20578 => "0000110001101011",
20579 => "0000110001101100",
20580 => "0000110001101101",
20581 => "0000110001101110",
20582 => "0000110001101110",
20583 => "0000110001101111",
20584 => "0000110001110000",
20585 => "0000110001110001",
20586 => "0000110001110001",
20587 => "0000110001110010",
20588 => "0000110001110011",
20589 => "0000110001110100",
20590 => "0000110001110100",
20591 => "0000110001110101",
20592 => "0000110001110110",
20593 => "0000110001110111",
20594 => "0000110001110111",
20595 => "0000110001111000",
20596 => "0000110001111001",
20597 => "0000110001111010",
20598 => "0000110001111010",
20599 => "0000110001111011",
20600 => "0000110001111100",
20601 => "0000110001111100",
20602 => "0000110001111101",
20603 => "0000110001111110",
20604 => "0000110001111111",
20605 => "0000110001111111",
20606 => "0000110010000000",
20607 => "0000110010000001",
20608 => "0000110010000010",
20609 => "0000110010000010",
20610 => "0000110010000011",
20611 => "0000110010000100",
20612 => "0000110010000101",
20613 => "0000110010000101",
20614 => "0000110010000110",
20615 => "0000110010000111",
20616 => "0000110010001000",
20617 => "0000110010001000",
20618 => "0000110010001001",
20619 => "0000110010001010",
20620 => "0000110010001011",
20621 => "0000110010001011",
20622 => "0000110010001100",
20623 => "0000110010001101",
20624 => "0000110010001110",
20625 => "0000110010001110",
20626 => "0000110010001111",
20627 => "0000110010010000",
20628 => "0000110010010001",
20629 => "0000110010010001",
20630 => "0000110010010010",
20631 => "0000110010010011",
20632 => "0000110010010100",
20633 => "0000110010010100",
20634 => "0000110010010101",
20635 => "0000110010010110",
20636 => "0000110010010111",
20637 => "0000110010010111",
20638 => "0000110010011000",
20639 => "0000110010011001",
20640 => "0000110010011010",
20641 => "0000110010011010",
20642 => "0000110010011011",
20643 => "0000110010011100",
20644 => "0000110010011101",
20645 => "0000110010011101",
20646 => "0000110010011110",
20647 => "0000110010011111",
20648 => "0000110010100000",
20649 => "0000110010100000",
20650 => "0000110010100001",
20651 => "0000110010100010",
20652 => "0000110010100011",
20653 => "0000110010100011",
20654 => "0000110010100100",
20655 => "0000110010100101",
20656 => "0000110010100110",
20657 => "0000110010100110",
20658 => "0000110010100111",
20659 => "0000110010101000",
20660 => "0000110010101001",
20661 => "0000110010101001",
20662 => "0000110010101010",
20663 => "0000110010101011",
20664 => "0000110010101100",
20665 => "0000110010101100",
20666 => "0000110010101101",
20667 => "0000110010101110",
20668 => "0000110010101111",
20669 => "0000110010101111",
20670 => "0000110010110000",
20671 => "0000110010110001",
20672 => "0000110010110010",
20673 => "0000110010110010",
20674 => "0000110010110011",
20675 => "0000110010110100",
20676 => "0000110010110101",
20677 => "0000110010110101",
20678 => "0000110010110110",
20679 => "0000110010110111",
20680 => "0000110010111000",
20681 => "0000110010111000",
20682 => "0000110010111001",
20683 => "0000110010111010",
20684 => "0000110010111011",
20685 => "0000110010111011",
20686 => "0000110010111100",
20687 => "0000110010111101",
20688 => "0000110010111110",
20689 => "0000110010111110",
20690 => "0000110010111111",
20691 => "0000110011000000",
20692 => "0000110011000001",
20693 => "0000110011000001",
20694 => "0000110011000010",
20695 => "0000110011000011",
20696 => "0000110011000100",
20697 => "0000110011000101",
20698 => "0000110011000101",
20699 => "0000110011000110",
20700 => "0000110011000111",
20701 => "0000110011001000",
20702 => "0000110011001000",
20703 => "0000110011001001",
20704 => "0000110011001010",
20705 => "0000110011001011",
20706 => "0000110011001011",
20707 => "0000110011001100",
20708 => "0000110011001101",
20709 => "0000110011001110",
20710 => "0000110011001110",
20711 => "0000110011001111",
20712 => "0000110011010000",
20713 => "0000110011010001",
20714 => "0000110011010001",
20715 => "0000110011010010",
20716 => "0000110011010011",
20717 => "0000110011010100",
20718 => "0000110011010100",
20719 => "0000110011010101",
20720 => "0000110011010110",
20721 => "0000110011010111",
20722 => "0000110011011000",
20723 => "0000110011011000",
20724 => "0000110011011001",
20725 => "0000110011011010",
20726 => "0000110011011011",
20727 => "0000110011011011",
20728 => "0000110011011100",
20729 => "0000110011011101",
20730 => "0000110011011110",
20731 => "0000110011011110",
20732 => "0000110011011111",
20733 => "0000110011100000",
20734 => "0000110011100001",
20735 => "0000110011100001",
20736 => "0000110011100010",
20737 => "0000110011100011",
20738 => "0000110011100100",
20739 => "0000110011100101",
20740 => "0000110011100101",
20741 => "0000110011100110",
20742 => "0000110011100111",
20743 => "0000110011101000",
20744 => "0000110011101000",
20745 => "0000110011101001",
20746 => "0000110011101010",
20747 => "0000110011101011",
20748 => "0000110011101011",
20749 => "0000110011101100",
20750 => "0000110011101101",
20751 => "0000110011101110",
20752 => "0000110011101110",
20753 => "0000110011101111",
20754 => "0000110011110000",
20755 => "0000110011110001",
20756 => "0000110011110010",
20757 => "0000110011110010",
20758 => "0000110011110011",
20759 => "0000110011110100",
20760 => "0000110011110101",
20761 => "0000110011110101",
20762 => "0000110011110110",
20763 => "0000110011110111",
20764 => "0000110011111000",
20765 => "0000110011111000",
20766 => "0000110011111001",
20767 => "0000110011111010",
20768 => "0000110011111011",
20769 => "0000110011111100",
20770 => "0000110011111100",
20771 => "0000110011111101",
20772 => "0000110011111110",
20773 => "0000110011111111",
20774 => "0000110011111111",
20775 => "0000110100000000",
20776 => "0000110100000001",
20777 => "0000110100000010",
20778 => "0000110100000010",
20779 => "0000110100000011",
20780 => "0000110100000100",
20781 => "0000110100000101",
20782 => "0000110100000110",
20783 => "0000110100000110",
20784 => "0000110100000111",
20785 => "0000110100001000",
20786 => "0000110100001001",
20787 => "0000110100001001",
20788 => "0000110100001010",
20789 => "0000110100001011",
20790 => "0000110100001100",
20791 => "0000110100001101",
20792 => "0000110100001101",
20793 => "0000110100001110",
20794 => "0000110100001111",
20795 => "0000110100010000",
20796 => "0000110100010000",
20797 => "0000110100010001",
20798 => "0000110100010010",
20799 => "0000110100010011",
20800 => "0000110100010100",
20801 => "0000110100010100",
20802 => "0000110100010101",
20803 => "0000110100010110",
20804 => "0000110100010111",
20805 => "0000110100010111",
20806 => "0000110100011000",
20807 => "0000110100011001",
20808 => "0000110100011010",
20809 => "0000110100011010",
20810 => "0000110100011011",
20811 => "0000110100011100",
20812 => "0000110100011101",
20813 => "0000110100011110",
20814 => "0000110100011110",
20815 => "0000110100011111",
20816 => "0000110100100000",
20817 => "0000110100100001",
20818 => "0000110100100001",
20819 => "0000110100100010",
20820 => "0000110100100011",
20821 => "0000110100100100",
20822 => "0000110100100101",
20823 => "0000110100100101",
20824 => "0000110100100110",
20825 => "0000110100100111",
20826 => "0000110100101000",
20827 => "0000110100101001",
20828 => "0000110100101001",
20829 => "0000110100101010",
20830 => "0000110100101011",
20831 => "0000110100101100",
20832 => "0000110100101100",
20833 => "0000110100101101",
20834 => "0000110100101110",
20835 => "0000110100101111",
20836 => "0000110100110000",
20837 => "0000110100110000",
20838 => "0000110100110001",
20839 => "0000110100110010",
20840 => "0000110100110011",
20841 => "0000110100110011",
20842 => "0000110100110100",
20843 => "0000110100110101",
20844 => "0000110100110110",
20845 => "0000110100110111",
20846 => "0000110100110111",
20847 => "0000110100111000",
20848 => "0000110100111001",
20849 => "0000110100111010",
20850 => "0000110100111010",
20851 => "0000110100111011",
20852 => "0000110100111100",
20853 => "0000110100111101",
20854 => "0000110100111110",
20855 => "0000110100111110",
20856 => "0000110100111111",
20857 => "0000110101000000",
20858 => "0000110101000001",
20859 => "0000110101000010",
20860 => "0000110101000010",
20861 => "0000110101000011",
20862 => "0000110101000100",
20863 => "0000110101000101",
20864 => "0000110101000101",
20865 => "0000110101000110",
20866 => "0000110101000111",
20867 => "0000110101001000",
20868 => "0000110101001001",
20869 => "0000110101001001",
20870 => "0000110101001010",
20871 => "0000110101001011",
20872 => "0000110101001100",
20873 => "0000110101001101",
20874 => "0000110101001101",
20875 => "0000110101001110",
20876 => "0000110101001111",
20877 => "0000110101010000",
20878 => "0000110101010001",
20879 => "0000110101010001",
20880 => "0000110101010010",
20881 => "0000110101010011",
20882 => "0000110101010100",
20883 => "0000110101010100",
20884 => "0000110101010101",
20885 => "0000110101010110",
20886 => "0000110101010111",
20887 => "0000110101011000",
20888 => "0000110101011000",
20889 => "0000110101011001",
20890 => "0000110101011010",
20891 => "0000110101011011",
20892 => "0000110101011100",
20893 => "0000110101011100",
20894 => "0000110101011101",
20895 => "0000110101011110",
20896 => "0000110101011111",
20897 => "0000110101100000",
20898 => "0000110101100000",
20899 => "0000110101100001",
20900 => "0000110101100010",
20901 => "0000110101100011",
20902 => "0000110101100100",
20903 => "0000110101100100",
20904 => "0000110101100101",
20905 => "0000110101100110",
20906 => "0000110101100111",
20907 => "0000110101100111",
20908 => "0000110101101000",
20909 => "0000110101101001",
20910 => "0000110101101010",
20911 => "0000110101101011",
20912 => "0000110101101011",
20913 => "0000110101101100",
20914 => "0000110101101101",
20915 => "0000110101101110",
20916 => "0000110101101111",
20917 => "0000110101101111",
20918 => "0000110101110000",
20919 => "0000110101110001",
20920 => "0000110101110010",
20921 => "0000110101110011",
20922 => "0000110101110011",
20923 => "0000110101110100",
20924 => "0000110101110101",
20925 => "0000110101110110",
20926 => "0000110101110111",
20927 => "0000110101110111",
20928 => "0000110101111000",
20929 => "0000110101111001",
20930 => "0000110101111010",
20931 => "0000110101111011",
20932 => "0000110101111011",
20933 => "0000110101111100",
20934 => "0000110101111101",
20935 => "0000110101111110",
20936 => "0000110101111111",
20937 => "0000110101111111",
20938 => "0000110110000000",
20939 => "0000110110000001",
20940 => "0000110110000010",
20941 => "0000110110000011",
20942 => "0000110110000011",
20943 => "0000110110000100",
20944 => "0000110110000101",
20945 => "0000110110000110",
20946 => "0000110110000111",
20947 => "0000110110000111",
20948 => "0000110110001000",
20949 => "0000110110001001",
20950 => "0000110110001010",
20951 => "0000110110001011",
20952 => "0000110110001011",
20953 => "0000110110001100",
20954 => "0000110110001101",
20955 => "0000110110001110",
20956 => "0000110110001111",
20957 => "0000110110001111",
20958 => "0000110110010000",
20959 => "0000110110010001",
20960 => "0000110110010010",
20961 => "0000110110010011",
20962 => "0000110110010011",
20963 => "0000110110010100",
20964 => "0000110110010101",
20965 => "0000110110010110",
20966 => "0000110110010111",
20967 => "0000110110010111",
20968 => "0000110110011000",
20969 => "0000110110011001",
20970 => "0000110110011010",
20971 => "0000110110011011",
20972 => "0000110110011011",
20973 => "0000110110011100",
20974 => "0000110110011101",
20975 => "0000110110011110",
20976 => "0000110110011111",
20977 => "0000110110011111",
20978 => "0000110110100000",
20979 => "0000110110100001",
20980 => "0000110110100010",
20981 => "0000110110100011",
20982 => "0000110110100100",
20983 => "0000110110100100",
20984 => "0000110110100101",
20985 => "0000110110100110",
20986 => "0000110110100111",
20987 => "0000110110101000",
20988 => "0000110110101000",
20989 => "0000110110101001",
20990 => "0000110110101010",
20991 => "0000110110101011",
20992 => "0000110110101100",
20993 => "0000110110101100",
20994 => "0000110110101101",
20995 => "0000110110101110",
20996 => "0000110110101111",
20997 => "0000110110110000",
20998 => "0000110110110000",
20999 => "0000110110110001",
21000 => "0000110110110010",
21001 => "0000110110110011",
21002 => "0000110110110100",
21003 => "0000110110110101",
21004 => "0000110110110101",
21005 => "0000110110110110",
21006 => "0000110110110111",
21007 => "0000110110111000",
21008 => "0000110110111001",
21009 => "0000110110111001",
21010 => "0000110110111010",
21011 => "0000110110111011",
21012 => "0000110110111100",
21013 => "0000110110111101",
21014 => "0000110110111101",
21015 => "0000110110111110",
21016 => "0000110110111111",
21017 => "0000110111000000",
21018 => "0000110111000001",
21019 => "0000110111000010",
21020 => "0000110111000010",
21021 => "0000110111000011",
21022 => "0000110111000100",
21023 => "0000110111000101",
21024 => "0000110111000110",
21025 => "0000110111000110",
21026 => "0000110111000111",
21027 => "0000110111001000",
21028 => "0000110111001001",
21029 => "0000110111001010",
21030 => "0000110111001010",
21031 => "0000110111001011",
21032 => "0000110111001100",
21033 => "0000110111001101",
21034 => "0000110111001110",
21035 => "0000110111001111",
21036 => "0000110111001111",
21037 => "0000110111010000",
21038 => "0000110111010001",
21039 => "0000110111010010",
21040 => "0000110111010011",
21041 => "0000110111010011",
21042 => "0000110111010100",
21043 => "0000110111010101",
21044 => "0000110111010110",
21045 => "0000110111010111",
21046 => "0000110111011000",
21047 => "0000110111011000",
21048 => "0000110111011001",
21049 => "0000110111011010",
21050 => "0000110111011011",
21051 => "0000110111011100",
21052 => "0000110111011100",
21053 => "0000110111011101",
21054 => "0000110111011110",
21055 => "0000110111011111",
21056 => "0000110111100000",
21057 => "0000110111100001",
21058 => "0000110111100001",
21059 => "0000110111100010",
21060 => "0000110111100011",
21061 => "0000110111100100",
21062 => "0000110111100101",
21063 => "0000110111100101",
21064 => "0000110111100110",
21065 => "0000110111100111",
21066 => "0000110111101000",
21067 => "0000110111101001",
21068 => "0000110111101010",
21069 => "0000110111101010",
21070 => "0000110111101011",
21071 => "0000110111101100",
21072 => "0000110111101101",
21073 => "0000110111101110",
21074 => "0000110111101111",
21075 => "0000110111101111",
21076 => "0000110111110000",
21077 => "0000110111110001",
21078 => "0000110111110010",
21079 => "0000110111110011",
21080 => "0000110111110011",
21081 => "0000110111110100",
21082 => "0000110111110101",
21083 => "0000110111110110",
21084 => "0000110111110111",
21085 => "0000110111111000",
21086 => "0000110111111000",
21087 => "0000110111111001",
21088 => "0000110111111010",
21089 => "0000110111111011",
21090 => "0000110111111100",
21091 => "0000110111111101",
21092 => "0000110111111101",
21093 => "0000110111111110",
21094 => "0000110111111111",
21095 => "0000111000000000",
21096 => "0000111000000001",
21097 => "0000111000000010",
21098 => "0000111000000010",
21099 => "0000111000000011",
21100 => "0000111000000100",
21101 => "0000111000000101",
21102 => "0000111000000110",
21103 => "0000111000000110",
21104 => "0000111000000111",
21105 => "0000111000001000",
21106 => "0000111000001001",
21107 => "0000111000001010",
21108 => "0000111000001011",
21109 => "0000111000001011",
21110 => "0000111000001100",
21111 => "0000111000001101",
21112 => "0000111000001110",
21113 => "0000111000001111",
21114 => "0000111000010000",
21115 => "0000111000010000",
21116 => "0000111000010001",
21117 => "0000111000010010",
21118 => "0000111000010011",
21119 => "0000111000010100",
21120 => "0000111000010101",
21121 => "0000111000010101",
21122 => "0000111000010110",
21123 => "0000111000010111",
21124 => "0000111000011000",
21125 => "0000111000011001",
21126 => "0000111000011010",
21127 => "0000111000011010",
21128 => "0000111000011011",
21129 => "0000111000011100",
21130 => "0000111000011101",
21131 => "0000111000011110",
21132 => "0000111000011111",
21133 => "0000111000011111",
21134 => "0000111000100000",
21135 => "0000111000100001",
21136 => "0000111000100010",
21137 => "0000111000100011",
21138 => "0000111000100100",
21139 => "0000111000100100",
21140 => "0000111000100101",
21141 => "0000111000100110",
21142 => "0000111000100111",
21143 => "0000111000101000",
21144 => "0000111000101001",
21145 => "0000111000101001",
21146 => "0000111000101010",
21147 => "0000111000101011",
21148 => "0000111000101100",
21149 => "0000111000101101",
21150 => "0000111000101110",
21151 => "0000111000101110",
21152 => "0000111000101111",
21153 => "0000111000110000",
21154 => "0000111000110001",
21155 => "0000111000110010",
21156 => "0000111000110011",
21157 => "0000111000110011",
21158 => "0000111000110100",
21159 => "0000111000110101",
21160 => "0000111000110110",
21161 => "0000111000110111",
21162 => "0000111000111000",
21163 => "0000111000111001",
21164 => "0000111000111001",
21165 => "0000111000111010",
21166 => "0000111000111011",
21167 => "0000111000111100",
21168 => "0000111000111101",
21169 => "0000111000111110",
21170 => "0000111000111110",
21171 => "0000111000111111",
21172 => "0000111001000000",
21173 => "0000111001000001",
21174 => "0000111001000010",
21175 => "0000111001000011",
21176 => "0000111001000011",
21177 => "0000111001000100",
21178 => "0000111001000101",
21179 => "0000111001000110",
21180 => "0000111001000111",
21181 => "0000111001001000",
21182 => "0000111001001001",
21183 => "0000111001001001",
21184 => "0000111001001010",
21185 => "0000111001001011",
21186 => "0000111001001100",
21187 => "0000111001001101",
21188 => "0000111001001110",
21189 => "0000111001001110",
21190 => "0000111001001111",
21191 => "0000111001010000",
21192 => "0000111001010001",
21193 => "0000111001010010",
21194 => "0000111001010011",
21195 => "0000111001010011",
21196 => "0000111001010100",
21197 => "0000111001010101",
21198 => "0000111001010110",
21199 => "0000111001010111",
21200 => "0000111001011000",
21201 => "0000111001011001",
21202 => "0000111001011001",
21203 => "0000111001011010",
21204 => "0000111001011011",
21205 => "0000111001011100",
21206 => "0000111001011101",
21207 => "0000111001011110",
21208 => "0000111001011110",
21209 => "0000111001011111",
21210 => "0000111001100000",
21211 => "0000111001100001",
21212 => "0000111001100010",
21213 => "0000111001100011",
21214 => "0000111001100100",
21215 => "0000111001100100",
21216 => "0000111001100101",
21217 => "0000111001100110",
21218 => "0000111001100111",
21219 => "0000111001101000",
21220 => "0000111001101001",
21221 => "0000111001101010",
21222 => "0000111001101010",
21223 => "0000111001101011",
21224 => "0000111001101100",
21225 => "0000111001101101",
21226 => "0000111001101110",
21227 => "0000111001101111",
21228 => "0000111001101111",
21229 => "0000111001110000",
21230 => "0000111001110001",
21231 => "0000111001110010",
21232 => "0000111001110011",
21233 => "0000111001110100",
21234 => "0000111001110101",
21235 => "0000111001110101",
21236 => "0000111001110110",
21237 => "0000111001110111",
21238 => "0000111001111000",
21239 => "0000111001111001",
21240 => "0000111001111010",
21241 => "0000111001111011",
21242 => "0000111001111011",
21243 => "0000111001111100",
21244 => "0000111001111101",
21245 => "0000111001111110",
21246 => "0000111001111111",
21247 => "0000111010000000",
21248 => "0000111010000001",
21249 => "0000111010000001",
21250 => "0000111010000010",
21251 => "0000111010000011",
21252 => "0000111010000100",
21253 => "0000111010000101",
21254 => "0000111010000110",
21255 => "0000111010000111",
21256 => "0000111010000111",
21257 => "0000111010001000",
21258 => "0000111010001001",
21259 => "0000111010001010",
21260 => "0000111010001011",
21261 => "0000111010001100",
21262 => "0000111010001101",
21263 => "0000111010001101",
21264 => "0000111010001110",
21265 => "0000111010001111",
21266 => "0000111010010000",
21267 => "0000111010010001",
21268 => "0000111010010010",
21269 => "0000111010010011",
21270 => "0000111010010011",
21271 => "0000111010010100",
21272 => "0000111010010101",
21273 => "0000111010010110",
21274 => "0000111010010111",
21275 => "0000111010011000",
21276 => "0000111010011001",
21277 => "0000111010011001",
21278 => "0000111010011010",
21279 => "0000111010011011",
21280 => "0000111010011100",
21281 => "0000111010011101",
21282 => "0000111010011110",
21283 => "0000111010011111",
21284 => "0000111010011111",
21285 => "0000111010100000",
21286 => "0000111010100001",
21287 => "0000111010100010",
21288 => "0000111010100011",
21289 => "0000111010100100",
21290 => "0000111010100101",
21291 => "0000111010100101",
21292 => "0000111010100110",
21293 => "0000111010100111",
21294 => "0000111010101000",
21295 => "0000111010101001",
21296 => "0000111010101010",
21297 => "0000111010101011",
21298 => "0000111010101100",
21299 => "0000111010101100",
21300 => "0000111010101101",
21301 => "0000111010101110",
21302 => "0000111010101111",
21303 => "0000111010110000",
21304 => "0000111010110001",
21305 => "0000111010110010",
21306 => "0000111010110010",
21307 => "0000111010110011",
21308 => "0000111010110100",
21309 => "0000111010110101",
21310 => "0000111010110110",
21311 => "0000111010110111",
21312 => "0000111010111000",
21313 => "0000111010111001",
21314 => "0000111010111001",
21315 => "0000111010111010",
21316 => "0000111010111011",
21317 => "0000111010111100",
21318 => "0000111010111101",
21319 => "0000111010111110",
21320 => "0000111010111111",
21321 => "0000111010111111",
21322 => "0000111011000000",
21323 => "0000111011000001",
21324 => "0000111011000010",
21325 => "0000111011000011",
21326 => "0000111011000100",
21327 => "0000111011000101",
21328 => "0000111011000110",
21329 => "0000111011000110",
21330 => "0000111011000111",
21331 => "0000111011001000",
21332 => "0000111011001001",
21333 => "0000111011001010",
21334 => "0000111011001011",
21335 => "0000111011001100",
21336 => "0000111011001101",
21337 => "0000111011001101",
21338 => "0000111011001110",
21339 => "0000111011001111",
21340 => "0000111011010000",
21341 => "0000111011010001",
21342 => "0000111011010010",
21343 => "0000111011010011",
21344 => "0000111011010100",
21345 => "0000111011010100",
21346 => "0000111011010101",
21347 => "0000111011010110",
21348 => "0000111011010111",
21349 => "0000111011011000",
21350 => "0000111011011001",
21351 => "0000111011011010",
21352 => "0000111011011010",
21353 => "0000111011011011",
21354 => "0000111011011100",
21355 => "0000111011011101",
21356 => "0000111011011110",
21357 => "0000111011011111",
21358 => "0000111011100000",
21359 => "0000111011100001",
21360 => "0000111011100001",
21361 => "0000111011100010",
21362 => "0000111011100011",
21363 => "0000111011100100",
21364 => "0000111011100101",
21365 => "0000111011100110",
21366 => "0000111011100111",
21367 => "0000111011101000",
21368 => "0000111011101001",
21369 => "0000111011101001",
21370 => "0000111011101010",
21371 => "0000111011101011",
21372 => "0000111011101100",
21373 => "0000111011101101",
21374 => "0000111011101110",
21375 => "0000111011101111",
21376 => "0000111011110000",
21377 => "0000111011110000",
21378 => "0000111011110001",
21379 => "0000111011110010",
21380 => "0000111011110011",
21381 => "0000111011110100",
21382 => "0000111011110101",
21383 => "0000111011110110",
21384 => "0000111011110111",
21385 => "0000111011110111",
21386 => "0000111011111000",
21387 => "0000111011111001",
21388 => "0000111011111010",
21389 => "0000111011111011",
21390 => "0000111011111100",
21391 => "0000111011111101",
21392 => "0000111011111110",
21393 => "0000111011111111",
21394 => "0000111011111111",
21395 => "0000111100000000",
21396 => "0000111100000001",
21397 => "0000111100000010",
21398 => "0000111100000011",
21399 => "0000111100000100",
21400 => "0000111100000101",
21401 => "0000111100000110",
21402 => "0000111100000110",
21403 => "0000111100000111",
21404 => "0000111100001000",
21405 => "0000111100001001",
21406 => "0000111100001010",
21407 => "0000111100001011",
21408 => "0000111100001100",
21409 => "0000111100001101",
21410 => "0000111100001110",
21411 => "0000111100001110",
21412 => "0000111100001111",
21413 => "0000111100010000",
21414 => "0000111100010001",
21415 => "0000111100010010",
21416 => "0000111100010011",
21417 => "0000111100010100",
21418 => "0000111100010101",
21419 => "0000111100010110",
21420 => "0000111100010110",
21421 => "0000111100010111",
21422 => "0000111100011000",
21423 => "0000111100011001",
21424 => "0000111100011010",
21425 => "0000111100011011",
21426 => "0000111100011100",
21427 => "0000111100011101",
21428 => "0000111100011110",
21429 => "0000111100011110",
21430 => "0000111100011111",
21431 => "0000111100100000",
21432 => "0000111100100001",
21433 => "0000111100100010",
21434 => "0000111100100011",
21435 => "0000111100100100",
21436 => "0000111100100101",
21437 => "0000111100100110",
21438 => "0000111100100110",
21439 => "0000111100100111",
21440 => "0000111100101000",
21441 => "0000111100101001",
21442 => "0000111100101010",
21443 => "0000111100101011",
21444 => "0000111100101100",
21445 => "0000111100101101",
21446 => "0000111100101110",
21447 => "0000111100101110",
21448 => "0000111100101111",
21449 => "0000111100110000",
21450 => "0000111100110001",
21451 => "0000111100110010",
21452 => "0000111100110011",
21453 => "0000111100110100",
21454 => "0000111100110101",
21455 => "0000111100110110",
21456 => "0000111100110110",
21457 => "0000111100110111",
21458 => "0000111100111000",
21459 => "0000111100111001",
21460 => "0000111100111010",
21461 => "0000111100111011",
21462 => "0000111100111100",
21463 => "0000111100111101",
21464 => "0000111100111110",
21465 => "0000111100111111",
21466 => "0000111100111111",
21467 => "0000111101000000",
21468 => "0000111101000001",
21469 => "0000111101000010",
21470 => "0000111101000011",
21471 => "0000111101000100",
21472 => "0000111101000101",
21473 => "0000111101000110",
21474 => "0000111101000111",
21475 => "0000111101001000",
21476 => "0000111101001000",
21477 => "0000111101001001",
21478 => "0000111101001010",
21479 => "0000111101001011",
21480 => "0000111101001100",
21481 => "0000111101001101",
21482 => "0000111101001110",
21483 => "0000111101001111",
21484 => "0000111101010000",
21485 => "0000111101010000",
21486 => "0000111101010001",
21487 => "0000111101010010",
21488 => "0000111101010011",
21489 => "0000111101010100",
21490 => "0000111101010101",
21491 => "0000111101010110",
21492 => "0000111101010111",
21493 => "0000111101011000",
21494 => "0000111101011001",
21495 => "0000111101011010",
21496 => "0000111101011010",
21497 => "0000111101011011",
21498 => "0000111101011100",
21499 => "0000111101011101",
21500 => "0000111101011110",
21501 => "0000111101011111",
21502 => "0000111101100000",
21503 => "0000111101100001",
21504 => "0000111101100010",
21505 => "0000111101100011",
21506 => "0000111101100011",
21507 => "0000111101100100",
21508 => "0000111101100101",
21509 => "0000111101100110",
21510 => "0000111101100111",
21511 => "0000111101101000",
21512 => "0000111101101001",
21513 => "0000111101101010",
21514 => "0000111101101011",
21515 => "0000111101101100",
21516 => "0000111101101100",
21517 => "0000111101101101",
21518 => "0000111101101110",
21519 => "0000111101101111",
21520 => "0000111101110000",
21521 => "0000111101110001",
21522 => "0000111101110010",
21523 => "0000111101110011",
21524 => "0000111101110100",
21525 => "0000111101110101",
21526 => "0000111101110110",
21527 => "0000111101110110",
21528 => "0000111101110111",
21529 => "0000111101111000",
21530 => "0000111101111001",
21531 => "0000111101111010",
21532 => "0000111101111011",
21533 => "0000111101111100",
21534 => "0000111101111101",
21535 => "0000111101111110",
21536 => "0000111101111111",
21537 => "0000111110000000",
21538 => "0000111110000000",
21539 => "0000111110000001",
21540 => "0000111110000010",
21541 => "0000111110000011",
21542 => "0000111110000100",
21543 => "0000111110000101",
21544 => "0000111110000110",
21545 => "0000111110000111",
21546 => "0000111110001000",
21547 => "0000111110001001",
21548 => "0000111110001010",
21549 => "0000111110001010",
21550 => "0000111110001011",
21551 => "0000111110001100",
21552 => "0000111110001101",
21553 => "0000111110001110",
21554 => "0000111110001111",
21555 => "0000111110010000",
21556 => "0000111110010001",
21557 => "0000111110010010",
21558 => "0000111110010011",
21559 => "0000111110010100",
21560 => "0000111110010101",
21561 => "0000111110010101",
21562 => "0000111110010110",
21563 => "0000111110010111",
21564 => "0000111110011000",
21565 => "0000111110011001",
21566 => "0000111110011010",
21567 => "0000111110011011",
21568 => "0000111110011100",
21569 => "0000111110011101",
21570 => "0000111110011110",
21571 => "0000111110011111",
21572 => "0000111110100000",
21573 => "0000111110100000",
21574 => "0000111110100001",
21575 => "0000111110100010",
21576 => "0000111110100011",
21577 => "0000111110100100",
21578 => "0000111110100101",
21579 => "0000111110100110",
21580 => "0000111110100111",
21581 => "0000111110101000",
21582 => "0000111110101001",
21583 => "0000111110101010",
21584 => "0000111110101011",
21585 => "0000111110101011",
21586 => "0000111110101100",
21587 => "0000111110101101",
21588 => "0000111110101110",
21589 => "0000111110101111",
21590 => "0000111110110000",
21591 => "0000111110110001",
21592 => "0000111110110010",
21593 => "0000111110110011",
21594 => "0000111110110100",
21595 => "0000111110110101",
21596 => "0000111110110110",
21597 => "0000111110110111",
21598 => "0000111110110111",
21599 => "0000111110111000",
21600 => "0000111110111001",
21601 => "0000111110111010",
21602 => "0000111110111011",
21603 => "0000111110111100",
21604 => "0000111110111101",
21605 => "0000111110111110",
21606 => "0000111110111111",
21607 => "0000111111000000",
21608 => "0000111111000001",
21609 => "0000111111000010",
21610 => "0000111111000011",
21611 => "0000111111000011",
21612 => "0000111111000100",
21613 => "0000111111000101",
21614 => "0000111111000110",
21615 => "0000111111000111",
21616 => "0000111111001000",
21617 => "0000111111001001",
21618 => "0000111111001010",
21619 => "0000111111001011",
21620 => "0000111111001100",
21621 => "0000111111001101",
21622 => "0000111111001110",
21623 => "0000111111001111",
21624 => "0000111111001111",
21625 => "0000111111010000",
21626 => "0000111111010001",
21627 => "0000111111010010",
21628 => "0000111111010011",
21629 => "0000111111010100",
21630 => "0000111111010101",
21631 => "0000111111010110",
21632 => "0000111111010111",
21633 => "0000111111011000",
21634 => "0000111111011001",
21635 => "0000111111011010",
21636 => "0000111111011011",
21637 => "0000111111011100",
21638 => "0000111111011100",
21639 => "0000111111011101",
21640 => "0000111111011110",
21641 => "0000111111011111",
21642 => "0000111111100000",
21643 => "0000111111100001",
21644 => "0000111111100010",
21645 => "0000111111100011",
21646 => "0000111111100100",
21647 => "0000111111100101",
21648 => "0000111111100110",
21649 => "0000111111100111",
21650 => "0000111111101000",
21651 => "0000111111101001",
21652 => "0000111111101010",
21653 => "0000111111101010",
21654 => "0000111111101011",
21655 => "0000111111101100",
21656 => "0000111111101101",
21657 => "0000111111101110",
21658 => "0000111111101111",
21659 => "0000111111110000",
21660 => "0000111111110001",
21661 => "0000111111110010",
21662 => "0000111111110011",
21663 => "0000111111110100",
21664 => "0000111111110101",
21665 => "0000111111110110",
21666 => "0000111111110111",
21667 => "0000111111111000",
21668 => "0000111111111000",
21669 => "0000111111111001",
21670 => "0000111111111010",
21671 => "0000111111111011",
21672 => "0000111111111100",
21673 => "0000111111111101",
21674 => "0000111111111110",
21675 => "0000111111111111",
21676 => "0001000000000000",
21677 => "0001000000000001",
21678 => "0001000000000010",
21679 => "0001000000000011",
21680 => "0001000000000100",
21681 => "0001000000000101",
21682 => "0001000000000110",
21683 => "0001000000000111",
21684 => "0001000000000111",
21685 => "0001000000001000",
21686 => "0001000000001001",
21687 => "0001000000001010",
21688 => "0001000000001011",
21689 => "0001000000001100",
21690 => "0001000000001101",
21691 => "0001000000001110",
21692 => "0001000000001111",
21693 => "0001000000010000",
21694 => "0001000000010001",
21695 => "0001000000010010",
21696 => "0001000000010011",
21697 => "0001000000010100",
21698 => "0001000000010101",
21699 => "0001000000010110",
21700 => "0001000000010111",
21701 => "0001000000010111",
21702 => "0001000000011000",
21703 => "0001000000011001",
21704 => "0001000000011010",
21705 => "0001000000011011",
21706 => "0001000000011100",
21707 => "0001000000011101",
21708 => "0001000000011110",
21709 => "0001000000011111",
21710 => "0001000000100000",
21711 => "0001000000100001",
21712 => "0001000000100010",
21713 => "0001000000100011",
21714 => "0001000000100100",
21715 => "0001000000100101",
21716 => "0001000000100110",
21717 => "0001000000100111",
21718 => "0001000000101000",
21719 => "0001000000101000",
21720 => "0001000000101001",
21721 => "0001000000101010",
21722 => "0001000000101011",
21723 => "0001000000101100",
21724 => "0001000000101101",
21725 => "0001000000101110",
21726 => "0001000000101111",
21727 => "0001000000110000",
21728 => "0001000000110001",
21729 => "0001000000110010",
21730 => "0001000000110011",
21731 => "0001000000110100",
21732 => "0001000000110101",
21733 => "0001000000110110",
21734 => "0001000000110111",
21735 => "0001000000111000",
21736 => "0001000000111001",
21737 => "0001000000111010",
21738 => "0001000000111010",
21739 => "0001000000111011",
21740 => "0001000000111100",
21741 => "0001000000111101",
21742 => "0001000000111110",
21743 => "0001000000111111",
21744 => "0001000001000000",
21745 => "0001000001000001",
21746 => "0001000001000010",
21747 => "0001000001000011",
21748 => "0001000001000100",
21749 => "0001000001000101",
21750 => "0001000001000110",
21751 => "0001000001000111",
21752 => "0001000001001000",
21753 => "0001000001001001",
21754 => "0001000001001010",
21755 => "0001000001001011",
21756 => "0001000001001100",
21757 => "0001000001001101",
21758 => "0001000001001110",
21759 => "0001000001001110",
21760 => "0001000001001111",
21761 => "0001000001010000",
21762 => "0001000001010001",
21763 => "0001000001010010",
21764 => "0001000001010011",
21765 => "0001000001010100",
21766 => "0001000001010101",
21767 => "0001000001010110",
21768 => "0001000001010111",
21769 => "0001000001011000",
21770 => "0001000001011001",
21771 => "0001000001011010",
21772 => "0001000001011011",
21773 => "0001000001011100",
21774 => "0001000001011101",
21775 => "0001000001011110",
21776 => "0001000001011111",
21777 => "0001000001100000",
21778 => "0001000001100001",
21779 => "0001000001100010",
21780 => "0001000001100011",
21781 => "0001000001100100",
21782 => "0001000001100100",
21783 => "0001000001100101",
21784 => "0001000001100110",
21785 => "0001000001100111",
21786 => "0001000001101000",
21787 => "0001000001101001",
21788 => "0001000001101010",
21789 => "0001000001101011",
21790 => "0001000001101100",
21791 => "0001000001101101",
21792 => "0001000001101110",
21793 => "0001000001101111",
21794 => "0001000001110000",
21795 => "0001000001110001",
21796 => "0001000001110010",
21797 => "0001000001110011",
21798 => "0001000001110100",
21799 => "0001000001110101",
21800 => "0001000001110110",
21801 => "0001000001110111",
21802 => "0001000001111000",
21803 => "0001000001111001",
21804 => "0001000001111010",
21805 => "0001000001111011",
21806 => "0001000001111100",
21807 => "0001000001111101",
21808 => "0001000001111101",
21809 => "0001000001111110",
21810 => "0001000001111111",
21811 => "0001000010000000",
21812 => "0001000010000001",
21813 => "0001000010000010",
21814 => "0001000010000011",
21815 => "0001000010000100",
21816 => "0001000010000101",
21817 => "0001000010000110",
21818 => "0001000010000111",
21819 => "0001000010001000",
21820 => "0001000010001001",
21821 => "0001000010001010",
21822 => "0001000010001011",
21823 => "0001000010001100",
21824 => "0001000010001101",
21825 => "0001000010001110",
21826 => "0001000010001111",
21827 => "0001000010010000",
21828 => "0001000010010001",
21829 => "0001000010010010",
21830 => "0001000010010011",
21831 => "0001000010010100",
21832 => "0001000010010101",
21833 => "0001000010010110",
21834 => "0001000010010111",
21835 => "0001000010011000",
21836 => "0001000010011001",
21837 => "0001000010011010",
21838 => "0001000010011011",
21839 => "0001000010011011",
21840 => "0001000010011100",
21841 => "0001000010011101",
21842 => "0001000010011110",
21843 => "0001000010011111",
21844 => "0001000010100000",
21845 => "0001000010100001",
21846 => "0001000010100010",
21847 => "0001000010100011",
21848 => "0001000010100100",
21849 => "0001000010100101",
21850 => "0001000010100110",
21851 => "0001000010100111",
21852 => "0001000010101000",
21853 => "0001000010101001",
21854 => "0001000010101010",
21855 => "0001000010101011",
21856 => "0001000010101100",
21857 => "0001000010101101",
21858 => "0001000010101110",
21859 => "0001000010101111",
21860 => "0001000010110000",
21861 => "0001000010110001",
21862 => "0001000010110010",
21863 => "0001000010110011",
21864 => "0001000010110100",
21865 => "0001000010110101",
21866 => "0001000010110110",
21867 => "0001000010110111",
21868 => "0001000010111000",
21869 => "0001000010111001",
21870 => "0001000010111010",
21871 => "0001000010111011",
21872 => "0001000010111100",
21873 => "0001000010111101",
21874 => "0001000010111110",
21875 => "0001000010111111",
21876 => "0001000011000000",
21877 => "0001000011000001",
21878 => "0001000011000010",
21879 => "0001000011000010",
21880 => "0001000011000011",
21881 => "0001000011000100",
21882 => "0001000011000101",
21883 => "0001000011000110",
21884 => "0001000011000111",
21885 => "0001000011001000",
21886 => "0001000011001001",
21887 => "0001000011001010",
21888 => "0001000011001011",
21889 => "0001000011001100",
21890 => "0001000011001101",
21891 => "0001000011001110",
21892 => "0001000011001111",
21893 => "0001000011010000",
21894 => "0001000011010001",
21895 => "0001000011010010",
21896 => "0001000011010011",
21897 => "0001000011010100",
21898 => "0001000011010101",
21899 => "0001000011010110",
21900 => "0001000011010111",
21901 => "0001000011011000",
21902 => "0001000011011001",
21903 => "0001000011011010",
21904 => "0001000011011011",
21905 => "0001000011011100",
21906 => "0001000011011101",
21907 => "0001000011011110",
21908 => "0001000011011111",
21909 => "0001000011100000",
21910 => "0001000011100001",
21911 => "0001000011100010",
21912 => "0001000011100011",
21913 => "0001000011100100",
21914 => "0001000011100101",
21915 => "0001000011100110",
21916 => "0001000011100111",
21917 => "0001000011101000",
21918 => "0001000011101001",
21919 => "0001000011101010",
21920 => "0001000011101011",
21921 => "0001000011101100",
21922 => "0001000011101101",
21923 => "0001000011101110",
21924 => "0001000011101111",
21925 => "0001000011110000",
21926 => "0001000011110001",
21927 => "0001000011110010",
21928 => "0001000011110011",
21929 => "0001000011110100",
21930 => "0001000011110101",
21931 => "0001000011110110",
21932 => "0001000011110111",
21933 => "0001000011111000",
21934 => "0001000011111001",
21935 => "0001000011111010",
21936 => "0001000011111011",
21937 => "0001000011111100",
21938 => "0001000011111101",
21939 => "0001000011111110",
21940 => "0001000011111111",
21941 => "0001000100000000",
21942 => "0001000100000001",
21943 => "0001000100000010",
21944 => "0001000100000011",
21945 => "0001000100000100",
21946 => "0001000100000101",
21947 => "0001000100000110",
21948 => "0001000100000111",
21949 => "0001000100001000",
21950 => "0001000100001001",
21951 => "0001000100001010",
21952 => "0001000100001011",
21953 => "0001000100001100",
21954 => "0001000100001101",
21955 => "0001000100001101",
21956 => "0001000100001110",
21957 => "0001000100001111",
21958 => "0001000100010000",
21959 => "0001000100010001",
21960 => "0001000100010010",
21961 => "0001000100010011",
21962 => "0001000100010100",
21963 => "0001000100010101",
21964 => "0001000100010110",
21965 => "0001000100010111",
21966 => "0001000100011000",
21967 => "0001000100011001",
21968 => "0001000100011010",
21969 => "0001000100011011",
21970 => "0001000100011100",
21971 => "0001000100011101",
21972 => "0001000100011110",
21973 => "0001000100011111",
21974 => "0001000100100000",
21975 => "0001000100100001",
21976 => "0001000100100010",
21977 => "0001000100100011",
21978 => "0001000100100100",
21979 => "0001000100100101",
21980 => "0001000100100110",
21981 => "0001000100100111",
21982 => "0001000100101000",
21983 => "0001000100101001",
21984 => "0001000100101010",
21985 => "0001000100101011",
21986 => "0001000100101100",
21987 => "0001000100101101",
21988 => "0001000100101110",
21989 => "0001000100101111",
21990 => "0001000100110000",
21991 => "0001000100110001",
21992 => "0001000100110010",
21993 => "0001000100110011",
21994 => "0001000100110100",
21995 => "0001000100110101",
21996 => "0001000100110110",
21997 => "0001000100110111",
21998 => "0001000100111000",
21999 => "0001000100111001",
22000 => "0001000100111010",
22001 => "0001000100111011",
22002 => "0001000100111100",
22003 => "0001000100111101",
22004 => "0001000100111110",
22005 => "0001000101000000",
22006 => "0001000101000001",
22007 => "0001000101000010",
22008 => "0001000101000011",
22009 => "0001000101000100",
22010 => "0001000101000101",
22011 => "0001000101000110",
22012 => "0001000101000111",
22013 => "0001000101001000",
22014 => "0001000101001001",
22015 => "0001000101001010",
22016 => "0001000101001011",
22017 => "0001000101001100",
22018 => "0001000101001101",
22019 => "0001000101001110",
22020 => "0001000101001111",
22021 => "0001000101010000",
22022 => "0001000101010001",
22023 => "0001000101010010",
22024 => "0001000101010011",
22025 => "0001000101010100",
22026 => "0001000101010101",
22027 => "0001000101010110",
22028 => "0001000101010111",
22029 => "0001000101011000",
22030 => "0001000101011001",
22031 => "0001000101011010",
22032 => "0001000101011011",
22033 => "0001000101011100",
22034 => "0001000101011101",
22035 => "0001000101011110",
22036 => "0001000101011111",
22037 => "0001000101100000",
22038 => "0001000101100001",
22039 => "0001000101100010",
22040 => "0001000101100011",
22041 => "0001000101100100",
22042 => "0001000101100101",
22043 => "0001000101100110",
22044 => "0001000101100111",
22045 => "0001000101101000",
22046 => "0001000101101001",
22047 => "0001000101101010",
22048 => "0001000101101011",
22049 => "0001000101101100",
22050 => "0001000101101101",
22051 => "0001000101101110",
22052 => "0001000101101111",
22053 => "0001000101110000",
22054 => "0001000101110001",
22055 => "0001000101110010",
22056 => "0001000101110011",
22057 => "0001000101110100",
22058 => "0001000101110101",
22059 => "0001000101110110",
22060 => "0001000101110111",
22061 => "0001000101111000",
22062 => "0001000101111001",
22063 => "0001000101111010",
22064 => "0001000101111011",
22065 => "0001000101111100",
22066 => "0001000101111101",
22067 => "0001000101111110",
22068 => "0001000101111111",
22069 => "0001000110000000",
22070 => "0001000110000001",
22071 => "0001000110000010",
22072 => "0001000110000011",
22073 => "0001000110000100",
22074 => "0001000110000101",
22075 => "0001000110000110",
22076 => "0001000110000111",
22077 => "0001000110001000",
22078 => "0001000110001001",
22079 => "0001000110001010",
22080 => "0001000110001100",
22081 => "0001000110001101",
22082 => "0001000110001110",
22083 => "0001000110001111",
22084 => "0001000110010000",
22085 => "0001000110010001",
22086 => "0001000110010010",
22087 => "0001000110010011",
22088 => "0001000110010100",
22089 => "0001000110010101",
22090 => "0001000110010110",
22091 => "0001000110010111",
22092 => "0001000110011000",
22093 => "0001000110011001",
22094 => "0001000110011010",
22095 => "0001000110011011",
22096 => "0001000110011100",
22097 => "0001000110011101",
22098 => "0001000110011110",
22099 => "0001000110011111",
22100 => "0001000110100000",
22101 => "0001000110100001",
22102 => "0001000110100010",
22103 => "0001000110100011",
22104 => "0001000110100100",
22105 => "0001000110100101",
22106 => "0001000110100110",
22107 => "0001000110100111",
22108 => "0001000110101000",
22109 => "0001000110101001",
22110 => "0001000110101010",
22111 => "0001000110101011",
22112 => "0001000110101100",
22113 => "0001000110101101",
22114 => "0001000110101110",
22115 => "0001000110101111",
22116 => "0001000110110000",
22117 => "0001000110110001",
22118 => "0001000110110010",
22119 => "0001000110110100",
22120 => "0001000110110101",
22121 => "0001000110110110",
22122 => "0001000110110111",
22123 => "0001000110111000",
22124 => "0001000110111001",
22125 => "0001000110111010",
22126 => "0001000110111011",
22127 => "0001000110111100",
22128 => "0001000110111101",
22129 => "0001000110111110",
22130 => "0001000110111111",
22131 => "0001000111000000",
22132 => "0001000111000001",
22133 => "0001000111000010",
22134 => "0001000111000011",
22135 => "0001000111000100",
22136 => "0001000111000101",
22137 => "0001000111000110",
22138 => "0001000111000111",
22139 => "0001000111001000",
22140 => "0001000111001001",
22141 => "0001000111001010",
22142 => "0001000111001011",
22143 => "0001000111001100",
22144 => "0001000111001101",
22145 => "0001000111001110",
22146 => "0001000111001111",
22147 => "0001000111010000",
22148 => "0001000111010001",
22149 => "0001000111010011",
22150 => "0001000111010100",
22151 => "0001000111010101",
22152 => "0001000111010110",
22153 => "0001000111010111",
22154 => "0001000111011000",
22155 => "0001000111011001",
22156 => "0001000111011010",
22157 => "0001000111011011",
22158 => "0001000111011100",
22159 => "0001000111011101",
22160 => "0001000111011110",
22161 => "0001000111011111",
22162 => "0001000111100000",
22163 => "0001000111100001",
22164 => "0001000111100010",
22165 => "0001000111100011",
22166 => "0001000111100100",
22167 => "0001000111100101",
22168 => "0001000111100110",
22169 => "0001000111100111",
22170 => "0001000111101000",
22171 => "0001000111101001",
22172 => "0001000111101010",
22173 => "0001000111101011",
22174 => "0001000111101100",
22175 => "0001000111101110",
22176 => "0001000111101111",
22177 => "0001000111110000",
22178 => "0001000111110001",
22179 => "0001000111110010",
22180 => "0001000111110011",
22181 => "0001000111110100",
22182 => "0001000111110101",
22183 => "0001000111110110",
22184 => "0001000111110111",
22185 => "0001000111111000",
22186 => "0001000111111001",
22187 => "0001000111111010",
22188 => "0001000111111011",
22189 => "0001000111111100",
22190 => "0001000111111101",
22191 => "0001000111111110",
22192 => "0001000111111111",
22193 => "0001001000000000",
22194 => "0001001000000001",
22195 => "0001001000000010",
22196 => "0001001000000011",
22197 => "0001001000000101",
22198 => "0001001000000110",
22199 => "0001001000000111",
22200 => "0001001000001000",
22201 => "0001001000001001",
22202 => "0001001000001010",
22203 => "0001001000001011",
22204 => "0001001000001100",
22205 => "0001001000001101",
22206 => "0001001000001110",
22207 => "0001001000001111",
22208 => "0001001000010000",
22209 => "0001001000010001",
22210 => "0001001000010010",
22211 => "0001001000010011",
22212 => "0001001000010100",
22213 => "0001001000010101",
22214 => "0001001000010110",
22215 => "0001001000010111",
22216 => "0001001000011000",
22217 => "0001001000011010",
22218 => "0001001000011011",
22219 => "0001001000011100",
22220 => "0001001000011101",
22221 => "0001001000011110",
22222 => "0001001000011111",
22223 => "0001001000100000",
22224 => "0001001000100001",
22225 => "0001001000100010",
22226 => "0001001000100011",
22227 => "0001001000100100",
22228 => "0001001000100101",
22229 => "0001001000100110",
22230 => "0001001000100111",
22231 => "0001001000101000",
22232 => "0001001000101001",
22233 => "0001001000101010",
22234 => "0001001000101011",
22235 => "0001001000101100",
22236 => "0001001000101110",
22237 => "0001001000101111",
22238 => "0001001000110000",
22239 => "0001001000110001",
22240 => "0001001000110010",
22241 => "0001001000110011",
22242 => "0001001000110100",
22243 => "0001001000110101",
22244 => "0001001000110110",
22245 => "0001001000110111",
22246 => "0001001000111000",
22247 => "0001001000111001",
22248 => "0001001000111010",
22249 => "0001001000111011",
22250 => "0001001000111100",
22251 => "0001001000111101",
22252 => "0001001000111110",
22253 => "0001001000111111",
22254 => "0001001001000001",
22255 => "0001001001000010",
22256 => "0001001001000011",
22257 => "0001001001000100",
22258 => "0001001001000101",
22259 => "0001001001000110",
22260 => "0001001001000111",
22261 => "0001001001001000",
22262 => "0001001001001001",
22263 => "0001001001001010",
22264 => "0001001001001011",
22265 => "0001001001001100",
22266 => "0001001001001101",
22267 => "0001001001001110",
22268 => "0001001001001111",
22269 => "0001001001010000",
22270 => "0001001001010010",
22271 => "0001001001010011",
22272 => "0001001001010100",
22273 => "0001001001010101",
22274 => "0001001001010110",
22275 => "0001001001010111",
22276 => "0001001001011000",
22277 => "0001001001011001",
22278 => "0001001001011010",
22279 => "0001001001011011",
22280 => "0001001001011100",
22281 => "0001001001011101",
22282 => "0001001001011110",
22283 => "0001001001011111",
22284 => "0001001001100000",
22285 => "0001001001100010",
22286 => "0001001001100011",
22287 => "0001001001100100",
22288 => "0001001001100101",
22289 => "0001001001100110",
22290 => "0001001001100111",
22291 => "0001001001101000",
22292 => "0001001001101001",
22293 => "0001001001101010",
22294 => "0001001001101011",
22295 => "0001001001101100",
22296 => "0001001001101101",
22297 => "0001001001101110",
22298 => "0001001001101111",
22299 => "0001001001110000",
22300 => "0001001001110010",
22301 => "0001001001110011",
22302 => "0001001001110100",
22303 => "0001001001110101",
22304 => "0001001001110110",
22305 => "0001001001110111",
22306 => "0001001001111000",
22307 => "0001001001111001",
22308 => "0001001001111010",
22309 => "0001001001111011",
22310 => "0001001001111100",
22311 => "0001001001111101",
22312 => "0001001001111110",
22313 => "0001001001111111",
22314 => "0001001010000001",
22315 => "0001001010000010",
22316 => "0001001010000011",
22317 => "0001001010000100",
22318 => "0001001010000101",
22319 => "0001001010000110",
22320 => "0001001010000111",
22321 => "0001001010001000",
22322 => "0001001010001001",
22323 => "0001001010001010",
22324 => "0001001010001011",
22325 => "0001001010001100",
22326 => "0001001010001101",
22327 => "0001001010001110",
22328 => "0001001010010000",
22329 => "0001001010010001",
22330 => "0001001010010010",
22331 => "0001001010010011",
22332 => "0001001010010100",
22333 => "0001001010010101",
22334 => "0001001010010110",
22335 => "0001001010010111",
22336 => "0001001010011000",
22337 => "0001001010011001",
22338 => "0001001010011010",
22339 => "0001001010011011",
22340 => "0001001010011100",
22341 => "0001001010011110",
22342 => "0001001010011111",
22343 => "0001001010100000",
22344 => "0001001010100001",
22345 => "0001001010100010",
22346 => "0001001010100011",
22347 => "0001001010100100",
22348 => "0001001010100101",
22349 => "0001001010100110",
22350 => "0001001010100111",
22351 => "0001001010101000",
22352 => "0001001010101001",
22353 => "0001001010101011",
22354 => "0001001010101100",
22355 => "0001001010101101",
22356 => "0001001010101110",
22357 => "0001001010101111",
22358 => "0001001010110000",
22359 => "0001001010110001",
22360 => "0001001010110010",
22361 => "0001001010110011",
22362 => "0001001010110100",
22363 => "0001001010110101",
22364 => "0001001010110110",
22365 => "0001001010111000",
22366 => "0001001010111001",
22367 => "0001001010111010",
22368 => "0001001010111011",
22369 => "0001001010111100",
22370 => "0001001010111101",
22371 => "0001001010111110",
22372 => "0001001010111111",
22373 => "0001001011000000",
22374 => "0001001011000001",
22375 => "0001001011000010",
22376 => "0001001011000011",
22377 => "0001001011000101",
22378 => "0001001011000110",
22379 => "0001001011000111",
22380 => "0001001011001000",
22381 => "0001001011001001",
22382 => "0001001011001010",
22383 => "0001001011001011",
22384 => "0001001011001100",
22385 => "0001001011001101",
22386 => "0001001011001110",
22387 => "0001001011001111",
22388 => "0001001011010001",
22389 => "0001001011010010",
22390 => "0001001011010011",
22391 => "0001001011010100",
22392 => "0001001011010101",
22393 => "0001001011010110",
22394 => "0001001011010111",
22395 => "0001001011011000",
22396 => "0001001011011001",
22397 => "0001001011011010",
22398 => "0001001011011011",
22399 => "0001001011011101",
22400 => "0001001011011110",
22401 => "0001001011011111",
22402 => "0001001011100000",
22403 => "0001001011100001",
22404 => "0001001011100010",
22405 => "0001001011100011",
22406 => "0001001011100100",
22407 => "0001001011100101",
22408 => "0001001011100110",
22409 => "0001001011100111",
22410 => "0001001011101001",
22411 => "0001001011101010",
22412 => "0001001011101011",
22413 => "0001001011101100",
22414 => "0001001011101101",
22415 => "0001001011101110",
22416 => "0001001011101111",
22417 => "0001001011110000",
22418 => "0001001011110001",
22419 => "0001001011110010",
22420 => "0001001011110100",
22421 => "0001001011110101",
22422 => "0001001011110110",
22423 => "0001001011110111",
22424 => "0001001011111000",
22425 => "0001001011111001",
22426 => "0001001011111010",
22427 => "0001001011111011",
22428 => "0001001011111100",
22429 => "0001001011111101",
22430 => "0001001011111111",
22431 => "0001001100000000",
22432 => "0001001100000001",
22433 => "0001001100000010",
22434 => "0001001100000011",
22435 => "0001001100000100",
22436 => "0001001100000101",
22437 => "0001001100000110",
22438 => "0001001100000111",
22439 => "0001001100001000",
22440 => "0001001100001010",
22441 => "0001001100001011",
22442 => "0001001100001100",
22443 => "0001001100001101",
22444 => "0001001100001110",
22445 => "0001001100001111",
22446 => "0001001100010000",
22447 => "0001001100010001",
22448 => "0001001100010010",
22449 => "0001001100010011",
22450 => "0001001100010101",
22451 => "0001001100010110",
22452 => "0001001100010111",
22453 => "0001001100011000",
22454 => "0001001100011001",
22455 => "0001001100011010",
22456 => "0001001100011011",
22457 => "0001001100011100",
22458 => "0001001100011101",
22459 => "0001001100011110",
22460 => "0001001100100000",
22461 => "0001001100100001",
22462 => "0001001100100010",
22463 => "0001001100100011",
22464 => "0001001100100100",
22465 => "0001001100100101",
22466 => "0001001100100110",
22467 => "0001001100100111",
22468 => "0001001100101000",
22469 => "0001001100101010",
22470 => "0001001100101011",
22471 => "0001001100101100",
22472 => "0001001100101101",
22473 => "0001001100101110",
22474 => "0001001100101111",
22475 => "0001001100110000",
22476 => "0001001100110001",
22477 => "0001001100110010",
22478 => "0001001100110100",
22479 => "0001001100110101",
22480 => "0001001100110110",
22481 => "0001001100110111",
22482 => "0001001100111000",
22483 => "0001001100111001",
22484 => "0001001100111010",
22485 => "0001001100111011",
22486 => "0001001100111100",
22487 => "0001001100111110",
22488 => "0001001100111111",
22489 => "0001001101000000",
22490 => "0001001101000001",
22491 => "0001001101000010",
22492 => "0001001101000011",
22493 => "0001001101000100",
22494 => "0001001101000101",
22495 => "0001001101000110",
22496 => "0001001101001000",
22497 => "0001001101001001",
22498 => "0001001101001010",
22499 => "0001001101001011",
22500 => "0001001101001100",
22501 => "0001001101001101",
22502 => "0001001101001110",
22503 => "0001001101001111",
22504 => "0001001101010000",
22505 => "0001001101010010",
22506 => "0001001101010011",
22507 => "0001001101010100",
22508 => "0001001101010101",
22509 => "0001001101010110",
22510 => "0001001101010111",
22511 => "0001001101011000",
22512 => "0001001101011001",
22513 => "0001001101011011",
22514 => "0001001101011100",
22515 => "0001001101011101",
22516 => "0001001101011110",
22517 => "0001001101011111",
22518 => "0001001101100000",
22519 => "0001001101100001",
22520 => "0001001101100010",
22521 => "0001001101100011",
22522 => "0001001101100101",
22523 => "0001001101100110",
22524 => "0001001101100111",
22525 => "0001001101101000",
22526 => "0001001101101001",
22527 => "0001001101101010",
22528 => "0001001101101011",
22529 => "0001001101101100",
22530 => "0001001101101110",
22531 => "0001001101101111",
22532 => "0001001101110000",
22533 => "0001001101110001",
22534 => "0001001101110010",
22535 => "0001001101110011",
22536 => "0001001101110100",
22537 => "0001001101110101",
22538 => "0001001101110111",
22539 => "0001001101111000",
22540 => "0001001101111001",
22541 => "0001001101111010",
22542 => "0001001101111011",
22543 => "0001001101111100",
22544 => "0001001101111101",
22545 => "0001001101111110",
22546 => "0001001110000000",
22547 => "0001001110000001",
22548 => "0001001110000010",
22549 => "0001001110000011",
22550 => "0001001110000100",
22551 => "0001001110000101",
22552 => "0001001110000110",
22553 => "0001001110000111",
22554 => "0001001110001001",
22555 => "0001001110001010",
22556 => "0001001110001011",
22557 => "0001001110001100",
22558 => "0001001110001101",
22559 => "0001001110001110",
22560 => "0001001110001111",
22561 => "0001001110010000",
22562 => "0001001110010010",
22563 => "0001001110010011",
22564 => "0001001110010100",
22565 => "0001001110010101",
22566 => "0001001110010110",
22567 => "0001001110010111",
22568 => "0001001110011000",
22569 => "0001001110011010",
22570 => "0001001110011011",
22571 => "0001001110011100",
22572 => "0001001110011101",
22573 => "0001001110011110",
22574 => "0001001110011111",
22575 => "0001001110100000",
22576 => "0001001110100001",
22577 => "0001001110100011",
22578 => "0001001110100100",
22579 => "0001001110100101",
22580 => "0001001110100110",
22581 => "0001001110100111",
22582 => "0001001110101000",
22583 => "0001001110101001",
22584 => "0001001110101011",
22585 => "0001001110101100",
22586 => "0001001110101101",
22587 => "0001001110101110",
22588 => "0001001110101111",
22589 => "0001001110110000",
22590 => "0001001110110001",
22591 => "0001001110110010",
22592 => "0001001110110100",
22593 => "0001001110110101",
22594 => "0001001110110110",
22595 => "0001001110110111",
22596 => "0001001110111000",
22597 => "0001001110111001",
22598 => "0001001110111010",
22599 => "0001001110111100",
22600 => "0001001110111101",
22601 => "0001001110111110",
22602 => "0001001110111111",
22603 => "0001001111000000",
22604 => "0001001111000001",
22605 => "0001001111000010",
22606 => "0001001111000100",
22607 => "0001001111000101",
22608 => "0001001111000110",
22609 => "0001001111000111",
22610 => "0001001111001000",
22611 => "0001001111001001",
22612 => "0001001111001010",
22613 => "0001001111001100",
22614 => "0001001111001101",
22615 => "0001001111001110",
22616 => "0001001111001111",
22617 => "0001001111010000",
22618 => "0001001111010001",
22619 => "0001001111010010",
22620 => "0001001111010100",
22621 => "0001001111010101",
22622 => "0001001111010110",
22623 => "0001001111010111",
22624 => "0001001111011000",
22625 => "0001001111011001",
22626 => "0001001111011010",
22627 => "0001001111011100",
22628 => "0001001111011101",
22629 => "0001001111011110",
22630 => "0001001111011111",
22631 => "0001001111100000",
22632 => "0001001111100001",
22633 => "0001001111100010",
22634 => "0001001111100100",
22635 => "0001001111100101",
22636 => "0001001111100110",
22637 => "0001001111100111",
22638 => "0001001111101000",
22639 => "0001001111101001",
22640 => "0001001111101010",
22641 => "0001001111101100",
22642 => "0001001111101101",
22643 => "0001001111101110",
22644 => "0001001111101111",
22645 => "0001001111110000",
22646 => "0001001111110001",
22647 => "0001001111110010",
22648 => "0001001111110100",
22649 => "0001001111110101",
22650 => "0001001111110110",
22651 => "0001001111110111",
22652 => "0001001111111000",
22653 => "0001001111111001",
22654 => "0001001111111011",
22655 => "0001001111111100",
22656 => "0001001111111101",
22657 => "0001001111111110",
22658 => "0001001111111111",
22659 => "0001010000000000",
22660 => "0001010000000001",
22661 => "0001010000000011",
22662 => "0001010000000100",
22663 => "0001010000000101",
22664 => "0001010000000110",
22665 => "0001010000000111",
22666 => "0001010000001000",
22667 => "0001010000001010",
22668 => "0001010000001011",
22669 => "0001010000001100",
22670 => "0001010000001101",
22671 => "0001010000001110",
22672 => "0001010000001111",
22673 => "0001010000010000",
22674 => "0001010000010010",
22675 => "0001010000010011",
22676 => "0001010000010100",
22677 => "0001010000010101",
22678 => "0001010000010110",
22679 => "0001010000010111",
22680 => "0001010000011001",
22681 => "0001010000011010",
22682 => "0001010000011011",
22683 => "0001010000011100",
22684 => "0001010000011101",
22685 => "0001010000011110",
22686 => "0001010000011111",
22687 => "0001010000100001",
22688 => "0001010000100010",
22689 => "0001010000100011",
22690 => "0001010000100100",
22691 => "0001010000100101",
22692 => "0001010000100110",
22693 => "0001010000101000",
22694 => "0001010000101001",
22695 => "0001010000101010",
22696 => "0001010000101011",
22697 => "0001010000101100",
22698 => "0001010000101101",
22699 => "0001010000101111",
22700 => "0001010000110000",
22701 => "0001010000110001",
22702 => "0001010000110010",
22703 => "0001010000110011",
22704 => "0001010000110100",
22705 => "0001010000110110",
22706 => "0001010000110111",
22707 => "0001010000111000",
22708 => "0001010000111001",
22709 => "0001010000111010",
22710 => "0001010000111011",
22711 => "0001010000111101",
22712 => "0001010000111110",
22713 => "0001010000111111",
22714 => "0001010001000000",
22715 => "0001010001000001",
22716 => "0001010001000010",
22717 => "0001010001000100",
22718 => "0001010001000101",
22719 => "0001010001000110",
22720 => "0001010001000111",
22721 => "0001010001001000",
22722 => "0001010001001001",
22723 => "0001010001001011",
22724 => "0001010001001100",
22725 => "0001010001001101",
22726 => "0001010001001110",
22727 => "0001010001001111",
22728 => "0001010001010000",
22729 => "0001010001010010",
22730 => "0001010001010011",
22731 => "0001010001010100",
22732 => "0001010001010101",
22733 => "0001010001010110",
22734 => "0001010001010111",
22735 => "0001010001011001",
22736 => "0001010001011010",
22737 => "0001010001011011",
22738 => "0001010001011100",
22739 => "0001010001011101",
22740 => "0001010001011110",
22741 => "0001010001100000",
22742 => "0001010001100001",
22743 => "0001010001100010",
22744 => "0001010001100011",
22745 => "0001010001100100",
22746 => "0001010001100101",
22747 => "0001010001100111",
22748 => "0001010001101000",
22749 => "0001010001101001",
22750 => "0001010001101010",
22751 => "0001010001101011",
22752 => "0001010001101101",
22753 => "0001010001101110",
22754 => "0001010001101111",
22755 => "0001010001110000",
22756 => "0001010001110001",
22757 => "0001010001110010",
22758 => "0001010001110100",
22759 => "0001010001110101",
22760 => "0001010001110110",
22761 => "0001010001110111",
22762 => "0001010001111000",
22763 => "0001010001111001",
22764 => "0001010001111011",
22765 => "0001010001111100",
22766 => "0001010001111101",
22767 => "0001010001111110",
22768 => "0001010001111111",
22769 => "0001010010000001",
22770 => "0001010010000010",
22771 => "0001010010000011",
22772 => "0001010010000100",
22773 => "0001010010000101",
22774 => "0001010010000110",
22775 => "0001010010001000",
22776 => "0001010010001001",
22777 => "0001010010001010",
22778 => "0001010010001011",
22779 => "0001010010001100",
22780 => "0001010010001101",
22781 => "0001010010001111",
22782 => "0001010010010000",
22783 => "0001010010010001",
22784 => "0001010010010010",
22785 => "0001010010010011",
22786 => "0001010010010101",
22787 => "0001010010010110",
22788 => "0001010010010111",
22789 => "0001010010011000",
22790 => "0001010010011001",
22791 => "0001010010011011",
22792 => "0001010010011100",
22793 => "0001010010011101",
22794 => "0001010010011110",
22795 => "0001010010011111",
22796 => "0001010010100000",
22797 => "0001010010100010",
22798 => "0001010010100011",
22799 => "0001010010100100",
22800 => "0001010010100101",
22801 => "0001010010100110",
22802 => "0001010010101000",
22803 => "0001010010101001",
22804 => "0001010010101010",
22805 => "0001010010101011",
22806 => "0001010010101100",
22807 => "0001010010101101",
22808 => "0001010010101111",
22809 => "0001010010110000",
22810 => "0001010010110001",
22811 => "0001010010110010",
22812 => "0001010010110011",
22813 => "0001010010110101",
22814 => "0001010010110110",
22815 => "0001010010110111",
22816 => "0001010010111000",
22817 => "0001010010111001",
22818 => "0001010010111011",
22819 => "0001010010111100",
22820 => "0001010010111101",
22821 => "0001010010111110",
22822 => "0001010010111111",
22823 => "0001010011000001",
22824 => "0001010011000010",
22825 => "0001010011000011",
22826 => "0001010011000100",
22827 => "0001010011000101",
22828 => "0001010011000110",
22829 => "0001010011001000",
22830 => "0001010011001001",
22831 => "0001010011001010",
22832 => "0001010011001011",
22833 => "0001010011001100",
22834 => "0001010011001110",
22835 => "0001010011001111",
22836 => "0001010011010000",
22837 => "0001010011010001",
22838 => "0001010011010010",
22839 => "0001010011010100",
22840 => "0001010011010101",
22841 => "0001010011010110",
22842 => "0001010011010111",
22843 => "0001010011011000",
22844 => "0001010011011010",
22845 => "0001010011011011",
22846 => "0001010011011100",
22847 => "0001010011011101",
22848 => "0001010011011110",
22849 => "0001010011100000",
22850 => "0001010011100001",
22851 => "0001010011100010",
22852 => "0001010011100011",
22853 => "0001010011100100",
22854 => "0001010011100110",
22855 => "0001010011100111",
22856 => "0001010011101000",
22857 => "0001010011101001",
22858 => "0001010011101010",
22859 => "0001010011101100",
22860 => "0001010011101101",
22861 => "0001010011101110",
22862 => "0001010011101111",
22863 => "0001010011110000",
22864 => "0001010011110010",
22865 => "0001010011110011",
22866 => "0001010011110100",
22867 => "0001010011110101",
22868 => "0001010011110110",
22869 => "0001010011111000",
22870 => "0001010011111001",
22871 => "0001010011111010",
22872 => "0001010011111011",
22873 => "0001010011111100",
22874 => "0001010011111110",
22875 => "0001010011111111",
22876 => "0001010100000000",
22877 => "0001010100000001",
22878 => "0001010100000010",
22879 => "0001010100000100",
22880 => "0001010100000101",
22881 => "0001010100000110",
22882 => "0001010100000111",
22883 => "0001010100001000",
22884 => "0001010100001010",
22885 => "0001010100001011",
22886 => "0001010100001100",
22887 => "0001010100001101",
22888 => "0001010100001111",
22889 => "0001010100010000",
22890 => "0001010100010001",
22891 => "0001010100010010",
22892 => "0001010100010011",
22893 => "0001010100010101",
22894 => "0001010100010110",
22895 => "0001010100010111",
22896 => "0001010100011000",
22897 => "0001010100011001",
22898 => "0001010100011011",
22899 => "0001010100011100",
22900 => "0001010100011101",
22901 => "0001010100011110",
22902 => "0001010100011111",
22903 => "0001010100100001",
22904 => "0001010100100010",
22905 => "0001010100100011",
22906 => "0001010100100100",
22907 => "0001010100100110",
22908 => "0001010100100111",
22909 => "0001010100101000",
22910 => "0001010100101001",
22911 => "0001010100101010",
22912 => "0001010100101100",
22913 => "0001010100101101",
22914 => "0001010100101110",
22915 => "0001010100101111",
22916 => "0001010100110000",
22917 => "0001010100110010",
22918 => "0001010100110011",
22919 => "0001010100110100",
22920 => "0001010100110101",
22921 => "0001010100110111",
22922 => "0001010100111000",
22923 => "0001010100111001",
22924 => "0001010100111010",
22925 => "0001010100111011",
22926 => "0001010100111101",
22927 => "0001010100111110",
22928 => "0001010100111111",
22929 => "0001010101000000",
22930 => "0001010101000001",
22931 => "0001010101000011",
22932 => "0001010101000100",
22933 => "0001010101000101",
22934 => "0001010101000110",
22935 => "0001010101001000",
22936 => "0001010101001001",
22937 => "0001010101001010",
22938 => "0001010101001011",
22939 => "0001010101001100",
22940 => "0001010101001110",
22941 => "0001010101001111",
22942 => "0001010101010000",
22943 => "0001010101010001",
22944 => "0001010101010011",
22945 => "0001010101010100",
22946 => "0001010101010101",
22947 => "0001010101010110",
22948 => "0001010101010111",
22949 => "0001010101011001",
22950 => "0001010101011010",
22951 => "0001010101011011",
22952 => "0001010101011100",
22953 => "0001010101011110",
22954 => "0001010101011111",
22955 => "0001010101100000",
22956 => "0001010101100001",
22957 => "0001010101100010",
22958 => "0001010101100100",
22959 => "0001010101100101",
22960 => "0001010101100110",
22961 => "0001010101100111",
22962 => "0001010101101001",
22963 => "0001010101101010",
22964 => "0001010101101011",
22965 => "0001010101101100",
22966 => "0001010101101101",
22967 => "0001010101101111",
22968 => "0001010101110000",
22969 => "0001010101110001",
22970 => "0001010101110010",
22971 => "0001010101110100",
22972 => "0001010101110101",
22973 => "0001010101110110",
22974 => "0001010101110111",
22975 => "0001010101111001",
22976 => "0001010101111010",
22977 => "0001010101111011",
22978 => "0001010101111100",
22979 => "0001010101111101",
22980 => "0001010101111111",
22981 => "0001010110000000",
22982 => "0001010110000001",
22983 => "0001010110000010",
22984 => "0001010110000100",
22985 => "0001010110000101",
22986 => "0001010110000110",
22987 => "0001010110000111",
22988 => "0001010110001001",
22989 => "0001010110001010",
22990 => "0001010110001011",
22991 => "0001010110001100",
22992 => "0001010110001101",
22993 => "0001010110001111",
22994 => "0001010110010000",
22995 => "0001010110010001",
22996 => "0001010110010010",
22997 => "0001010110010100",
22998 => "0001010110010101",
22999 => "0001010110010110",
23000 => "0001010110010111",
23001 => "0001010110011001",
23002 => "0001010110011010",
23003 => "0001010110011011",
23004 => "0001010110011100",
23005 => "0001010110011110",
23006 => "0001010110011111",
23007 => "0001010110100000",
23008 => "0001010110100001",
23009 => "0001010110100010",
23010 => "0001010110100100",
23011 => "0001010110100101",
23012 => "0001010110100110",
23013 => "0001010110100111",
23014 => "0001010110101001",
23015 => "0001010110101010",
23016 => "0001010110101011",
23017 => "0001010110101100",
23018 => "0001010110101110",
23019 => "0001010110101111",
23020 => "0001010110110000",
23021 => "0001010110110001",
23022 => "0001010110110011",
23023 => "0001010110110100",
23024 => "0001010110110101",
23025 => "0001010110110110",
23026 => "0001010110111000",
23027 => "0001010110111001",
23028 => "0001010110111010",
23029 => "0001010110111011",
23030 => "0001010110111101",
23031 => "0001010110111110",
23032 => "0001010110111111",
23033 => "0001010111000000",
23034 => "0001010111000010",
23035 => "0001010111000011",
23036 => "0001010111000100",
23037 => "0001010111000101",
23038 => "0001010111000110",
23039 => "0001010111001000",
23040 => "0001010111001001",
23041 => "0001010111001010",
23042 => "0001010111001011",
23043 => "0001010111001101",
23044 => "0001010111001110",
23045 => "0001010111001111",
23046 => "0001010111010000",
23047 => "0001010111010010",
23048 => "0001010111010011",
23049 => "0001010111010100",
23050 => "0001010111010101",
23051 => "0001010111010111",
23052 => "0001010111011000",
23053 => "0001010111011001",
23054 => "0001010111011010",
23055 => "0001010111011100",
23056 => "0001010111011101",
23057 => "0001010111011110",
23058 => "0001010111011111",
23059 => "0001010111100001",
23060 => "0001010111100010",
23061 => "0001010111100011",
23062 => "0001010111100100",
23063 => "0001010111100110",
23064 => "0001010111100111",
23065 => "0001010111101000",
23066 => "0001010111101001",
23067 => "0001010111101011",
23068 => "0001010111101100",
23069 => "0001010111101101",
23070 => "0001010111101110",
23071 => "0001010111110000",
23072 => "0001010111110001",
23073 => "0001010111110010",
23074 => "0001010111110011",
23075 => "0001010111110101",
23076 => "0001010111110110",
23077 => "0001010111110111",
23078 => "0001010111111001",
23079 => "0001010111111010",
23080 => "0001010111111011",
23081 => "0001010111111100",
23082 => "0001010111111110",
23083 => "0001010111111111",
23084 => "0001011000000000",
23085 => "0001011000000001",
23086 => "0001011000000011",
23087 => "0001011000000100",
23088 => "0001011000000101",
23089 => "0001011000000110",
23090 => "0001011000001000",
23091 => "0001011000001001",
23092 => "0001011000001010",
23093 => "0001011000001011",
23094 => "0001011000001101",
23095 => "0001011000001110",
23096 => "0001011000001111",
23097 => "0001011000010000",
23098 => "0001011000010010",
23099 => "0001011000010011",
23100 => "0001011000010100",
23101 => "0001011000010101",
23102 => "0001011000010111",
23103 => "0001011000011000",
23104 => "0001011000011001",
23105 => "0001011000011011",
23106 => "0001011000011100",
23107 => "0001011000011101",
23108 => "0001011000011110",
23109 => "0001011000100000",
23110 => "0001011000100001",
23111 => "0001011000100010",
23112 => "0001011000100011",
23113 => "0001011000100101",
23114 => "0001011000100110",
23115 => "0001011000100111",
23116 => "0001011000101000",
23117 => "0001011000101010",
23118 => "0001011000101011",
23119 => "0001011000101100",
23120 => "0001011000101101",
23121 => "0001011000101111",
23122 => "0001011000110000",
23123 => "0001011000110001",
23124 => "0001011000110011",
23125 => "0001011000110100",
23126 => "0001011000110101",
23127 => "0001011000110110",
23128 => "0001011000111000",
23129 => "0001011000111001",
23130 => "0001011000111010",
23131 => "0001011000111011",
23132 => "0001011000111101",
23133 => "0001011000111110",
23134 => "0001011000111111",
23135 => "0001011001000000",
23136 => "0001011001000010",
23137 => "0001011001000011",
23138 => "0001011001000100",
23139 => "0001011001000110",
23140 => "0001011001000111",
23141 => "0001011001001000",
23142 => "0001011001001001",
23143 => "0001011001001011",
23144 => "0001011001001100",
23145 => "0001011001001101",
23146 => "0001011001001110",
23147 => "0001011001010000",
23148 => "0001011001010001",
23149 => "0001011001010010",
23150 => "0001011001010100",
23151 => "0001011001010101",
23152 => "0001011001010110",
23153 => "0001011001010111",
23154 => "0001011001011001",
23155 => "0001011001011010",
23156 => "0001011001011011",
23157 => "0001011001011100",
23158 => "0001011001011110",
23159 => "0001011001011111",
23160 => "0001011001100000",
23161 => "0001011001100010",
23162 => "0001011001100011",
23163 => "0001011001100100",
23164 => "0001011001100101",
23165 => "0001011001100111",
23166 => "0001011001101000",
23167 => "0001011001101001",
23168 => "0001011001101011",
23169 => "0001011001101100",
23170 => "0001011001101101",
23171 => "0001011001101110",
23172 => "0001011001110000",
23173 => "0001011001110001",
23174 => "0001011001110010",
23175 => "0001011001110011",
23176 => "0001011001110101",
23177 => "0001011001110110",
23178 => "0001011001110111",
23179 => "0001011001111001",
23180 => "0001011001111010",
23181 => "0001011001111011",
23182 => "0001011001111100",
23183 => "0001011001111110",
23184 => "0001011001111111",
23185 => "0001011010000000",
23186 => "0001011010000010",
23187 => "0001011010000011",
23188 => "0001011010000100",
23189 => "0001011010000101",
23190 => "0001011010000111",
23191 => "0001011010001000",
23192 => "0001011010001001",
23193 => "0001011010001011",
23194 => "0001011010001100",
23195 => "0001011010001101",
23196 => "0001011010001110",
23197 => "0001011010010000",
23198 => "0001011010010001",
23199 => "0001011010010010",
23200 => "0001011010010100",
23201 => "0001011010010101",
23202 => "0001011010010110",
23203 => "0001011010010111",
23204 => "0001011010011001",
23205 => "0001011010011010",
23206 => "0001011010011011",
23207 => "0001011010011101",
23208 => "0001011010011110",
23209 => "0001011010011111",
23210 => "0001011010100000",
23211 => "0001011010100010",
23212 => "0001011010100011",
23213 => "0001011010100100",
23214 => "0001011010100110",
23215 => "0001011010100111",
23216 => "0001011010101000",
23217 => "0001011010101001",
23218 => "0001011010101011",
23219 => "0001011010101100",
23220 => "0001011010101101",
23221 => "0001011010101111",
23222 => "0001011010110000",
23223 => "0001011010110001",
23224 => "0001011010110011",
23225 => "0001011010110100",
23226 => "0001011010110101",
23227 => "0001011010110110",
23228 => "0001011010111000",
23229 => "0001011010111001",
23230 => "0001011010111010",
23231 => "0001011010111100",
23232 => "0001011010111101",
23233 => "0001011010111110",
23234 => "0001011010111111",
23235 => "0001011011000001",
23236 => "0001011011000010",
23237 => "0001011011000011",
23238 => "0001011011000101",
23239 => "0001011011000110",
23240 => "0001011011000111",
23241 => "0001011011001001",
23242 => "0001011011001010",
23243 => "0001011011001011",
23244 => "0001011011001100",
23245 => "0001011011001110",
23246 => "0001011011001111",
23247 => "0001011011010000",
23248 => "0001011011010010",
23249 => "0001011011010011",
23250 => "0001011011010100",
23251 => "0001011011010110",
23252 => "0001011011010111",
23253 => "0001011011011000",
23254 => "0001011011011001",
23255 => "0001011011011011",
23256 => "0001011011011100",
23257 => "0001011011011101",
23258 => "0001011011011111",
23259 => "0001011011100000",
23260 => "0001011011100001",
23261 => "0001011011100011",
23262 => "0001011011100100",
23263 => "0001011011100101",
23264 => "0001011011100110",
23265 => "0001011011101000",
23266 => "0001011011101001",
23267 => "0001011011101010",
23268 => "0001011011101100",
23269 => "0001011011101101",
23270 => "0001011011101110",
23271 => "0001011011110000",
23272 => "0001011011110001",
23273 => "0001011011110010",
23274 => "0001011011110100",
23275 => "0001011011110101",
23276 => "0001011011110110",
23277 => "0001011011110111",
23278 => "0001011011111001",
23279 => "0001011011111010",
23280 => "0001011011111011",
23281 => "0001011011111101",
23282 => "0001011011111110",
23283 => "0001011011111111",
23284 => "0001011100000001",
23285 => "0001011100000010",
23286 => "0001011100000011",
23287 => "0001011100000101",
23288 => "0001011100000110",
23289 => "0001011100000111",
23290 => "0001011100001000",
23291 => "0001011100001010",
23292 => "0001011100001011",
23293 => "0001011100001100",
23294 => "0001011100001110",
23295 => "0001011100001111",
23296 => "0001011100010000",
23297 => "0001011100010010",
23298 => "0001011100010011",
23299 => "0001011100010100",
23300 => "0001011100010110",
23301 => "0001011100010111",
23302 => "0001011100011000",
23303 => "0001011100011001",
23304 => "0001011100011011",
23305 => "0001011100011100",
23306 => "0001011100011101",
23307 => "0001011100011111",
23308 => "0001011100100000",
23309 => "0001011100100001",
23310 => "0001011100100011",
23311 => "0001011100100100",
23312 => "0001011100100101",
23313 => "0001011100100111",
23314 => "0001011100101000",
23315 => "0001011100101001",
23316 => "0001011100101011",
23317 => "0001011100101100",
23318 => "0001011100101101",
23319 => "0001011100101111",
23320 => "0001011100110000",
23321 => "0001011100110001",
23322 => "0001011100110010",
23323 => "0001011100110100",
23324 => "0001011100110101",
23325 => "0001011100110110",
23326 => "0001011100111000",
23327 => "0001011100111001",
23328 => "0001011100111010",
23329 => "0001011100111100",
23330 => "0001011100111101",
23331 => "0001011100111110",
23332 => "0001011101000000",
23333 => "0001011101000001",
23334 => "0001011101000010",
23335 => "0001011101000100",
23336 => "0001011101000101",
23337 => "0001011101000110",
23338 => "0001011101001000",
23339 => "0001011101001001",
23340 => "0001011101001010",
23341 => "0001011101001100",
23342 => "0001011101001101",
23343 => "0001011101001110",
23344 => "0001011101010000",
23345 => "0001011101010001",
23346 => "0001011101010010",
23347 => "0001011101010100",
23348 => "0001011101010101",
23349 => "0001011101010110",
23350 => "0001011101011000",
23351 => "0001011101011001",
23352 => "0001011101011010",
23353 => "0001011101011011",
23354 => "0001011101011101",
23355 => "0001011101011110",
23356 => "0001011101011111",
23357 => "0001011101100001",
23358 => "0001011101100010",
23359 => "0001011101100011",
23360 => "0001011101100101",
23361 => "0001011101100110",
23362 => "0001011101100111",
23363 => "0001011101101001",
23364 => "0001011101101010",
23365 => "0001011101101011",
23366 => "0001011101101101",
23367 => "0001011101101110",
23368 => "0001011101101111",
23369 => "0001011101110001",
23370 => "0001011101110010",
23371 => "0001011101110011",
23372 => "0001011101110101",
23373 => "0001011101110110",
23374 => "0001011101110111",
23375 => "0001011101111001",
23376 => "0001011101111010",
23377 => "0001011101111011",
23378 => "0001011101111101",
23379 => "0001011101111110",
23380 => "0001011101111111",
23381 => "0001011110000001",
23382 => "0001011110000010",
23383 => "0001011110000011",
23384 => "0001011110000101",
23385 => "0001011110000110",
23386 => "0001011110000111",
23387 => "0001011110001001",
23388 => "0001011110001010",
23389 => "0001011110001011",
23390 => "0001011110001101",
23391 => "0001011110001110",
23392 => "0001011110001111",
23393 => "0001011110010001",
23394 => "0001011110010010",
23395 => "0001011110010011",
23396 => "0001011110010101",
23397 => "0001011110010110",
23398 => "0001011110010111",
23399 => "0001011110011001",
23400 => "0001011110011010",
23401 => "0001011110011011",
23402 => "0001011110011101",
23403 => "0001011110011110",
23404 => "0001011110100000",
23405 => "0001011110100001",
23406 => "0001011110100010",
23407 => "0001011110100100",
23408 => "0001011110100101",
23409 => "0001011110100110",
23410 => "0001011110101000",
23411 => "0001011110101001",
23412 => "0001011110101010",
23413 => "0001011110101100",
23414 => "0001011110101101",
23415 => "0001011110101110",
23416 => "0001011110110000",
23417 => "0001011110110001",
23418 => "0001011110110010",
23419 => "0001011110110100",
23420 => "0001011110110101",
23421 => "0001011110110110",
23422 => "0001011110111000",
23423 => "0001011110111001",
23424 => "0001011110111010",
23425 => "0001011110111100",
23426 => "0001011110111101",
23427 => "0001011110111110",
23428 => "0001011111000000",
23429 => "0001011111000001",
23430 => "0001011111000010",
23431 => "0001011111000100",
23432 => "0001011111000101",
23433 => "0001011111000110",
23434 => "0001011111001000",
23435 => "0001011111001001",
23436 => "0001011111001011",
23437 => "0001011111001100",
23438 => "0001011111001101",
23439 => "0001011111001111",
23440 => "0001011111010000",
23441 => "0001011111010001",
23442 => "0001011111010011",
23443 => "0001011111010100",
23444 => "0001011111010101",
23445 => "0001011111010111",
23446 => "0001011111011000",
23447 => "0001011111011001",
23448 => "0001011111011011",
23449 => "0001011111011100",
23450 => "0001011111011101",
23451 => "0001011111011111",
23452 => "0001011111100000",
23453 => "0001011111100010",
23454 => "0001011111100011",
23455 => "0001011111100100",
23456 => "0001011111100110",
23457 => "0001011111100111",
23458 => "0001011111101000",
23459 => "0001011111101010",
23460 => "0001011111101011",
23461 => "0001011111101100",
23462 => "0001011111101110",
23463 => "0001011111101111",
23464 => "0001011111110000",
23465 => "0001011111110010",
23466 => "0001011111110011",
23467 => "0001011111110100",
23468 => "0001011111110110",
23469 => "0001011111110111",
23470 => "0001011111111001",
23471 => "0001011111111010",
23472 => "0001011111111011",
23473 => "0001011111111101",
23474 => "0001011111111110",
23475 => "0001011111111111",
23476 => "0001100000000001",
23477 => "0001100000000010",
23478 => "0001100000000011",
23479 => "0001100000000101",
23480 => "0001100000000110",
23481 => "0001100000001000",
23482 => "0001100000001001",
23483 => "0001100000001010",
23484 => "0001100000001100",
23485 => "0001100000001101",
23486 => "0001100000001110",
23487 => "0001100000010000",
23488 => "0001100000010001",
23489 => "0001100000010010",
23490 => "0001100000010100",
23491 => "0001100000010101",
23492 => "0001100000010110",
23493 => "0001100000011000",
23494 => "0001100000011001",
23495 => "0001100000011011",
23496 => "0001100000011100",
23497 => "0001100000011101",
23498 => "0001100000011111",
23499 => "0001100000100000",
23500 => "0001100000100001",
23501 => "0001100000100011",
23502 => "0001100000100100",
23503 => "0001100000100110",
23504 => "0001100000100111",
23505 => "0001100000101000",
23506 => "0001100000101010",
23507 => "0001100000101011",
23508 => "0001100000101100",
23509 => "0001100000101110",
23510 => "0001100000101111",
23511 => "0001100000110000",
23512 => "0001100000110010",
23513 => "0001100000110011",
23514 => "0001100000110101",
23515 => "0001100000110110",
23516 => "0001100000110111",
23517 => "0001100000111001",
23518 => "0001100000111010",
23519 => "0001100000111011",
23520 => "0001100000111101",
23521 => "0001100000111110",
23522 => "0001100001000000",
23523 => "0001100001000001",
23524 => "0001100001000010",
23525 => "0001100001000100",
23526 => "0001100001000101",
23527 => "0001100001000110",
23528 => "0001100001001000",
23529 => "0001100001001001",
23530 => "0001100001001011",
23531 => "0001100001001100",
23532 => "0001100001001101",
23533 => "0001100001001111",
23534 => "0001100001010000",
23535 => "0001100001010001",
23536 => "0001100001010011",
23537 => "0001100001010100",
23538 => "0001100001010110",
23539 => "0001100001010111",
23540 => "0001100001011000",
23541 => "0001100001011010",
23542 => "0001100001011011",
23543 => "0001100001011100",
23544 => "0001100001011110",
23545 => "0001100001011111",
23546 => "0001100001100001",
23547 => "0001100001100010",
23548 => "0001100001100011",
23549 => "0001100001100101",
23550 => "0001100001100110",
23551 => "0001100001100111",
23552 => "0001100001101001",
23553 => "0001100001101010",
23554 => "0001100001101100",
23555 => "0001100001101101",
23556 => "0001100001101110",
23557 => "0001100001110000",
23558 => "0001100001110001",
23559 => "0001100001110010",
23560 => "0001100001110100",
23561 => "0001100001110101",
23562 => "0001100001110111",
23563 => "0001100001111000",
23564 => "0001100001111001",
23565 => "0001100001111011",
23566 => "0001100001111100",
23567 => "0001100001111110",
23568 => "0001100001111111",
23569 => "0001100010000000",
23570 => "0001100010000010",
23571 => "0001100010000011",
23572 => "0001100010000100",
23573 => "0001100010000110",
23574 => "0001100010000111",
23575 => "0001100010001001",
23576 => "0001100010001010",
23577 => "0001100010001011",
23578 => "0001100010001101",
23579 => "0001100010001110",
23580 => "0001100010010000",
23581 => "0001100010010001",
23582 => "0001100010010010",
23583 => "0001100010010100",
23584 => "0001100010010101",
23585 => "0001100010010111",
23586 => "0001100010011000",
23587 => "0001100010011001",
23588 => "0001100010011011",
23589 => "0001100010011100",
23590 => "0001100010011101",
23591 => "0001100010011111",
23592 => "0001100010100000",
23593 => "0001100010100010",
23594 => "0001100010100011",
23595 => "0001100010100100",
23596 => "0001100010100110",
23597 => "0001100010100111",
23598 => "0001100010101001",
23599 => "0001100010101010",
23600 => "0001100010101011",
23601 => "0001100010101101",
23602 => "0001100010101110",
23603 => "0001100010110000",
23604 => "0001100010110001",
23605 => "0001100010110010",
23606 => "0001100010110100",
23607 => "0001100010110101",
23608 => "0001100010110111",
23609 => "0001100010111000",
23610 => "0001100010111001",
23611 => "0001100010111011",
23612 => "0001100010111100",
23613 => "0001100010111110",
23614 => "0001100010111111",
23615 => "0001100011000000",
23616 => "0001100011000010",
23617 => "0001100011000011",
23618 => "0001100011000101",
23619 => "0001100011000110",
23620 => "0001100011000111",
23621 => "0001100011001001",
23622 => "0001100011001010",
23623 => "0001100011001100",
23624 => "0001100011001101",
23625 => "0001100011001110",
23626 => "0001100011010000",
23627 => "0001100011010001",
23628 => "0001100011010011",
23629 => "0001100011010100",
23630 => "0001100011010101",
23631 => "0001100011010111",
23632 => "0001100011011000",
23633 => "0001100011011010",
23634 => "0001100011011011",
23635 => "0001100011011100",
23636 => "0001100011011110",
23637 => "0001100011011111",
23638 => "0001100011100001",
23639 => "0001100011100010",
23640 => "0001100011100011",
23641 => "0001100011100101",
23642 => "0001100011100110",
23643 => "0001100011101000",
23644 => "0001100011101001",
23645 => "0001100011101010",
23646 => "0001100011101100",
23647 => "0001100011101101",
23648 => "0001100011101111",
23649 => "0001100011110000",
23650 => "0001100011110001",
23651 => "0001100011110011",
23652 => "0001100011110100",
23653 => "0001100011110110",
23654 => "0001100011110111",
23655 => "0001100011111000",
23656 => "0001100011111010",
23657 => "0001100011111011",
23658 => "0001100011111101",
23659 => "0001100011111110",
23660 => "0001100011111111",
23661 => "0001100100000001",
23662 => "0001100100000010",
23663 => "0001100100000100",
23664 => "0001100100000101",
23665 => "0001100100000111",
23666 => "0001100100001000",
23667 => "0001100100001001",
23668 => "0001100100001011",
23669 => "0001100100001100",
23670 => "0001100100001110",
23671 => "0001100100001111",
23672 => "0001100100010000",
23673 => "0001100100010010",
23674 => "0001100100010011",
23675 => "0001100100010101",
23676 => "0001100100010110",
23677 => "0001100100010111",
23678 => "0001100100011001",
23679 => "0001100100011010",
23680 => "0001100100011100",
23681 => "0001100100011101",
23682 => "0001100100011111",
23683 => "0001100100100000",
23684 => "0001100100100001",
23685 => "0001100100100011",
23686 => "0001100100100100",
23687 => "0001100100100110",
23688 => "0001100100100111",
23689 => "0001100100101000",
23690 => "0001100100101010",
23691 => "0001100100101011",
23692 => "0001100100101101",
23693 => "0001100100101110",
23694 => "0001100100110000",
23695 => "0001100100110001",
23696 => "0001100100110010",
23697 => "0001100100110100",
23698 => "0001100100110101",
23699 => "0001100100110111",
23700 => "0001100100111000",
23701 => "0001100100111010",
23702 => "0001100100111011",
23703 => "0001100100111100",
23704 => "0001100100111110",
23705 => "0001100100111111",
23706 => "0001100101000001",
23707 => "0001100101000010",
23708 => "0001100101000011",
23709 => "0001100101000101",
23710 => "0001100101000110",
23711 => "0001100101001000",
23712 => "0001100101001001",
23713 => "0001100101001011",
23714 => "0001100101001100",
23715 => "0001100101001101",
23716 => "0001100101001111",
23717 => "0001100101010000",
23718 => "0001100101010010",
23719 => "0001100101010011",
23720 => "0001100101010101",
23721 => "0001100101010110",
23722 => "0001100101010111",
23723 => "0001100101011001",
23724 => "0001100101011010",
23725 => "0001100101011100",
23726 => "0001100101011101",
23727 => "0001100101011111",
23728 => "0001100101100000",
23729 => "0001100101100001",
23730 => "0001100101100011",
23731 => "0001100101100100",
23732 => "0001100101100110",
23733 => "0001100101100111",
23734 => "0001100101101001",
23735 => "0001100101101010",
23736 => "0001100101101011",
23737 => "0001100101101101",
23738 => "0001100101101110",
23739 => "0001100101110000",
23740 => "0001100101110001",
23741 => "0001100101110011",
23742 => "0001100101110100",
23743 => "0001100101110101",
23744 => "0001100101110111",
23745 => "0001100101111000",
23746 => "0001100101111010",
23747 => "0001100101111011",
23748 => "0001100101111101",
23749 => "0001100101111110",
23750 => "0001100110000000",
23751 => "0001100110000001",
23752 => "0001100110000010",
23753 => "0001100110000100",
23754 => "0001100110000101",
23755 => "0001100110000111",
23756 => "0001100110001000",
23757 => "0001100110001010",
23758 => "0001100110001011",
23759 => "0001100110001100",
23760 => "0001100110001110",
23761 => "0001100110001111",
23762 => "0001100110010001",
23763 => "0001100110010010",
23764 => "0001100110010100",
23765 => "0001100110010101",
23766 => "0001100110010111",
23767 => "0001100110011000",
23768 => "0001100110011001",
23769 => "0001100110011011",
23770 => "0001100110011100",
23771 => "0001100110011110",
23772 => "0001100110011111",
23773 => "0001100110100001",
23774 => "0001100110100010",
23775 => "0001100110100011",
23776 => "0001100110100101",
23777 => "0001100110100110",
23778 => "0001100110101000",
23779 => "0001100110101001",
23780 => "0001100110101011",
23781 => "0001100110101100",
23782 => "0001100110101110",
23783 => "0001100110101111",
23784 => "0001100110110000",
23785 => "0001100110110010",
23786 => "0001100110110011",
23787 => "0001100110110101",
23788 => "0001100110110110",
23789 => "0001100110111000",
23790 => "0001100110111001",
23791 => "0001100110111011",
23792 => "0001100110111100",
23793 => "0001100110111101",
23794 => "0001100110111111",
23795 => "0001100111000000",
23796 => "0001100111000010",
23797 => "0001100111000011",
23798 => "0001100111000101",
23799 => "0001100111000110",
23800 => "0001100111001000",
23801 => "0001100111001001",
23802 => "0001100111001011",
23803 => "0001100111001100",
23804 => "0001100111001101",
23805 => "0001100111001111",
23806 => "0001100111010000",
23807 => "0001100111010010",
23808 => "0001100111010011",
23809 => "0001100111010101",
23810 => "0001100111010110",
23811 => "0001100111011000",
23812 => "0001100111011001",
23813 => "0001100111011010",
23814 => "0001100111011100",
23815 => "0001100111011101",
23816 => "0001100111011111",
23817 => "0001100111100000",
23818 => "0001100111100010",
23819 => "0001100111100011",
23820 => "0001100111100101",
23821 => "0001100111100110",
23822 => "0001100111101000",
23823 => "0001100111101001",
23824 => "0001100111101010",
23825 => "0001100111101100",
23826 => "0001100111101101",
23827 => "0001100111101111",
23828 => "0001100111110000",
23829 => "0001100111110010",
23830 => "0001100111110011",
23831 => "0001100111110101",
23832 => "0001100111110110",
23833 => "0001100111111000",
23834 => "0001100111111001",
23835 => "0001100111111010",
23836 => "0001100111111100",
23837 => "0001100111111101",
23838 => "0001100111111111",
23839 => "0001101000000000",
23840 => "0001101000000010",
23841 => "0001101000000011",
23842 => "0001101000000101",
23843 => "0001101000000110",
23844 => "0001101000001000",
23845 => "0001101000001001",
23846 => "0001101000001011",
23847 => "0001101000001100",
23848 => "0001101000001101",
23849 => "0001101000001111",
23850 => "0001101000010000",
23851 => "0001101000010010",
23852 => "0001101000010011",
23853 => "0001101000010101",
23854 => "0001101000010110",
23855 => "0001101000011000",
23856 => "0001101000011001",
23857 => "0001101000011011",
23858 => "0001101000011100",
23859 => "0001101000011110",
23860 => "0001101000011111",
23861 => "0001101000100001",
23862 => "0001101000100010",
23863 => "0001101000100011",
23864 => "0001101000100101",
23865 => "0001101000100110",
23866 => "0001101000101000",
23867 => "0001101000101001",
23868 => "0001101000101011",
23869 => "0001101000101100",
23870 => "0001101000101110",
23871 => "0001101000101111",
23872 => "0001101000110001",
23873 => "0001101000110010",
23874 => "0001101000110100",
23875 => "0001101000110101",
23876 => "0001101000110111",
23877 => "0001101000111000",
23878 => "0001101000111001",
23879 => "0001101000111011",
23880 => "0001101000111100",
23881 => "0001101000111110",
23882 => "0001101000111111",
23883 => "0001101001000001",
23884 => "0001101001000010",
23885 => "0001101001000100",
23886 => "0001101001000101",
23887 => "0001101001000111",
23888 => "0001101001001000",
23889 => "0001101001001010",
23890 => "0001101001001011",
23891 => "0001101001001101",
23892 => "0001101001001110",
23893 => "0001101001010000",
23894 => "0001101001010001",
23895 => "0001101001010011",
23896 => "0001101001010100",
23897 => "0001101001010110",
23898 => "0001101001010111",
23899 => "0001101001011000",
23900 => "0001101001011010",
23901 => "0001101001011011",
23902 => "0001101001011101",
23903 => "0001101001011110",
23904 => "0001101001100000",
23905 => "0001101001100001",
23906 => "0001101001100011",
23907 => "0001101001100100",
23908 => "0001101001100110",
23909 => "0001101001100111",
23910 => "0001101001101001",
23911 => "0001101001101010",
23912 => "0001101001101100",
23913 => "0001101001101101",
23914 => "0001101001101111",
23915 => "0001101001110000",
23916 => "0001101001110010",
23917 => "0001101001110011",
23918 => "0001101001110101",
23919 => "0001101001110110",
23920 => "0001101001111000",
23921 => "0001101001111001",
23922 => "0001101001111011",
23923 => "0001101001111100",
23924 => "0001101001111101",
23925 => "0001101001111111",
23926 => "0001101010000000",
23927 => "0001101010000010",
23928 => "0001101010000011",
23929 => "0001101010000101",
23930 => "0001101010000110",
23931 => "0001101010001000",
23932 => "0001101010001001",
23933 => "0001101010001011",
23934 => "0001101010001100",
23935 => "0001101010001110",
23936 => "0001101010001111",
23937 => "0001101010010001",
23938 => "0001101010010010",
23939 => "0001101010010100",
23940 => "0001101010010101",
23941 => "0001101010010111",
23942 => "0001101010011000",
23943 => "0001101010011010",
23944 => "0001101010011011",
23945 => "0001101010011101",
23946 => "0001101010011110",
23947 => "0001101010100000",
23948 => "0001101010100001",
23949 => "0001101010100011",
23950 => "0001101010100100",
23951 => "0001101010100110",
23952 => "0001101010100111",
23953 => "0001101010101001",
23954 => "0001101010101010",
23955 => "0001101010101100",
23956 => "0001101010101101",
23957 => "0001101010101111",
23958 => "0001101010110000",
23959 => "0001101010110010",
23960 => "0001101010110011",
23961 => "0001101010110101",
23962 => "0001101010110110",
23963 => "0001101010111000",
23964 => "0001101010111001",
23965 => "0001101010111011",
23966 => "0001101010111100",
23967 => "0001101010111110",
23968 => "0001101010111111",
23969 => "0001101011000001",
23970 => "0001101011000010",
23971 => "0001101011000100",
23972 => "0001101011000101",
23973 => "0001101011000111",
23974 => "0001101011001000",
23975 => "0001101011001010",
23976 => "0001101011001011",
23977 => "0001101011001101",
23978 => "0001101011001110",
23979 => "0001101011010000",
23980 => "0001101011010001",
23981 => "0001101011010011",
23982 => "0001101011010100",
23983 => "0001101011010110",
23984 => "0001101011010111",
23985 => "0001101011011001",
23986 => "0001101011011010",
23987 => "0001101011011100",
23988 => "0001101011011101",
23989 => "0001101011011111",
23990 => "0001101011100000",
23991 => "0001101011100010",
23992 => "0001101011100011",
23993 => "0001101011100101",
23994 => "0001101011100110",
23995 => "0001101011101000",
23996 => "0001101011101001",
23997 => "0001101011101011",
23998 => "0001101011101100",
23999 => "0001101011101110",
24000 => "0001101011101111",
24001 => "0001101011110001",
24002 => "0001101011110010",
24003 => "0001101011110100",
24004 => "0001101011110101",
24005 => "0001101011110111",
24006 => "0001101011111000",
24007 => "0001101011111010",
24008 => "0001101011111011",
24009 => "0001101011111101",
24010 => "0001101011111110",
24011 => "0001101100000000",
24012 => "0001101100000001",
24013 => "0001101100000011",
24014 => "0001101100000100",
24015 => "0001101100000110",
24016 => "0001101100000111",
24017 => "0001101100001001",
24018 => "0001101100001010",
24019 => "0001101100001100",
24020 => "0001101100001101",
24021 => "0001101100001111",
24022 => "0001101100010000",
24023 => "0001101100010010",
24024 => "0001101100010011",
24025 => "0001101100010101",
24026 => "0001101100010110",
24027 => "0001101100011000",
24028 => "0001101100011001",
24029 => "0001101100011011",
24030 => "0001101100011100",
24031 => "0001101100011110",
24032 => "0001101100011111",
24033 => "0001101100100001",
24034 => "0001101100100011",
24035 => "0001101100100100",
24036 => "0001101100100110",
24037 => "0001101100100111",
24038 => "0001101100101001",
24039 => "0001101100101010",
24040 => "0001101100101100",
24041 => "0001101100101101",
24042 => "0001101100101111",
24043 => "0001101100110000",
24044 => "0001101100110010",
24045 => "0001101100110011",
24046 => "0001101100110101",
24047 => "0001101100110110",
24048 => "0001101100111000",
24049 => "0001101100111001",
24050 => "0001101100111011",
24051 => "0001101100111100",
24052 => "0001101100111110",
24053 => "0001101100111111",
24054 => "0001101101000001",
24055 => "0001101101000010",
24056 => "0001101101000100",
24057 => "0001101101000101",
24058 => "0001101101000111",
24059 => "0001101101001001",
24060 => "0001101101001010",
24061 => "0001101101001100",
24062 => "0001101101001101",
24063 => "0001101101001111",
24064 => "0001101101010000",
24065 => "0001101101010010",
24066 => "0001101101010011",
24067 => "0001101101010101",
24068 => "0001101101010110",
24069 => "0001101101011000",
24070 => "0001101101011001",
24071 => "0001101101011011",
24072 => "0001101101011100",
24073 => "0001101101011110",
24074 => "0001101101011111",
24075 => "0001101101100001",
24076 => "0001101101100010",
24077 => "0001101101100100",
24078 => "0001101101100110",
24079 => "0001101101100111",
24080 => "0001101101101001",
24081 => "0001101101101010",
24082 => "0001101101101100",
24083 => "0001101101101101",
24084 => "0001101101101111",
24085 => "0001101101110000",
24086 => "0001101101110010",
24087 => "0001101101110011",
24088 => "0001101101110101",
24089 => "0001101101110110",
24090 => "0001101101111000",
24091 => "0001101101111001",
24092 => "0001101101111011",
24093 => "0001101101111100",
24094 => "0001101101111110",
24095 => "0001101110000000",
24096 => "0001101110000001",
24097 => "0001101110000011",
24098 => "0001101110000100",
24099 => "0001101110000110",
24100 => "0001101110000111",
24101 => "0001101110001001",
24102 => "0001101110001010",
24103 => "0001101110001100",
24104 => "0001101110001101",
24105 => "0001101110001111",
24106 => "0001101110010000",
24107 => "0001101110010010",
24108 => "0001101110010100",
24109 => "0001101110010101",
24110 => "0001101110010111",
24111 => "0001101110011000",
24112 => "0001101110011010",
24113 => "0001101110011011",
24114 => "0001101110011101",
24115 => "0001101110011110",
24116 => "0001101110100000",
24117 => "0001101110100001",
24118 => "0001101110100011",
24119 => "0001101110100100",
24120 => "0001101110100110",
24121 => "0001101110101000",
24122 => "0001101110101001",
24123 => "0001101110101011",
24124 => "0001101110101100",
24125 => "0001101110101110",
24126 => "0001101110101111",
24127 => "0001101110110001",
24128 => "0001101110110010",
24129 => "0001101110110100",
24130 => "0001101110110101",
24131 => "0001101110110111",
24132 => "0001101110111001",
24133 => "0001101110111010",
24134 => "0001101110111100",
24135 => "0001101110111101",
24136 => "0001101110111111",
24137 => "0001101111000000",
24138 => "0001101111000010",
24139 => "0001101111000011",
24140 => "0001101111000101",
24141 => "0001101111000110",
24142 => "0001101111001000",
24143 => "0001101111001010",
24144 => "0001101111001011",
24145 => "0001101111001101",
24146 => "0001101111001110",
24147 => "0001101111010000",
24148 => "0001101111010001",
24149 => "0001101111010011",
24150 => "0001101111010100",
24151 => "0001101111010110",
24152 => "0001101111010111",
24153 => "0001101111011001",
24154 => "0001101111011011",
24155 => "0001101111011100",
24156 => "0001101111011110",
24157 => "0001101111011111",
24158 => "0001101111100001",
24159 => "0001101111100010",
24160 => "0001101111100100",
24161 => "0001101111100101",
24162 => "0001101111100111",
24163 => "0001101111101001",
24164 => "0001101111101010",
24165 => "0001101111101100",
24166 => "0001101111101101",
24167 => "0001101111101111",
24168 => "0001101111110000",
24169 => "0001101111110010",
24170 => "0001101111110011",
24171 => "0001101111110101",
24172 => "0001101111110111",
24173 => "0001101111111000",
24174 => "0001101111111010",
24175 => "0001101111111011",
24176 => "0001101111111101",
24177 => "0001101111111110",
24178 => "0001110000000000",
24179 => "0001110000000001",
24180 => "0001110000000011",
24181 => "0001110000000101",
24182 => "0001110000000110",
24183 => "0001110000001000",
24184 => "0001110000001001",
24185 => "0001110000001011",
24186 => "0001110000001100",
24187 => "0001110000001110",
24188 => "0001110000010000",
24189 => "0001110000010001",
24190 => "0001110000010011",
24191 => "0001110000010100",
24192 => "0001110000010110",
24193 => "0001110000010111",
24194 => "0001110000011001",
24195 => "0001110000011010",
24196 => "0001110000011100",
24197 => "0001110000011110",
24198 => "0001110000011111",
24199 => "0001110000100001",
24200 => "0001110000100010",
24201 => "0001110000100100",
24202 => "0001110000100101",
24203 => "0001110000100111",
24204 => "0001110000101001",
24205 => "0001110000101010",
24206 => "0001110000101100",
24207 => "0001110000101101",
24208 => "0001110000101111",
24209 => "0001110000110000",
24210 => "0001110000110010",
24211 => "0001110000110100",
24212 => "0001110000110101",
24213 => "0001110000110111",
24214 => "0001110000111000",
24215 => "0001110000111010",
24216 => "0001110000111011",
24217 => "0001110000111101",
24218 => "0001110000111110",
24219 => "0001110001000000",
24220 => "0001110001000010",
24221 => "0001110001000011",
24222 => "0001110001000101",
24223 => "0001110001000110",
24224 => "0001110001001000",
24225 => "0001110001001001",
24226 => "0001110001001011",
24227 => "0001110001001101",
24228 => "0001110001001110",
24229 => "0001110001010000",
24230 => "0001110001010001",
24231 => "0001110001010011",
24232 => "0001110001010101",
24233 => "0001110001010110",
24234 => "0001110001011000",
24235 => "0001110001011001",
24236 => "0001110001011011",
24237 => "0001110001011100",
24238 => "0001110001011110",
24239 => "0001110001100000",
24240 => "0001110001100001",
24241 => "0001110001100011",
24242 => "0001110001100100",
24243 => "0001110001100110",
24244 => "0001110001100111",
24245 => "0001110001101001",
24246 => "0001110001101011",
24247 => "0001110001101100",
24248 => "0001110001101110",
24249 => "0001110001101111",
24250 => "0001110001110001",
24251 => "0001110001110010",
24252 => "0001110001110100",
24253 => "0001110001110110",
24254 => "0001110001110111",
24255 => "0001110001111001",
24256 => "0001110001111010",
24257 => "0001110001111100",
24258 => "0001110001111110",
24259 => "0001110001111111",
24260 => "0001110010000001",
24261 => "0001110010000010",
24262 => "0001110010000100",
24263 => "0001110010000101",
24264 => "0001110010000111",
24265 => "0001110010001001",
24266 => "0001110010001010",
24267 => "0001110010001100",
24268 => "0001110010001101",
24269 => "0001110010001111",
24270 => "0001110010010001",
24271 => "0001110010010010",
24272 => "0001110010010100",
24273 => "0001110010010101",
24274 => "0001110010010111",
24275 => "0001110010011001",
24276 => "0001110010011010",
24277 => "0001110010011100",
24278 => "0001110010011101",
24279 => "0001110010011111",
24280 => "0001110010100000",
24281 => "0001110010100010",
24282 => "0001110010100100",
24283 => "0001110010100101",
24284 => "0001110010100111",
24285 => "0001110010101000",
24286 => "0001110010101010",
24287 => "0001110010101100",
24288 => "0001110010101101",
24289 => "0001110010101111",
24290 => "0001110010110000",
24291 => "0001110010110010",
24292 => "0001110010110100",
24293 => "0001110010110101",
24294 => "0001110010110111",
24295 => "0001110010111000",
24296 => "0001110010111010",
24297 => "0001110010111100",
24298 => "0001110010111101",
24299 => "0001110010111111",
24300 => "0001110011000000",
24301 => "0001110011000010",
24302 => "0001110011000011",
24303 => "0001110011000101",
24304 => "0001110011000111",
24305 => "0001110011001000",
24306 => "0001110011001010",
24307 => "0001110011001011",
24308 => "0001110011001101",
24309 => "0001110011001111",
24310 => "0001110011010000",
24311 => "0001110011010010",
24312 => "0001110011010011",
24313 => "0001110011010101",
24314 => "0001110011010111",
24315 => "0001110011011000",
24316 => "0001110011011010",
24317 => "0001110011011011",
24318 => "0001110011011101",
24319 => "0001110011011111",
24320 => "0001110011100000",
24321 => "0001110011100010",
24322 => "0001110011100011",
24323 => "0001110011100101",
24324 => "0001110011100111",
24325 => "0001110011101000",
24326 => "0001110011101010",
24327 => "0001110011101011",
24328 => "0001110011101101",
24329 => "0001110011101111",
24330 => "0001110011110000",
24331 => "0001110011110010",
24332 => "0001110011110011",
24333 => "0001110011110101",
24334 => "0001110011110111",
24335 => "0001110011111000",
24336 => "0001110011111010",
24337 => "0001110011111100",
24338 => "0001110011111101",
24339 => "0001110011111111",
24340 => "0001110100000000",
24341 => "0001110100000010",
24342 => "0001110100000100",
24343 => "0001110100000101",
24344 => "0001110100000111",
24345 => "0001110100001000",
24346 => "0001110100001010",
24347 => "0001110100001100",
24348 => "0001110100001101",
24349 => "0001110100001111",
24350 => "0001110100010000",
24351 => "0001110100010010",
24352 => "0001110100010100",
24353 => "0001110100010101",
24354 => "0001110100010111",
24355 => "0001110100011000",
24356 => "0001110100011010",
24357 => "0001110100011100",
24358 => "0001110100011101",
24359 => "0001110100011111",
24360 => "0001110100100001",
24361 => "0001110100100010",
24362 => "0001110100100100",
24363 => "0001110100100101",
24364 => "0001110100100111",
24365 => "0001110100101001",
24366 => "0001110100101010",
24367 => "0001110100101100",
24368 => "0001110100101101",
24369 => "0001110100101111",
24370 => "0001110100110001",
24371 => "0001110100110010",
24372 => "0001110100110100",
24373 => "0001110100110110",
24374 => "0001110100110111",
24375 => "0001110100111001",
24376 => "0001110100111010",
24377 => "0001110100111100",
24378 => "0001110100111110",
24379 => "0001110100111111",
24380 => "0001110101000001",
24381 => "0001110101000010",
24382 => "0001110101000100",
24383 => "0001110101000110",
24384 => "0001110101000111",
24385 => "0001110101001001",
24386 => "0001110101001011",
24387 => "0001110101001100",
24388 => "0001110101001110",
24389 => "0001110101001111",
24390 => "0001110101010001",
24391 => "0001110101010011",
24392 => "0001110101010100",
24393 => "0001110101010110",
24394 => "0001110101011000",
24395 => "0001110101011001",
24396 => "0001110101011011",
24397 => "0001110101011100",
24398 => "0001110101011110",
24399 => "0001110101100000",
24400 => "0001110101100001",
24401 => "0001110101100011",
24402 => "0001110101100101",
24403 => "0001110101100110",
24404 => "0001110101101000",
24405 => "0001110101101001",
24406 => "0001110101101011",
24407 => "0001110101101101",
24408 => "0001110101101110",
24409 => "0001110101110000",
24410 => "0001110101110010",
24411 => "0001110101110011",
24412 => "0001110101110101",
24413 => "0001110101110110",
24414 => "0001110101111000",
24415 => "0001110101111010",
24416 => "0001110101111011",
24417 => "0001110101111101",
24418 => "0001110101111111",
24419 => "0001110110000000",
24420 => "0001110110000010",
24421 => "0001110110000100",
24422 => "0001110110000101",
24423 => "0001110110000111",
24424 => "0001110110001000",
24425 => "0001110110001010",
24426 => "0001110110001100",
24427 => "0001110110001101",
24428 => "0001110110001111",
24429 => "0001110110010001",
24430 => "0001110110010010",
24431 => "0001110110010100",
24432 => "0001110110010110",
24433 => "0001110110010111",
24434 => "0001110110011001",
24435 => "0001110110011010",
24436 => "0001110110011100",
24437 => "0001110110011110",
24438 => "0001110110011111",
24439 => "0001110110100001",
24440 => "0001110110100011",
24441 => "0001110110100100",
24442 => "0001110110100110",
24443 => "0001110110101000",
24444 => "0001110110101001",
24445 => "0001110110101011",
24446 => "0001110110101100",
24447 => "0001110110101110",
24448 => "0001110110110000",
24449 => "0001110110110001",
24450 => "0001110110110011",
24451 => "0001110110110101",
24452 => "0001110110110110",
24453 => "0001110110111000",
24454 => "0001110110111010",
24455 => "0001110110111011",
24456 => "0001110110111101",
24457 => "0001110110111110",
24458 => "0001110111000000",
24459 => "0001110111000010",
24460 => "0001110111000011",
24461 => "0001110111000101",
24462 => "0001110111000111",
24463 => "0001110111001000",
24464 => "0001110111001010",
24465 => "0001110111001100",
24466 => "0001110111001101",
24467 => "0001110111001111",
24468 => "0001110111010001",
24469 => "0001110111010010",
24470 => "0001110111010100",
24471 => "0001110111010110",
24472 => "0001110111010111",
24473 => "0001110111011001",
24474 => "0001110111011010",
24475 => "0001110111011100",
24476 => "0001110111011110",
24477 => "0001110111011111",
24478 => "0001110111100001",
24479 => "0001110111100011",
24480 => "0001110111100100",
24481 => "0001110111100110",
24482 => "0001110111101000",
24483 => "0001110111101001",
24484 => "0001110111101011",
24485 => "0001110111101101",
24486 => "0001110111101110",
24487 => "0001110111110000",
24488 => "0001110111110010",
24489 => "0001110111110011",
24490 => "0001110111110101",
24491 => "0001110111110111",
24492 => "0001110111111000",
24493 => "0001110111111010",
24494 => "0001110111111011",
24495 => "0001110111111101",
24496 => "0001110111111111",
24497 => "0001111000000000",
24498 => "0001111000000010",
24499 => "0001111000000100",
24500 => "0001111000000101",
24501 => "0001111000000111",
24502 => "0001111000001001",
24503 => "0001111000001010",
24504 => "0001111000001100",
24505 => "0001111000001110",
24506 => "0001111000001111",
24507 => "0001111000010001",
24508 => "0001111000010011",
24509 => "0001111000010100",
24510 => "0001111000010110",
24511 => "0001111000011000",
24512 => "0001111000011001",
24513 => "0001111000011011",
24514 => "0001111000011101",
24515 => "0001111000011110",
24516 => "0001111000100000",
24517 => "0001111000100010",
24518 => "0001111000100011",
24519 => "0001111000100101",
24520 => "0001111000100111",
24521 => "0001111000101000",
24522 => "0001111000101010",
24523 => "0001111000101100",
24524 => "0001111000101101",
24525 => "0001111000101111",
24526 => "0001111000110001",
24527 => "0001111000110010",
24528 => "0001111000110100",
24529 => "0001111000110110",
24530 => "0001111000110111",
24531 => "0001111000111001",
24532 => "0001111000111011",
24533 => "0001111000111100",
24534 => "0001111000111110",
24535 => "0001111001000000",
24536 => "0001111001000001",
24537 => "0001111001000011",
24538 => "0001111001000101",
24539 => "0001111001000110",
24540 => "0001111001001000",
24541 => "0001111001001010",
24542 => "0001111001001011",
24543 => "0001111001001101",
24544 => "0001111001001111",
24545 => "0001111001010000",
24546 => "0001111001010010",
24547 => "0001111001010100",
24548 => "0001111001010101",
24549 => "0001111001010111",
24550 => "0001111001011001",
24551 => "0001111001011010",
24552 => "0001111001011100",
24553 => "0001111001011110",
24554 => "0001111001011111",
24555 => "0001111001100001",
24556 => "0001111001100011",
24557 => "0001111001100100",
24558 => "0001111001100110",
24559 => "0001111001101000",
24560 => "0001111001101001",
24561 => "0001111001101011",
24562 => "0001111001101101",
24563 => "0001111001101110",
24564 => "0001111001110000",
24565 => "0001111001110010",
24566 => "0001111001110011",
24567 => "0001111001110101",
24568 => "0001111001110111",
24569 => "0001111001111000",
24570 => "0001111001111010",
24571 => "0001111001111100",
24572 => "0001111001111101",
24573 => "0001111001111111",
24574 => "0001111010000001",
24575 => "0001111010000011",
24576 => "0001111010000100",
24577 => "0001111010000110",
24578 => "0001111010001000",
24579 => "0001111010001001",
24580 => "0001111010001011",
24581 => "0001111010001101",
24582 => "0001111010001110",
24583 => "0001111010010000",
24584 => "0001111010010010",
24585 => "0001111010010011",
24586 => "0001111010010101",
24587 => "0001111010010111",
24588 => "0001111010011000",
24589 => "0001111010011010",
24590 => "0001111010011100",
24591 => "0001111010011101",
24592 => "0001111010011111",
24593 => "0001111010100001",
24594 => "0001111010100011",
24595 => "0001111010100100",
24596 => "0001111010100110",
24597 => "0001111010101000",
24598 => "0001111010101001",
24599 => "0001111010101011",
24600 => "0001111010101101",
24601 => "0001111010101110",
24602 => "0001111010110000",
24603 => "0001111010110010",
24604 => "0001111010110011",
24605 => "0001111010110101",
24606 => "0001111010110111",
24607 => "0001111010111000",
24608 => "0001111010111010",
24609 => "0001111010111100",
24610 => "0001111010111110",
24611 => "0001111010111111",
24612 => "0001111011000001",
24613 => "0001111011000011",
24614 => "0001111011000100",
24615 => "0001111011000110",
24616 => "0001111011001000",
24617 => "0001111011001001",
24618 => "0001111011001011",
24619 => "0001111011001101",
24620 => "0001111011001110",
24621 => "0001111011010000",
24622 => "0001111011010010",
24623 => "0001111011010100",
24624 => "0001111011010101",
24625 => "0001111011010111",
24626 => "0001111011011001",
24627 => "0001111011011010",
24628 => "0001111011011100",
24629 => "0001111011011110",
24630 => "0001111011011111",
24631 => "0001111011100001",
24632 => "0001111011100011",
24633 => "0001111011100100",
24634 => "0001111011100110",
24635 => "0001111011101000",
24636 => "0001111011101010",
24637 => "0001111011101011",
24638 => "0001111011101101",
24639 => "0001111011101111",
24640 => "0001111011110000",
24641 => "0001111011110010",
24642 => "0001111011110100",
24643 => "0001111011110101",
24644 => "0001111011110111",
24645 => "0001111011111001",
24646 => "0001111011111011",
24647 => "0001111011111100",
24648 => "0001111011111110",
24649 => "0001111100000000",
24650 => "0001111100000001",
24651 => "0001111100000011",
24652 => "0001111100000101",
24653 => "0001111100000111",
24654 => "0001111100001000",
24655 => "0001111100001010",
24656 => "0001111100001100",
24657 => "0001111100001101",
24658 => "0001111100001111",
24659 => "0001111100010001",
24660 => "0001111100010010",
24661 => "0001111100010100",
24662 => "0001111100010110",
24663 => "0001111100011000",
24664 => "0001111100011001",
24665 => "0001111100011011",
24666 => "0001111100011101",
24667 => "0001111100011110",
24668 => "0001111100100000",
24669 => "0001111100100010",
24670 => "0001111100100100",
24671 => "0001111100100101",
24672 => "0001111100100111",
24673 => "0001111100101001",
24674 => "0001111100101010",
24675 => "0001111100101100",
24676 => "0001111100101110",
24677 => "0001111100101111",
24678 => "0001111100110001",
24679 => "0001111100110011",
24680 => "0001111100110101",
24681 => "0001111100110110",
24682 => "0001111100111000",
24683 => "0001111100111010",
24684 => "0001111100111011",
24685 => "0001111100111101",
24686 => "0001111100111111",
24687 => "0001111101000001",
24688 => "0001111101000010",
24689 => "0001111101000100",
24690 => "0001111101000110",
24691 => "0001111101000111",
24692 => "0001111101001001",
24693 => "0001111101001011",
24694 => "0001111101001101",
24695 => "0001111101001110",
24696 => "0001111101010000",
24697 => "0001111101010010",
24698 => "0001111101010100",
24699 => "0001111101010101",
24700 => "0001111101010111",
24701 => "0001111101011001",
24702 => "0001111101011010",
24703 => "0001111101011100",
24704 => "0001111101011110",
24705 => "0001111101100000",
24706 => "0001111101100001",
24707 => "0001111101100011",
24708 => "0001111101100101",
24709 => "0001111101100110",
24710 => "0001111101101000",
24711 => "0001111101101010",
24712 => "0001111101101100",
24713 => "0001111101101101",
24714 => "0001111101101111",
24715 => "0001111101110001",
24716 => "0001111101110010",
24717 => "0001111101110100",
24718 => "0001111101110110",
24719 => "0001111101111000",
24720 => "0001111101111001",
24721 => "0001111101111011",
24722 => "0001111101111101",
24723 => "0001111101111111",
24724 => "0001111110000000",
24725 => "0001111110000010",
24726 => "0001111110000100",
24727 => "0001111110000101",
24728 => "0001111110000111",
24729 => "0001111110001001",
24730 => "0001111110001011",
24731 => "0001111110001100",
24732 => "0001111110001110",
24733 => "0001111110010000",
24734 => "0001111110010010",
24735 => "0001111110010011",
24736 => "0001111110010101",
24737 => "0001111110010111",
24738 => "0001111110011001",
24739 => "0001111110011010",
24740 => "0001111110011100",
24741 => "0001111110011110",
24742 => "0001111110011111",
24743 => "0001111110100001",
24744 => "0001111110100011",
24745 => "0001111110100101",
24746 => "0001111110100110",
24747 => "0001111110101000",
24748 => "0001111110101010",
24749 => "0001111110101100",
24750 => "0001111110101101",
24751 => "0001111110101111",
24752 => "0001111110110001",
24753 => "0001111110110011",
24754 => "0001111110110100",
24755 => "0001111110110110",
24756 => "0001111110111000",
24757 => "0001111110111001",
24758 => "0001111110111011",
24759 => "0001111110111101",
24760 => "0001111110111111",
24761 => "0001111111000000",
24762 => "0001111111000010",
24763 => "0001111111000100",
24764 => "0001111111000110",
24765 => "0001111111000111",
24766 => "0001111111001001",
24767 => "0001111111001011",
24768 => "0001111111001101",
24769 => "0001111111001110",
24770 => "0001111111010000",
24771 => "0001111111010010",
24772 => "0001111111010100",
24773 => "0001111111010101",
24774 => "0001111111010111",
24775 => "0001111111011001",
24776 => "0001111111011011",
24777 => "0001111111011100",
24778 => "0001111111011110",
24779 => "0001111111100000",
24780 => "0001111111100001",
24781 => "0001111111100011",
24782 => "0001111111100101",
24783 => "0001111111100111",
24784 => "0001111111101000",
24785 => "0001111111101010",
24786 => "0001111111101100",
24787 => "0001111111101110",
24788 => "0001111111101111",
24789 => "0001111111110001",
24790 => "0001111111110011",
24791 => "0001111111110101",
24792 => "0001111111110110",
24793 => "0001111111111000",
24794 => "0001111111111010",
24795 => "0001111111111100",
24796 => "0001111111111101",
24797 => "0001111111111111",
24798 => "0010000000000001",
24799 => "0010000000000011",
24800 => "0010000000000100",
24801 => "0010000000000110",
24802 => "0010000000001000",
24803 => "0010000000001010",
24804 => "0010000000001011",
24805 => "0010000000001101",
24806 => "0010000000001111",
24807 => "0010000000010001",
24808 => "0010000000010010",
24809 => "0010000000010100",
24810 => "0010000000010110",
24811 => "0010000000011000",
24812 => "0010000000011001",
24813 => "0010000000011011",
24814 => "0010000000011101",
24815 => "0010000000011111",
24816 => "0010000000100001",
24817 => "0010000000100010",
24818 => "0010000000100100",
24819 => "0010000000100110",
24820 => "0010000000101000",
24821 => "0010000000101001",
24822 => "0010000000101011",
24823 => "0010000000101101",
24824 => "0010000000101111",
24825 => "0010000000110000",
24826 => "0010000000110010",
24827 => "0010000000110100",
24828 => "0010000000110110",
24829 => "0010000000110111",
24830 => "0010000000111001",
24831 => "0010000000111011",
24832 => "0010000000111101",
24833 => "0010000000111110",
24834 => "0010000001000000",
24835 => "0010000001000010",
24836 => "0010000001000100",
24837 => "0010000001000101",
24838 => "0010000001000111",
24839 => "0010000001001001",
24840 => "0010000001001011",
24841 => "0010000001001101",
24842 => "0010000001001110",
24843 => "0010000001010000",
24844 => "0010000001010010",
24845 => "0010000001010100",
24846 => "0010000001010101",
24847 => "0010000001010111",
24848 => "0010000001011001",
24849 => "0010000001011011",
24850 => "0010000001011100",
24851 => "0010000001011110",
24852 => "0010000001100000",
24853 => "0010000001100010",
24854 => "0010000001100011",
24855 => "0010000001100101",
24856 => "0010000001100111",
24857 => "0010000001101001",
24858 => "0010000001101011",
24859 => "0010000001101100",
24860 => "0010000001101110",
24861 => "0010000001110000",
24862 => "0010000001110010",
24863 => "0010000001110011",
24864 => "0010000001110101",
24865 => "0010000001110111",
24866 => "0010000001111001",
24867 => "0010000001111010",
24868 => "0010000001111100",
24869 => "0010000001111110",
24870 => "0010000010000000",
24871 => "0010000010000010",
24872 => "0010000010000011",
24873 => "0010000010000101",
24874 => "0010000010000111",
24875 => "0010000010001001",
24876 => "0010000010001010",
24877 => "0010000010001100",
24878 => "0010000010001110",
24879 => "0010000010010000",
24880 => "0010000010010010",
24881 => "0010000010010011",
24882 => "0010000010010101",
24883 => "0010000010010111",
24884 => "0010000010011001",
24885 => "0010000010011010",
24886 => "0010000010011100",
24887 => "0010000010011110",
24888 => "0010000010100000",
24889 => "0010000010100010",
24890 => "0010000010100011",
24891 => "0010000010100101",
24892 => "0010000010100111",
24893 => "0010000010101001",
24894 => "0010000010101010",
24895 => "0010000010101100",
24896 => "0010000010101110",
24897 => "0010000010110000",
24898 => "0010000010110010",
24899 => "0010000010110011",
24900 => "0010000010110101",
24901 => "0010000010110111",
24902 => "0010000010111001",
24903 => "0010000010111011",
24904 => "0010000010111100",
24905 => "0010000010111110",
24906 => "0010000011000000",
24907 => "0010000011000010",
24908 => "0010000011000011",
24909 => "0010000011000101",
24910 => "0010000011000111",
24911 => "0010000011001001",
24912 => "0010000011001011",
24913 => "0010000011001100",
24914 => "0010000011001110",
24915 => "0010000011010000",
24916 => "0010000011010010",
24917 => "0010000011010100",
24918 => "0010000011010101",
24919 => "0010000011010111",
24920 => "0010000011011001",
24921 => "0010000011011011",
24922 => "0010000011011100",
24923 => "0010000011011110",
24924 => "0010000011100000",
24925 => "0010000011100010",
24926 => "0010000011100100",
24927 => "0010000011100101",
24928 => "0010000011100111",
24929 => "0010000011101001",
24930 => "0010000011101011",
24931 => "0010000011101101",
24932 => "0010000011101110",
24933 => "0010000011110000",
24934 => "0010000011110010",
24935 => "0010000011110100",
24936 => "0010000011110110",
24937 => "0010000011110111",
24938 => "0010000011111001",
24939 => "0010000011111011",
24940 => "0010000011111101",
24941 => "0010000011111111",
24942 => "0010000100000000",
24943 => "0010000100000010",
24944 => "0010000100000100",
24945 => "0010000100000110",
24946 => "0010000100001000",
24947 => "0010000100001001",
24948 => "0010000100001011",
24949 => "0010000100001101",
24950 => "0010000100001111",
24951 => "0010000100010001",
24952 => "0010000100010010",
24953 => "0010000100010100",
24954 => "0010000100010110",
24955 => "0010000100011000",
24956 => "0010000100011010",
24957 => "0010000100011011",
24958 => "0010000100011101",
24959 => "0010000100011111",
24960 => "0010000100100001",
24961 => "0010000100100011",
24962 => "0010000100100100",
24963 => "0010000100100110",
24964 => "0010000100101000",
24965 => "0010000100101010",
24966 => "0010000100101100",
24967 => "0010000100101101",
24968 => "0010000100101111",
24969 => "0010000100110001",
24970 => "0010000100110011",
24971 => "0010000100110101",
24972 => "0010000100110110",
24973 => "0010000100111000",
24974 => "0010000100111010",
24975 => "0010000100111100",
24976 => "0010000100111110",
24977 => "0010000100111111",
24978 => "0010000101000001",
24979 => "0010000101000011",
24980 => "0010000101000101",
24981 => "0010000101000111",
24982 => "0010000101001000",
24983 => "0010000101001010",
24984 => "0010000101001100",
24985 => "0010000101001110",
24986 => "0010000101010000",
24987 => "0010000101010010",
24988 => "0010000101010011",
24989 => "0010000101010101",
24990 => "0010000101010111",
24991 => "0010000101011001",
24992 => "0010000101011011",
24993 => "0010000101011100",
24994 => "0010000101011110",
24995 => "0010000101100000",
24996 => "0010000101100010",
24997 => "0010000101100100",
24998 => "0010000101100101",
24999 => "0010000101100111",
25000 => "0010000101101001",
25001 => "0010000101101011",
25002 => "0010000101101101",
25003 => "0010000101101111",
25004 => "0010000101110000",
25005 => "0010000101110010",
25006 => "0010000101110100",
25007 => "0010000101110110",
25008 => "0010000101111000",
25009 => "0010000101111001",
25010 => "0010000101111011",
25011 => "0010000101111101",
25012 => "0010000101111111",
25013 => "0010000110000001",
25014 => "0010000110000011",
25015 => "0010000110000100",
25016 => "0010000110000110",
25017 => "0010000110001000",
25018 => "0010000110001010",
25019 => "0010000110001100",
25020 => "0010000110001101",
25021 => "0010000110001111",
25022 => "0010000110010001",
25023 => "0010000110010011",
25024 => "0010000110010101",
25025 => "0010000110010111",
25026 => "0010000110011000",
25027 => "0010000110011010",
25028 => "0010000110011100",
25029 => "0010000110011110",
25030 => "0010000110100000",
25031 => "0010000110100010",
25032 => "0010000110100011",
25033 => "0010000110100101",
25034 => "0010000110100111",
25035 => "0010000110101001",
25036 => "0010000110101011",
25037 => "0010000110101100",
25038 => "0010000110101110",
25039 => "0010000110110000",
25040 => "0010000110110010",
25041 => "0010000110110100",
25042 => "0010000110110110",
25043 => "0010000110110111",
25044 => "0010000110111001",
25045 => "0010000110111011",
25046 => "0010000110111101",
25047 => "0010000110111111",
25048 => "0010000111000001",
25049 => "0010000111000010",
25050 => "0010000111000100",
25051 => "0010000111000110",
25052 => "0010000111001000",
25053 => "0010000111001010",
25054 => "0010000111001100",
25055 => "0010000111001101",
25056 => "0010000111001111",
25057 => "0010000111010001",
25058 => "0010000111010011",
25059 => "0010000111010101",
25060 => "0010000111010111",
25061 => "0010000111011000",
25062 => "0010000111011010",
25063 => "0010000111011100",
25064 => "0010000111011110",
25065 => "0010000111100000",
25066 => "0010000111100010",
25067 => "0010000111100011",
25068 => "0010000111100101",
25069 => "0010000111100111",
25070 => "0010000111101001",
25071 => "0010000111101011",
25072 => "0010000111101101",
25073 => "0010000111101111",
25074 => "0010000111110000",
25075 => "0010000111110010",
25076 => "0010000111110100",
25077 => "0010000111110110",
25078 => "0010000111111000",
25079 => "0010000111111010",
25080 => "0010000111111011",
25081 => "0010000111111101",
25082 => "0010000111111111",
25083 => "0010001000000001",
25084 => "0010001000000011",
25085 => "0010001000000101",
25086 => "0010001000000110",
25087 => "0010001000001000",
25088 => "0010001000001010",
25089 => "0010001000001100",
25090 => "0010001000001110",
25091 => "0010001000010000",
25092 => "0010001000010010",
25093 => "0010001000010011",
25094 => "0010001000010101",
25095 => "0010001000010111",
25096 => "0010001000011001",
25097 => "0010001000011011",
25098 => "0010001000011101",
25099 => "0010001000011110",
25100 => "0010001000100000",
25101 => "0010001000100010",
25102 => "0010001000100100",
25103 => "0010001000100110",
25104 => "0010001000101000",
25105 => "0010001000101010",
25106 => "0010001000101011",
25107 => "0010001000101101",
25108 => "0010001000101111",
25109 => "0010001000110001",
25110 => "0010001000110011",
25111 => "0010001000110101",
25112 => "0010001000110111",
25113 => "0010001000111000",
25114 => "0010001000111010",
25115 => "0010001000111100",
25116 => "0010001000111110",
25117 => "0010001001000000",
25118 => "0010001001000010",
25119 => "0010001001000011",
25120 => "0010001001000101",
25121 => "0010001001000111",
25122 => "0010001001001001",
25123 => "0010001001001011",
25124 => "0010001001001101",
25125 => "0010001001001111",
25126 => "0010001001010000",
25127 => "0010001001010010",
25128 => "0010001001010100",
25129 => "0010001001010110",
25130 => "0010001001011000",
25131 => "0010001001011010",
25132 => "0010001001011100",
25133 => "0010001001011101",
25134 => "0010001001011111",
25135 => "0010001001100001",
25136 => "0010001001100011",
25137 => "0010001001100101",
25138 => "0010001001100111",
25139 => "0010001001101001",
25140 => "0010001001101011",
25141 => "0010001001101100",
25142 => "0010001001101110",
25143 => "0010001001110000",
25144 => "0010001001110010",
25145 => "0010001001110100",
25146 => "0010001001110110",
25147 => "0010001001111000",
25148 => "0010001001111001",
25149 => "0010001001111011",
25150 => "0010001001111101",
25151 => "0010001001111111",
25152 => "0010001010000001",
25153 => "0010001010000011",
25154 => "0010001010000101",
25155 => "0010001010000110",
25156 => "0010001010001000",
25157 => "0010001010001010",
25158 => "0010001010001100",
25159 => "0010001010001110",
25160 => "0010001010010000",
25161 => "0010001010010010",
25162 => "0010001010010100",
25163 => "0010001010010101",
25164 => "0010001010010111",
25165 => "0010001010011001",
25166 => "0010001010011011",
25167 => "0010001010011101",
25168 => "0010001010011111",
25169 => "0010001010100001",
25170 => "0010001010100011",
25171 => "0010001010100100",
25172 => "0010001010100110",
25173 => "0010001010101000",
25174 => "0010001010101010",
25175 => "0010001010101100",
25176 => "0010001010101110",
25177 => "0010001010110000",
25178 => "0010001010110010",
25179 => "0010001010110011",
25180 => "0010001010110101",
25181 => "0010001010110111",
25182 => "0010001010111001",
25183 => "0010001010111011",
25184 => "0010001010111101",
25185 => "0010001010111111",
25186 => "0010001011000001",
25187 => "0010001011000010",
25188 => "0010001011000100",
25189 => "0010001011000110",
25190 => "0010001011001000",
25191 => "0010001011001010",
25192 => "0010001011001100",
25193 => "0010001011001110",
25194 => "0010001011010000",
25195 => "0010001011010001",
25196 => "0010001011010011",
25197 => "0010001011010101",
25198 => "0010001011010111",
25199 => "0010001011011001",
25200 => "0010001011011011",
25201 => "0010001011011101",
25202 => "0010001011011111",
25203 => "0010001011100000",
25204 => "0010001011100010",
25205 => "0010001011100100",
25206 => "0010001011100110",
25207 => "0010001011101000",
25208 => "0010001011101010",
25209 => "0010001011101100",
25210 => "0010001011101110",
25211 => "0010001011110000",
25212 => "0010001011110001",
25213 => "0010001011110011",
25214 => "0010001011110101",
25215 => "0010001011110111",
25216 => "0010001011111001",
25217 => "0010001011111011",
25218 => "0010001011111101",
25219 => "0010001011111111",
25220 => "0010001100000001",
25221 => "0010001100000010",
25222 => "0010001100000100",
25223 => "0010001100000110",
25224 => "0010001100001000",
25225 => "0010001100001010",
25226 => "0010001100001100",
25227 => "0010001100001110",
25228 => "0010001100010000",
25229 => "0010001100010010",
25230 => "0010001100010011",
25231 => "0010001100010101",
25232 => "0010001100010111",
25233 => "0010001100011001",
25234 => "0010001100011011",
25235 => "0010001100011101",
25236 => "0010001100011111",
25237 => "0010001100100001",
25238 => "0010001100100011",
25239 => "0010001100100100",
25240 => "0010001100100110",
25241 => "0010001100101000",
25242 => "0010001100101010",
25243 => "0010001100101100",
25244 => "0010001100101110",
25245 => "0010001100110000",
25246 => "0010001100110010",
25247 => "0010001100110100",
25248 => "0010001100110110",
25249 => "0010001100110111",
25250 => "0010001100111001",
25251 => "0010001100111011",
25252 => "0010001100111101",
25253 => "0010001100111111",
25254 => "0010001101000001",
25255 => "0010001101000011",
25256 => "0010001101000101",
25257 => "0010001101000111",
25258 => "0010001101001001",
25259 => "0010001101001010",
25260 => "0010001101001100",
25261 => "0010001101001110",
25262 => "0010001101010000",
25263 => "0010001101010010",
25264 => "0010001101010100",
25265 => "0010001101010110",
25266 => "0010001101011000",
25267 => "0010001101011010",
25268 => "0010001101011100",
25269 => "0010001101011101",
25270 => "0010001101011111",
25271 => "0010001101100001",
25272 => "0010001101100011",
25273 => "0010001101100101",
25274 => "0010001101100111",
25275 => "0010001101101001",
25276 => "0010001101101011",
25277 => "0010001101101101",
25278 => "0010001101101111",
25279 => "0010001101110001",
25280 => "0010001101110010",
25281 => "0010001101110100",
25282 => "0010001101110110",
25283 => "0010001101111000",
25284 => "0010001101111010",
25285 => "0010001101111100",
25286 => "0010001101111110",
25287 => "0010001110000000",
25288 => "0010001110000010",
25289 => "0010001110000100",
25290 => "0010001110000110",
25291 => "0010001110000111",
25292 => "0010001110001001",
25293 => "0010001110001011",
25294 => "0010001110001101",
25295 => "0010001110001111",
25296 => "0010001110010001",
25297 => "0010001110010011",
25298 => "0010001110010101",
25299 => "0010001110010111",
25300 => "0010001110011001",
25301 => "0010001110011011",
25302 => "0010001110011101",
25303 => "0010001110011110",
25304 => "0010001110100000",
25305 => "0010001110100010",
25306 => "0010001110100100",
25307 => "0010001110100110",
25308 => "0010001110101000",
25309 => "0010001110101010",
25310 => "0010001110101100",
25311 => "0010001110101110",
25312 => "0010001110110000",
25313 => "0010001110110010",
25314 => "0010001110110100",
25315 => "0010001110110101",
25316 => "0010001110110111",
25317 => "0010001110111001",
25318 => "0010001110111011",
25319 => "0010001110111101",
25320 => "0010001110111111",
25321 => "0010001111000001",
25322 => "0010001111000011",
25323 => "0010001111000101",
25324 => "0010001111000111",
25325 => "0010001111001001",
25326 => "0010001111001011",
25327 => "0010001111001101",
25328 => "0010001111001110",
25329 => "0010001111010000",
25330 => "0010001111010010",
25331 => "0010001111010100",
25332 => "0010001111010110",
25333 => "0010001111011000",
25334 => "0010001111011010",
25335 => "0010001111011100",
25336 => "0010001111011110",
25337 => "0010001111100000",
25338 => "0010001111100010",
25339 => "0010001111100100",
25340 => "0010001111100110",
25341 => "0010001111101000",
25342 => "0010001111101001",
25343 => "0010001111101011",
25344 => "0010001111101101",
25345 => "0010001111101111",
25346 => "0010001111110001",
25347 => "0010001111110011",
25348 => "0010001111110101",
25349 => "0010001111110111",
25350 => "0010001111111001",
25351 => "0010001111111011",
25352 => "0010001111111101",
25353 => "0010001111111111",
25354 => "0010010000000001",
25355 => "0010010000000011",
25356 => "0010010000000101",
25357 => "0010010000000110",
25358 => "0010010000001000",
25359 => "0010010000001010",
25360 => "0010010000001100",
25361 => "0010010000001110",
25362 => "0010010000010000",
25363 => "0010010000010010",
25364 => "0010010000010100",
25365 => "0010010000010110",
25366 => "0010010000011000",
25367 => "0010010000011010",
25368 => "0010010000011100",
25369 => "0010010000011110",
25370 => "0010010000100000",
25371 => "0010010000100010",
25372 => "0010010000100100",
25373 => "0010010000100101",
25374 => "0010010000100111",
25375 => "0010010000101001",
25376 => "0010010000101011",
25377 => "0010010000101101",
25378 => "0010010000101111",
25379 => "0010010000110001",
25380 => "0010010000110011",
25381 => "0010010000110101",
25382 => "0010010000110111",
25383 => "0010010000111001",
25384 => "0010010000111011",
25385 => "0010010000111101",
25386 => "0010010000111111",
25387 => "0010010001000001",
25388 => "0010010001000011",
25389 => "0010010001000101",
25390 => "0010010001000110",
25391 => "0010010001001000",
25392 => "0010010001001010",
25393 => "0010010001001100",
25394 => "0010010001001110",
25395 => "0010010001010000",
25396 => "0010010001010010",
25397 => "0010010001010100",
25398 => "0010010001010110",
25399 => "0010010001011000",
25400 => "0010010001011010",
25401 => "0010010001011100",
25402 => "0010010001011110",
25403 => "0010010001100000",
25404 => "0010010001100010",
25405 => "0010010001100100",
25406 => "0010010001100110",
25407 => "0010010001101000",
25408 => "0010010001101010",
25409 => "0010010001101100",
25410 => "0010010001101101",
25411 => "0010010001101111",
25412 => "0010010001110001",
25413 => "0010010001110011",
25414 => "0010010001110101",
25415 => "0010010001110111",
25416 => "0010010001111001",
25417 => "0010010001111011",
25418 => "0010010001111101",
25419 => "0010010001111111",
25420 => "0010010010000001",
25421 => "0010010010000011",
25422 => "0010010010000101",
25423 => "0010010010000111",
25424 => "0010010010001001",
25425 => "0010010010001011",
25426 => "0010010010001101",
25427 => "0010010010001111",
25428 => "0010010010010001",
25429 => "0010010010010011",
25430 => "0010010010010101",
25431 => "0010010010010111",
25432 => "0010010010011001",
25433 => "0010010010011010",
25434 => "0010010010011100",
25435 => "0010010010011110",
25436 => "0010010010100000",
25437 => "0010010010100010",
25438 => "0010010010100100",
25439 => "0010010010100110",
25440 => "0010010010101000",
25441 => "0010010010101010",
25442 => "0010010010101100",
25443 => "0010010010101110",
25444 => "0010010010110000",
25445 => "0010010010110010",
25446 => "0010010010110100",
25447 => "0010010010110110",
25448 => "0010010010111000",
25449 => "0010010010111010",
25450 => "0010010010111100",
25451 => "0010010010111110",
25452 => "0010010011000000",
25453 => "0010010011000010",
25454 => "0010010011000100",
25455 => "0010010011000110",
25456 => "0010010011001000",
25457 => "0010010011001010",
25458 => "0010010011001100",
25459 => "0010010011001110",
25460 => "0010010011010000",
25461 => "0010010011010010",
25462 => "0010010011010011",
25463 => "0010010011010101",
25464 => "0010010011010111",
25465 => "0010010011011001",
25466 => "0010010011011011",
25467 => "0010010011011101",
25468 => "0010010011011111",
25469 => "0010010011100001",
25470 => "0010010011100011",
25471 => "0010010011100101",
25472 => "0010010011100111",
25473 => "0010010011101001",
25474 => "0010010011101011",
25475 => "0010010011101101",
25476 => "0010010011101111",
25477 => "0010010011110001",
25478 => "0010010011110011",
25479 => "0010010011110101",
25480 => "0010010011110111",
25481 => "0010010011111001",
25482 => "0010010011111011",
25483 => "0010010011111101",
25484 => "0010010011111111",
25485 => "0010010100000001",
25486 => "0010010100000011",
25487 => "0010010100000101",
25488 => "0010010100000111",
25489 => "0010010100001001",
25490 => "0010010100001011",
25491 => "0010010100001101",
25492 => "0010010100001111",
25493 => "0010010100010001",
25494 => "0010010100010011",
25495 => "0010010100010101",
25496 => "0010010100010111",
25497 => "0010010100011001",
25498 => "0010010100011011",
25499 => "0010010100011101",
25500 => "0010010100011111",
25501 => "0010010100100001",
25502 => "0010010100100011",
25503 => "0010010100100101",
25504 => "0010010100100111",
25505 => "0010010100101001",
25506 => "0010010100101011",
25507 => "0010010100101101",
25508 => "0010010100101110",
25509 => "0010010100110000",
25510 => "0010010100110010",
25511 => "0010010100110100",
25512 => "0010010100110110",
25513 => "0010010100111000",
25514 => "0010010100111010",
25515 => "0010010100111100",
25516 => "0010010100111110",
25517 => "0010010101000000",
25518 => "0010010101000010",
25519 => "0010010101000100",
25520 => "0010010101000110",
25521 => "0010010101001000",
25522 => "0010010101001010",
25523 => "0010010101001100",
25524 => "0010010101001110",
25525 => "0010010101010000",
25526 => "0010010101010010",
25527 => "0010010101010100",
25528 => "0010010101010110",
25529 => "0010010101011000",
25530 => "0010010101011010",
25531 => "0010010101011100",
25532 => "0010010101011110",
25533 => "0010010101100000",
25534 => "0010010101100010",
25535 => "0010010101100100",
25536 => "0010010101100110",
25537 => "0010010101101000",
25538 => "0010010101101010",
25539 => "0010010101101100",
25540 => "0010010101101110",
25541 => "0010010101110000",
25542 => "0010010101110010",
25543 => "0010010101110100",
25544 => "0010010101110110",
25545 => "0010010101111000",
25546 => "0010010101111010",
25547 => "0010010101111100",
25548 => "0010010101111110",
25549 => "0010010110000000",
25550 => "0010010110000010",
25551 => "0010010110000100",
25552 => "0010010110000110",
25553 => "0010010110001000",
25554 => "0010010110001010",
25555 => "0010010110001100",
25556 => "0010010110001110",
25557 => "0010010110010000",
25558 => "0010010110010010",
25559 => "0010010110010100",
25560 => "0010010110010110",
25561 => "0010010110011000",
25562 => "0010010110011010",
25563 => "0010010110011100",
25564 => "0010010110011110",
25565 => "0010010110100000",
25566 => "0010010110100010",
25567 => "0010010110100100",
25568 => "0010010110100110",
25569 => "0010010110101000",
25570 => "0010010110101010",
25571 => "0010010110101100",
25572 => "0010010110101110",
25573 => "0010010110110000",
25574 => "0010010110110010",
25575 => "0010010110110100",
25576 => "0010010110110110",
25577 => "0010010110111000",
25578 => "0010010110111010",
25579 => "0010010110111100",
25580 => "0010010110111110",
25581 => "0010010111000000",
25582 => "0010010111000010",
25583 => "0010010111000100",
25584 => "0010010111000110",
25585 => "0010010111001000",
25586 => "0010010111001010",
25587 => "0010010111001101",
25588 => "0010010111001111",
25589 => "0010010111010001",
25590 => "0010010111010011",
25591 => "0010010111010101",
25592 => "0010010111010111",
25593 => "0010010111011001",
25594 => "0010010111011011",
25595 => "0010010111011101",
25596 => "0010010111011111",
25597 => "0010010111100001",
25598 => "0010010111100011",
25599 => "0010010111100101",
25600 => "0010010111100111",
25601 => "0010010111101001",
25602 => "0010010111101011",
25603 => "0010010111101101",
25604 => "0010010111101111",
25605 => "0010010111110001",
25606 => "0010010111110011",
25607 => "0010010111110101",
25608 => "0010010111110111",
25609 => "0010010111111001",
25610 => "0010010111111011",
25611 => "0010010111111101",
25612 => "0010010111111111",
25613 => "0010011000000001",
25614 => "0010011000000011",
25615 => "0010011000000101",
25616 => "0010011000000111",
25617 => "0010011000001001",
25618 => "0010011000001011",
25619 => "0010011000001101",
25620 => "0010011000001111",
25621 => "0010011000010001",
25622 => "0010011000010011",
25623 => "0010011000010101",
25624 => "0010011000010111",
25625 => "0010011000011001",
25626 => "0010011000011011",
25627 => "0010011000011101",
25628 => "0010011000011111",
25629 => "0010011000100001",
25630 => "0010011000100011",
25631 => "0010011000100101",
25632 => "0010011000100111",
25633 => "0010011000101010",
25634 => "0010011000101100",
25635 => "0010011000101110",
25636 => "0010011000110000",
25637 => "0010011000110010",
25638 => "0010011000110100",
25639 => "0010011000110110",
25640 => "0010011000111000",
25641 => "0010011000111010",
25642 => "0010011000111100",
25643 => "0010011000111110",
25644 => "0010011001000000",
25645 => "0010011001000010",
25646 => "0010011001000100",
25647 => "0010011001000110",
25648 => "0010011001001000",
25649 => "0010011001001010",
25650 => "0010011001001100",
25651 => "0010011001001110",
25652 => "0010011001010000",
25653 => "0010011001010010",
25654 => "0010011001010100",
25655 => "0010011001010110",
25656 => "0010011001011000",
25657 => "0010011001011010",
25658 => "0010011001011100",
25659 => "0010011001011110",
25660 => "0010011001100000",
25661 => "0010011001100010",
25662 => "0010011001100101",
25663 => "0010011001100111",
25664 => "0010011001101001",
25665 => "0010011001101011",
25666 => "0010011001101101",
25667 => "0010011001101111",
25668 => "0010011001110001",
25669 => "0010011001110011",
25670 => "0010011001110101",
25671 => "0010011001110111",
25672 => "0010011001111001",
25673 => "0010011001111011",
25674 => "0010011001111101",
25675 => "0010011001111111",
25676 => "0010011010000001",
25677 => "0010011010000011",
25678 => "0010011010000101",
25679 => "0010011010000111",
25680 => "0010011010001001",
25681 => "0010011010001011",
25682 => "0010011010001101",
25683 => "0010011010001111",
25684 => "0010011010010001",
25685 => "0010011010010100",
25686 => "0010011010010110",
25687 => "0010011010011000",
25688 => "0010011010011010",
25689 => "0010011010011100",
25690 => "0010011010011110",
25691 => "0010011010100000",
25692 => "0010011010100010",
25693 => "0010011010100100",
25694 => "0010011010100110",
25695 => "0010011010101000",
25696 => "0010011010101010",
25697 => "0010011010101100",
25698 => "0010011010101110",
25699 => "0010011010110000",
25700 => "0010011010110010",
25701 => "0010011010110100",
25702 => "0010011010110110",
25703 => "0010011010111000",
25704 => "0010011010111010",
25705 => "0010011010111101",
25706 => "0010011010111111",
25707 => "0010011011000001",
25708 => "0010011011000011",
25709 => "0010011011000101",
25710 => "0010011011000111",
25711 => "0010011011001001",
25712 => "0010011011001011",
25713 => "0010011011001101",
25714 => "0010011011001111",
25715 => "0010011011010001",
25716 => "0010011011010011",
25717 => "0010011011010101",
25718 => "0010011011010111",
25719 => "0010011011011001",
25720 => "0010011011011011",
25721 => "0010011011011101",
25722 => "0010011011100000",
25723 => "0010011011100010",
25724 => "0010011011100100",
25725 => "0010011011100110",
25726 => "0010011011101000",
25727 => "0010011011101010",
25728 => "0010011011101100",
25729 => "0010011011101110",
25730 => "0010011011110000",
25731 => "0010011011110010",
25732 => "0010011011110100",
25733 => "0010011011110110",
25734 => "0010011011111000",
25735 => "0010011011111010",
25736 => "0010011011111100",
25737 => "0010011011111110",
25738 => "0010011100000001",
25739 => "0010011100000011",
25740 => "0010011100000101",
25741 => "0010011100000111",
25742 => "0010011100001001",
25743 => "0010011100001011",
25744 => "0010011100001101",
25745 => "0010011100001111",
25746 => "0010011100010001",
25747 => "0010011100010011",
25748 => "0010011100010101",
25749 => "0010011100010111",
25750 => "0010011100011001",
25751 => "0010011100011011",
25752 => "0010011100011110",
25753 => "0010011100100000",
25754 => "0010011100100010",
25755 => "0010011100100100",
25756 => "0010011100100110",
25757 => "0010011100101000",
25758 => "0010011100101010",
25759 => "0010011100101100",
25760 => "0010011100101110",
25761 => "0010011100110000",
25762 => "0010011100110010",
25763 => "0010011100110100",
25764 => "0010011100110110",
25765 => "0010011100111000",
25766 => "0010011100111011",
25767 => "0010011100111101",
25768 => "0010011100111111",
25769 => "0010011101000001",
25770 => "0010011101000011",
25771 => "0010011101000101",
25772 => "0010011101000111",
25773 => "0010011101001001",
25774 => "0010011101001011",
25775 => "0010011101001101",
25776 => "0010011101001111",
25777 => "0010011101010001",
25778 => "0010011101010011",
25779 => "0010011101010110",
25780 => "0010011101011000",
25781 => "0010011101011010",
25782 => "0010011101011100",
25783 => "0010011101011110",
25784 => "0010011101100000",
25785 => "0010011101100010",
25786 => "0010011101100100",
25787 => "0010011101100110",
25788 => "0010011101101000",
25789 => "0010011101101010",
25790 => "0010011101101100",
25791 => "0010011101101111",
25792 => "0010011101110001",
25793 => "0010011101110011",
25794 => "0010011101110101",
25795 => "0010011101110111",
25796 => "0010011101111001",
25797 => "0010011101111011",
25798 => "0010011101111101",
25799 => "0010011101111111",
25800 => "0010011110000001",
25801 => "0010011110000011",
25802 => "0010011110000110",
25803 => "0010011110001000",
25804 => "0010011110001010",
25805 => "0010011110001100",
25806 => "0010011110001110",
25807 => "0010011110010000",
25808 => "0010011110010010",
25809 => "0010011110010100",
25810 => "0010011110010110",
25811 => "0010011110011000",
25812 => "0010011110011010",
25813 => "0010011110011101",
25814 => "0010011110011111",
25815 => "0010011110100001",
25816 => "0010011110100011",
25817 => "0010011110100101",
25818 => "0010011110100111",
25819 => "0010011110101001",
25820 => "0010011110101011",
25821 => "0010011110101101",
25822 => "0010011110101111",
25823 => "0010011110110001",
25824 => "0010011110110100",
25825 => "0010011110110110",
25826 => "0010011110111000",
25827 => "0010011110111010",
25828 => "0010011110111100",
25829 => "0010011110111110",
25830 => "0010011111000000",
25831 => "0010011111000010",
25832 => "0010011111000100",
25833 => "0010011111000110",
25834 => "0010011111001001",
25835 => "0010011111001011",
25836 => "0010011111001101",
25837 => "0010011111001111",
25838 => "0010011111010001",
25839 => "0010011111010011",
25840 => "0010011111010101",
25841 => "0010011111010111",
25842 => "0010011111011001",
25843 => "0010011111011011",
25844 => "0010011111011110",
25845 => "0010011111100000",
25846 => "0010011111100010",
25847 => "0010011111100100",
25848 => "0010011111100110",
25849 => "0010011111101000",
25850 => "0010011111101010",
25851 => "0010011111101100",
25852 => "0010011111101110",
25853 => "0010011111110000",
25854 => "0010011111110011",
25855 => "0010011111110101",
25856 => "0010011111110111",
25857 => "0010011111111001",
25858 => "0010011111111011",
25859 => "0010011111111101",
25860 => "0010011111111111",
25861 => "0010100000000001",
25862 => "0010100000000011",
25863 => "0010100000000110",
25864 => "0010100000001000",
25865 => "0010100000001010",
25866 => "0010100000001100",
25867 => "0010100000001110",
25868 => "0010100000010000",
25869 => "0010100000010010",
25870 => "0010100000010100",
25871 => "0010100000010110",
25872 => "0010100000011001",
25873 => "0010100000011011",
25874 => "0010100000011101",
25875 => "0010100000011111",
25876 => "0010100000100001",
25877 => "0010100000100011",
25878 => "0010100000100101",
25879 => "0010100000100111",
25880 => "0010100000101010",
25881 => "0010100000101100",
25882 => "0010100000101110",
25883 => "0010100000110000",
25884 => "0010100000110010",
25885 => "0010100000110100",
25886 => "0010100000110110",
25887 => "0010100000111000",
25888 => "0010100000111010",
25889 => "0010100000111101",
25890 => "0010100000111111",
25891 => "0010100001000001",
25892 => "0010100001000011",
25893 => "0010100001000101",
25894 => "0010100001000111",
25895 => "0010100001001001",
25896 => "0010100001001011",
25897 => "0010100001001110",
25898 => "0010100001010000",
25899 => "0010100001010010",
25900 => "0010100001010100",
25901 => "0010100001010110",
25902 => "0010100001011000",
25903 => "0010100001011010",
25904 => "0010100001011100",
25905 => "0010100001011111",
25906 => "0010100001100001",
25907 => "0010100001100011",
25908 => "0010100001100101",
25909 => "0010100001100111",
25910 => "0010100001101001",
25911 => "0010100001101011",
25912 => "0010100001101101",
25913 => "0010100001110000",
25914 => "0010100001110010",
25915 => "0010100001110100",
25916 => "0010100001110110",
25917 => "0010100001111000",
25918 => "0010100001111010",
25919 => "0010100001111100",
25920 => "0010100001111110",
25921 => "0010100010000001",
25922 => "0010100010000011",
25923 => "0010100010000101",
25924 => "0010100010000111",
25925 => "0010100010001001",
25926 => "0010100010001011",
25927 => "0010100010001101",
25928 => "0010100010010000",
25929 => "0010100010010010",
25930 => "0010100010010100",
25931 => "0010100010010110",
25932 => "0010100010011000",
25933 => "0010100010011010",
25934 => "0010100010011100",
25935 => "0010100010011110",
25936 => "0010100010100001",
25937 => "0010100010100011",
25938 => "0010100010100101",
25939 => "0010100010100111",
25940 => "0010100010101001",
25941 => "0010100010101011",
25942 => "0010100010101101",
25943 => "0010100010110000",
25944 => "0010100010110010",
25945 => "0010100010110100",
25946 => "0010100010110110",
25947 => "0010100010111000",
25948 => "0010100010111010",
25949 => "0010100010111100",
25950 => "0010100010111111",
25951 => "0010100011000001",
25952 => "0010100011000011",
25953 => "0010100011000101",
25954 => "0010100011000111",
25955 => "0010100011001001",
25956 => "0010100011001011",
25957 => "0010100011001110",
25958 => "0010100011010000",
25959 => "0010100011010010",
25960 => "0010100011010100",
25961 => "0010100011010110",
25962 => "0010100011011000",
25963 => "0010100011011010",
25964 => "0010100011011101",
25965 => "0010100011011111",
25966 => "0010100011100001",
25967 => "0010100011100011",
25968 => "0010100011100101",
25969 => "0010100011100111",
25970 => "0010100011101001",
25971 => "0010100011101100",
25972 => "0010100011101110",
25973 => "0010100011110000",
25974 => "0010100011110010",
25975 => "0010100011110100",
25976 => "0010100011110110",
25977 => "0010100011111000",
25978 => "0010100011111011",
25979 => "0010100011111101",
25980 => "0010100011111111",
25981 => "0010100100000001",
25982 => "0010100100000011",
25983 => "0010100100000101",
25984 => "0010100100001000",
25985 => "0010100100001010",
25986 => "0010100100001100",
25987 => "0010100100001110",
25988 => "0010100100010000",
25989 => "0010100100010010",
25990 => "0010100100010100",
25991 => "0010100100010111",
25992 => "0010100100011001",
25993 => "0010100100011011",
25994 => "0010100100011101",
25995 => "0010100100011111",
25996 => "0010100100100001",
25997 => "0010100100100100",
25998 => "0010100100100110",
25999 => "0010100100101000",
26000 => "0010100100101010",
26001 => "0010100100101100",
26002 => "0010100100101110",
26003 => "0010100100110001",
26004 => "0010100100110011",
26005 => "0010100100110101",
26006 => "0010100100110111",
26007 => "0010100100111001",
26008 => "0010100100111011",
26009 => "0010100100111101",
26010 => "0010100101000000",
26011 => "0010100101000010",
26012 => "0010100101000100",
26013 => "0010100101000110",
26014 => "0010100101001000",
26015 => "0010100101001010",
26016 => "0010100101001101",
26017 => "0010100101001111",
26018 => "0010100101010001",
26019 => "0010100101010011",
26020 => "0010100101010101",
26021 => "0010100101010111",
26022 => "0010100101011010",
26023 => "0010100101011100",
26024 => "0010100101011110",
26025 => "0010100101100000",
26026 => "0010100101100010",
26027 => "0010100101100100",
26028 => "0010100101100111",
26029 => "0010100101101001",
26030 => "0010100101101011",
26031 => "0010100101101101",
26032 => "0010100101101111",
26033 => "0010100101110001",
26034 => "0010100101110100",
26035 => "0010100101110110",
26036 => "0010100101111000",
26037 => "0010100101111010",
26038 => "0010100101111100",
26039 => "0010100101111111",
26040 => "0010100110000001",
26041 => "0010100110000011",
26042 => "0010100110000101",
26043 => "0010100110000111",
26044 => "0010100110001001",
26045 => "0010100110001100",
26046 => "0010100110001110",
26047 => "0010100110010000",
26048 => "0010100110010010",
26049 => "0010100110010100",
26050 => "0010100110010110",
26051 => "0010100110011001",
26052 => "0010100110011011",
26053 => "0010100110011101",
26054 => "0010100110011111",
26055 => "0010100110100001",
26056 => "0010100110100100",
26057 => "0010100110100110",
26058 => "0010100110101000",
26059 => "0010100110101010",
26060 => "0010100110101100",
26061 => "0010100110101110",
26062 => "0010100110110001",
26063 => "0010100110110011",
26064 => "0010100110110101",
26065 => "0010100110110111",
26066 => "0010100110111001",
26067 => "0010100110111100",
26068 => "0010100110111110",
26069 => "0010100111000000",
26070 => "0010100111000010",
26071 => "0010100111000100",
26072 => "0010100111000110",
26073 => "0010100111001001",
26074 => "0010100111001011",
26075 => "0010100111001101",
26076 => "0010100111001111",
26077 => "0010100111010001",
26078 => "0010100111010100",
26079 => "0010100111010110",
26080 => "0010100111011000",
26081 => "0010100111011010",
26082 => "0010100111011100",
26083 => "0010100111011110",
26084 => "0010100111100001",
26085 => "0010100111100011",
26086 => "0010100111100101",
26087 => "0010100111100111",
26088 => "0010100111101001",
26089 => "0010100111101100",
26090 => "0010100111101110",
26091 => "0010100111110000",
26092 => "0010100111110010",
26093 => "0010100111110100",
26094 => "0010100111110111",
26095 => "0010100111111001",
26096 => "0010100111111011",
26097 => "0010100111111101",
26098 => "0010100111111111",
26099 => "0010101000000010",
26100 => "0010101000000100",
26101 => "0010101000000110",
26102 => "0010101000001000",
26103 => "0010101000001010",
26104 => "0010101000001101",
26105 => "0010101000001111",
26106 => "0010101000010001",
26107 => "0010101000010011",
26108 => "0010101000010101",
26109 => "0010101000011000",
26110 => "0010101000011010",
26111 => "0010101000011100",
26112 => "0010101000011110",
26113 => "0010101000100000",
26114 => "0010101000100011",
26115 => "0010101000100101",
26116 => "0010101000100111",
26117 => "0010101000101001",
26118 => "0010101000101011",
26119 => "0010101000101110",
26120 => "0010101000110000",
26121 => "0010101000110010",
26122 => "0010101000110100",
26123 => "0010101000110110",
26124 => "0010101000111001",
26125 => "0010101000111011",
26126 => "0010101000111101",
26127 => "0010101000111111",
26128 => "0010101001000001",
26129 => "0010101001000100",
26130 => "0010101001000110",
26131 => "0010101001001000",
26132 => "0010101001001010",
26133 => "0010101001001100",
26134 => "0010101001001111",
26135 => "0010101001010001",
26136 => "0010101001010011",
26137 => "0010101001010101",
26138 => "0010101001010111",
26139 => "0010101001011010",
26140 => "0010101001011100",
26141 => "0010101001011110",
26142 => "0010101001100000",
26143 => "0010101001100010",
26144 => "0010101001100101",
26145 => "0010101001100111",
26146 => "0010101001101001",
26147 => "0010101001101011",
26148 => "0010101001101110",
26149 => "0010101001110000",
26150 => "0010101001110010",
26151 => "0010101001110100",
26152 => "0010101001110110",
26153 => "0010101001111001",
26154 => "0010101001111011",
26155 => "0010101001111101",
26156 => "0010101001111111",
26157 => "0010101010000001",
26158 => "0010101010000100",
26159 => "0010101010000110",
26160 => "0010101010001000",
26161 => "0010101010001010",
26162 => "0010101010001101",
26163 => "0010101010001111",
26164 => "0010101010010001",
26165 => "0010101010010011",
26166 => "0010101010010101",
26167 => "0010101010011000",
26168 => "0010101010011010",
26169 => "0010101010011100",
26170 => "0010101010011110",
26171 => "0010101010100001",
26172 => "0010101010100011",
26173 => "0010101010100101",
26174 => "0010101010100111",
26175 => "0010101010101001",
26176 => "0010101010101100",
26177 => "0010101010101110",
26178 => "0010101010110000",
26179 => "0010101010110010",
26180 => "0010101010110101",
26181 => "0010101010110111",
26182 => "0010101010111001",
26183 => "0010101010111011",
26184 => "0010101010111101",
26185 => "0010101011000000",
26186 => "0010101011000010",
26187 => "0010101011000100",
26188 => "0010101011000110",
26189 => "0010101011001001",
26190 => "0010101011001011",
26191 => "0010101011001101",
26192 => "0010101011001111",
26193 => "0010101011010001",
26194 => "0010101011010100",
26195 => "0010101011010110",
26196 => "0010101011011000",
26197 => "0010101011011010",
26198 => "0010101011011101",
26199 => "0010101011011111",
26200 => "0010101011100001",
26201 => "0010101011100011",
26202 => "0010101011100110",
26203 => "0010101011101000",
26204 => "0010101011101010",
26205 => "0010101011101100",
26206 => "0010101011101110",
26207 => "0010101011110001",
26208 => "0010101011110011",
26209 => "0010101011110101",
26210 => "0010101011110111",
26211 => "0010101011111010",
26212 => "0010101011111100",
26213 => "0010101011111110",
26214 => "0010101100000000",
26215 => "0010101100000011",
26216 => "0010101100000101",
26217 => "0010101100000111",
26218 => "0010101100001001",
26219 => "0010101100001100",
26220 => "0010101100001110",
26221 => "0010101100010000",
26222 => "0010101100010010",
26223 => "0010101100010100",
26224 => "0010101100010111",
26225 => "0010101100011001",
26226 => "0010101100011011",
26227 => "0010101100011101",
26228 => "0010101100100000",
26229 => "0010101100100010",
26230 => "0010101100100100",
26231 => "0010101100100110",
26232 => "0010101100101001",
26233 => "0010101100101011",
26234 => "0010101100101101",
26235 => "0010101100101111",
26236 => "0010101100110010",
26237 => "0010101100110100",
26238 => "0010101100110110",
26239 => "0010101100111000",
26240 => "0010101100111011",
26241 => "0010101100111101",
26242 => "0010101100111111",
26243 => "0010101101000001",
26244 => "0010101101000100",
26245 => "0010101101000110",
26246 => "0010101101001000",
26247 => "0010101101001010",
26248 => "0010101101001101",
26249 => "0010101101001111",
26250 => "0010101101010001",
26251 => "0010101101010011",
26252 => "0010101101010110",
26253 => "0010101101011000",
26254 => "0010101101011010",
26255 => "0010101101011100",
26256 => "0010101101011111",
26257 => "0010101101100001",
26258 => "0010101101100011",
26259 => "0010101101100101",
26260 => "0010101101101000",
26261 => "0010101101101010",
26262 => "0010101101101100",
26263 => "0010101101101110",
26264 => "0010101101110001",
26265 => "0010101101110011",
26266 => "0010101101110101",
26267 => "0010101101110111",
26268 => "0010101101111010",
26269 => "0010101101111100",
26270 => "0010101101111110",
26271 => "0010101110000000",
26272 => "0010101110000011",
26273 => "0010101110000101",
26274 => "0010101110000111",
26275 => "0010101110001001",
26276 => "0010101110001100",
26277 => "0010101110001110",
26278 => "0010101110010000",
26279 => "0010101110010010",
26280 => "0010101110010101",
26281 => "0010101110010111",
26282 => "0010101110011001",
26283 => "0010101110011100",
26284 => "0010101110011110",
26285 => "0010101110100000",
26286 => "0010101110100010",
26287 => "0010101110100101",
26288 => "0010101110100111",
26289 => "0010101110101001",
26290 => "0010101110101011",
26291 => "0010101110101110",
26292 => "0010101110110000",
26293 => "0010101110110010",
26294 => "0010101110110100",
26295 => "0010101110110111",
26296 => "0010101110111001",
26297 => "0010101110111011",
26298 => "0010101110111101",
26299 => "0010101111000000",
26300 => "0010101111000010",
26301 => "0010101111000100",
26302 => "0010101111000111",
26303 => "0010101111001001",
26304 => "0010101111001011",
26305 => "0010101111001101",
26306 => "0010101111010000",
26307 => "0010101111010010",
26308 => "0010101111010100",
26309 => "0010101111010110",
26310 => "0010101111011001",
26311 => "0010101111011011",
26312 => "0010101111011101",
26313 => "0010101111100000",
26314 => "0010101111100010",
26315 => "0010101111100100",
26316 => "0010101111100110",
26317 => "0010101111101001",
26318 => "0010101111101011",
26319 => "0010101111101101",
26320 => "0010101111101111",
26321 => "0010101111110010",
26322 => "0010101111110100",
26323 => "0010101111110110",
26324 => "0010101111111001",
26325 => "0010101111111011",
26326 => "0010101111111101",
26327 => "0010101111111111",
26328 => "0010110000000010",
26329 => "0010110000000100",
26330 => "0010110000000110",
26331 => "0010110000001000",
26332 => "0010110000001011",
26333 => "0010110000001101",
26334 => "0010110000001111",
26335 => "0010110000010010",
26336 => "0010110000010100",
26337 => "0010110000010110",
26338 => "0010110000011000",
26339 => "0010110000011011",
26340 => "0010110000011101",
26341 => "0010110000011111",
26342 => "0010110000100010",
26343 => "0010110000100100",
26344 => "0010110000100110",
26345 => "0010110000101000",
26346 => "0010110000101011",
26347 => "0010110000101101",
26348 => "0010110000101111",
26349 => "0010110000110010",
26350 => "0010110000110100",
26351 => "0010110000110110",
26352 => "0010110000111000",
26353 => "0010110000111011",
26354 => "0010110000111101",
26355 => "0010110000111111",
26356 => "0010110001000010",
26357 => "0010110001000100",
26358 => "0010110001000110",
26359 => "0010110001001000",
26360 => "0010110001001011",
26361 => "0010110001001101",
26362 => "0010110001001111",
26363 => "0010110001010010",
26364 => "0010110001010100",
26365 => "0010110001010110",
26366 => "0010110001011000",
26367 => "0010110001011011",
26368 => "0010110001011101",
26369 => "0010110001011111",
26370 => "0010110001100010",
26371 => "0010110001100100",
26372 => "0010110001100110",
26373 => "0010110001101001",
26374 => "0010110001101011",
26375 => "0010110001101101",
26376 => "0010110001101111",
26377 => "0010110001110010",
26378 => "0010110001110100",
26379 => "0010110001110110",
26380 => "0010110001111001",
26381 => "0010110001111011",
26382 => "0010110001111101",
26383 => "0010110001111111",
26384 => "0010110010000010",
26385 => "0010110010000100",
26386 => "0010110010000110",
26387 => "0010110010001001",
26388 => "0010110010001011",
26389 => "0010110010001101",
26390 => "0010110010010000",
26391 => "0010110010010010",
26392 => "0010110010010100",
26393 => "0010110010010110",
26394 => "0010110010011001",
26395 => "0010110010011011",
26396 => "0010110010011101",
26397 => "0010110010100000",
26398 => "0010110010100010",
26399 => "0010110010100100",
26400 => "0010110010100111",
26401 => "0010110010101001",
26402 => "0010110010101011",
26403 => "0010110010101101",
26404 => "0010110010110000",
26405 => "0010110010110010",
26406 => "0010110010110100",
26407 => "0010110010110111",
26408 => "0010110010111001",
26409 => "0010110010111011",
26410 => "0010110010111110",
26411 => "0010110011000000",
26412 => "0010110011000010",
26413 => "0010110011000101",
26414 => "0010110011000111",
26415 => "0010110011001001",
26416 => "0010110011001011",
26417 => "0010110011001110",
26418 => "0010110011010000",
26419 => "0010110011010010",
26420 => "0010110011010101",
26421 => "0010110011010111",
26422 => "0010110011011001",
26423 => "0010110011011100",
26424 => "0010110011011110",
26425 => "0010110011100000",
26426 => "0010110011100011",
26427 => "0010110011100101",
26428 => "0010110011100111",
26429 => "0010110011101010",
26430 => "0010110011101100",
26431 => "0010110011101110",
26432 => "0010110011110000",
26433 => "0010110011110011",
26434 => "0010110011110101",
26435 => "0010110011110111",
26436 => "0010110011111010",
26437 => "0010110011111100",
26438 => "0010110011111110",
26439 => "0010110100000001",
26440 => "0010110100000011",
26441 => "0010110100000101",
26442 => "0010110100001000",
26443 => "0010110100001010",
26444 => "0010110100001100",
26445 => "0010110100001111",
26446 => "0010110100010001",
26447 => "0010110100010011",
26448 => "0010110100010110",
26449 => "0010110100011000",
26450 => "0010110100011010",
26451 => "0010110100011101",
26452 => "0010110100011111",
26453 => "0010110100100001",
26454 => "0010110100100100",
26455 => "0010110100100110",
26456 => "0010110100101000",
26457 => "0010110100101011",
26458 => "0010110100101101",
26459 => "0010110100101111",
26460 => "0010110100110001",
26461 => "0010110100110100",
26462 => "0010110100110110",
26463 => "0010110100111000",
26464 => "0010110100111011",
26465 => "0010110100111101",
26466 => "0010110100111111",
26467 => "0010110101000010",
26468 => "0010110101000100",
26469 => "0010110101000110",
26470 => "0010110101001001",
26471 => "0010110101001011",
26472 => "0010110101001101",
26473 => "0010110101010000",
26474 => "0010110101010010",
26475 => "0010110101010100",
26476 => "0010110101010111",
26477 => "0010110101011001",
26478 => "0010110101011011",
26479 => "0010110101011110",
26480 => "0010110101100000",
26481 => "0010110101100010",
26482 => "0010110101100101",
26483 => "0010110101100111",
26484 => "0010110101101001",
26485 => "0010110101101100",
26486 => "0010110101101110",
26487 => "0010110101110000",
26488 => "0010110101110011",
26489 => "0010110101110101",
26490 => "0010110101110111",
26491 => "0010110101111010",
26492 => "0010110101111100",
26493 => "0010110101111110",
26494 => "0010110110000001",
26495 => "0010110110000011",
26496 => "0010110110000101",
26497 => "0010110110001000",
26498 => "0010110110001010",
26499 => "0010110110001100",
26500 => "0010110110001111",
26501 => "0010110110010001",
26502 => "0010110110010100",
26503 => "0010110110010110",
26504 => "0010110110011000",
26505 => "0010110110011011",
26506 => "0010110110011101",
26507 => "0010110110011111",
26508 => "0010110110100010",
26509 => "0010110110100100",
26510 => "0010110110100110",
26511 => "0010110110101001",
26512 => "0010110110101011",
26513 => "0010110110101101",
26514 => "0010110110110000",
26515 => "0010110110110010",
26516 => "0010110110110100",
26517 => "0010110110110111",
26518 => "0010110110111001",
26519 => "0010110110111011",
26520 => "0010110110111110",
26521 => "0010110111000000",
26522 => "0010110111000010",
26523 => "0010110111000101",
26524 => "0010110111000111",
26525 => "0010110111001001",
26526 => "0010110111001100",
26527 => "0010110111001110",
26528 => "0010110111010001",
26529 => "0010110111010011",
26530 => "0010110111010101",
26531 => "0010110111011000",
26532 => "0010110111011010",
26533 => "0010110111011100",
26534 => "0010110111011111",
26535 => "0010110111100001",
26536 => "0010110111100011",
26537 => "0010110111100110",
26538 => "0010110111101000",
26539 => "0010110111101010",
26540 => "0010110111101101",
26541 => "0010110111101111",
26542 => "0010110111110001",
26543 => "0010110111110100",
26544 => "0010110111110110",
26545 => "0010110111111001",
26546 => "0010110111111011",
26547 => "0010110111111101",
26548 => "0010111000000000",
26549 => "0010111000000010",
26550 => "0010111000000100",
26551 => "0010111000000111",
26552 => "0010111000001001",
26553 => "0010111000001011",
26554 => "0010111000001110",
26555 => "0010111000010000",
26556 => "0010111000010010",
26557 => "0010111000010101",
26558 => "0010111000010111",
26559 => "0010111000011010",
26560 => "0010111000011100",
26561 => "0010111000011110",
26562 => "0010111000100001",
26563 => "0010111000100011",
26564 => "0010111000100101",
26565 => "0010111000101000",
26566 => "0010111000101010",
26567 => "0010111000101100",
26568 => "0010111000101111",
26569 => "0010111000110001",
26570 => "0010111000110100",
26571 => "0010111000110110",
26572 => "0010111000111000",
26573 => "0010111000111011",
26574 => "0010111000111101",
26575 => "0010111000111111",
26576 => "0010111001000010",
26577 => "0010111001000100",
26578 => "0010111001000111",
26579 => "0010111001001001",
26580 => "0010111001001011",
26581 => "0010111001001110",
26582 => "0010111001010000",
26583 => "0010111001010010",
26584 => "0010111001010101",
26585 => "0010111001010111",
26586 => "0010111001011001",
26587 => "0010111001011100",
26588 => "0010111001011110",
26589 => "0010111001100001",
26590 => "0010111001100011",
26591 => "0010111001100101",
26592 => "0010111001101000",
26593 => "0010111001101010",
26594 => "0010111001101100",
26595 => "0010111001101111",
26596 => "0010111001110001",
26597 => "0010111001110100",
26598 => "0010111001110110",
26599 => "0010111001111000",
26600 => "0010111001111011",
26601 => "0010111001111101",
26602 => "0010111001111111",
26603 => "0010111010000010",
26604 => "0010111010000100",
26605 => "0010111010000111",
26606 => "0010111010001001",
26607 => "0010111010001011",
26608 => "0010111010001110",
26609 => "0010111010010000",
26610 => "0010111010010011",
26611 => "0010111010010101",
26612 => "0010111010010111",
26613 => "0010111010011010",
26614 => "0010111010011100",
26615 => "0010111010011110",
26616 => "0010111010100001",
26617 => "0010111010100011",
26618 => "0010111010100110",
26619 => "0010111010101000",
26620 => "0010111010101010",
26621 => "0010111010101101",
26622 => "0010111010101111",
26623 => "0010111010110010",
26624 => "0010111010110100",
26625 => "0010111010110110",
26626 => "0010111010111001",
26627 => "0010111010111011",
26628 => "0010111010111101",
26629 => "0010111011000000",
26630 => "0010111011000010",
26631 => "0010111011000101",
26632 => "0010111011000111",
26633 => "0010111011001001",
26634 => "0010111011001100",
26635 => "0010111011001110",
26636 => "0010111011010001",
26637 => "0010111011010011",
26638 => "0010111011010101",
26639 => "0010111011011000",
26640 => "0010111011011010",
26641 => "0010111011011101",
26642 => "0010111011011111",
26643 => "0010111011100001",
26644 => "0010111011100100",
26645 => "0010111011100110",
26646 => "0010111011101001",
26647 => "0010111011101011",
26648 => "0010111011101101",
26649 => "0010111011110000",
26650 => "0010111011110010",
26651 => "0010111011110100",
26652 => "0010111011110111",
26653 => "0010111011111001",
26654 => "0010111011111100",
26655 => "0010111011111110",
26656 => "0010111100000000",
26657 => "0010111100000011",
26658 => "0010111100000101",
26659 => "0010111100001000",
26660 => "0010111100001010",
26661 => "0010111100001100",
26662 => "0010111100001111",
26663 => "0010111100010001",
26664 => "0010111100010100",
26665 => "0010111100010110",
26666 => "0010111100011000",
26667 => "0010111100011011",
26668 => "0010111100011101",
26669 => "0010111100100000",
26670 => "0010111100100010",
26671 => "0010111100100100",
26672 => "0010111100100111",
26673 => "0010111100101001",
26674 => "0010111100101100",
26675 => "0010111100101110",
26676 => "0010111100110001",
26677 => "0010111100110011",
26678 => "0010111100110101",
26679 => "0010111100111000",
26680 => "0010111100111010",
26681 => "0010111100111101",
26682 => "0010111100111111",
26683 => "0010111101000001",
26684 => "0010111101000100",
26685 => "0010111101000110",
26686 => "0010111101001001",
26687 => "0010111101001011",
26688 => "0010111101001101",
26689 => "0010111101010000",
26690 => "0010111101010010",
26691 => "0010111101010101",
26692 => "0010111101010111",
26693 => "0010111101011001",
26694 => "0010111101011100",
26695 => "0010111101011110",
26696 => "0010111101100001",
26697 => "0010111101100011",
26698 => "0010111101100110",
26699 => "0010111101101000",
26700 => "0010111101101010",
26701 => "0010111101101101",
26702 => "0010111101101111",
26703 => "0010111101110010",
26704 => "0010111101110100",
26705 => "0010111101110110",
26706 => "0010111101111001",
26707 => "0010111101111011",
26708 => "0010111101111110",
26709 => "0010111110000000",
26710 => "0010111110000011",
26711 => "0010111110000101",
26712 => "0010111110000111",
26713 => "0010111110001010",
26714 => "0010111110001100",
26715 => "0010111110001111",
26716 => "0010111110010001",
26717 => "0010111110010011",
26718 => "0010111110010110",
26719 => "0010111110011000",
26720 => "0010111110011011",
26721 => "0010111110011101",
26722 => "0010111110100000",
26723 => "0010111110100010",
26724 => "0010111110100100",
26725 => "0010111110100111",
26726 => "0010111110101001",
26727 => "0010111110101100",
26728 => "0010111110101110",
26729 => "0010111110110001",
26730 => "0010111110110011",
26731 => "0010111110110101",
26732 => "0010111110111000",
26733 => "0010111110111010",
26734 => "0010111110111101",
26735 => "0010111110111111",
26736 => "0010111111000010",
26737 => "0010111111000100",
26738 => "0010111111000110",
26739 => "0010111111001001",
26740 => "0010111111001011",
26741 => "0010111111001110",
26742 => "0010111111010000",
26743 => "0010111111010011",
26744 => "0010111111010101",
26745 => "0010111111010111",
26746 => "0010111111011010",
26747 => "0010111111011100",
26748 => "0010111111011111",
26749 => "0010111111100001",
26750 => "0010111111100100",
26751 => "0010111111100110",
26752 => "0010111111101000",
26753 => "0010111111101011",
26754 => "0010111111101101",
26755 => "0010111111110000",
26756 => "0010111111110010",
26757 => "0010111111110101",
26758 => "0010111111110111",
26759 => "0010111111111001",
26760 => "0010111111111100",
26761 => "0010111111111110",
26762 => "0011000000000001",
26763 => "0011000000000011",
26764 => "0011000000000110",
26765 => "0011000000001000",
26766 => "0011000000001011",
26767 => "0011000000001101",
26768 => "0011000000001111",
26769 => "0011000000010010",
26770 => "0011000000010100",
26771 => "0011000000010111",
26772 => "0011000000011001",
26773 => "0011000000011100",
26774 => "0011000000011110",
26775 => "0011000000100001",
26776 => "0011000000100011",
26777 => "0011000000100101",
26778 => "0011000000101000",
26779 => "0011000000101010",
26780 => "0011000000101101",
26781 => "0011000000101111",
26782 => "0011000000110010",
26783 => "0011000000110100",
26784 => "0011000000110110",
26785 => "0011000000111001",
26786 => "0011000000111011",
26787 => "0011000000111110",
26788 => "0011000001000000",
26789 => "0011000001000011",
26790 => "0011000001000101",
26791 => "0011000001001000",
26792 => "0011000001001010",
26793 => "0011000001001101",
26794 => "0011000001001111",
26795 => "0011000001010001",
26796 => "0011000001010100",
26797 => "0011000001010110",
26798 => "0011000001011001",
26799 => "0011000001011011",
26800 => "0011000001011110",
26801 => "0011000001100000",
26802 => "0011000001100011",
26803 => "0011000001100101",
26804 => "0011000001100111",
26805 => "0011000001101010",
26806 => "0011000001101100",
26807 => "0011000001101111",
26808 => "0011000001110001",
26809 => "0011000001110100",
26810 => "0011000001110110",
26811 => "0011000001111001",
26812 => "0011000001111011",
26813 => "0011000001111110",
26814 => "0011000010000000",
26815 => "0011000010000011",
26816 => "0011000010000101",
26817 => "0011000010000111",
26818 => "0011000010001010",
26819 => "0011000010001100",
26820 => "0011000010001111",
26821 => "0011000010010001",
26822 => "0011000010010100",
26823 => "0011000010010110",
26824 => "0011000010011001",
26825 => "0011000010011011",
26826 => "0011000010011110",
26827 => "0011000010100000",
26828 => "0011000010100010",
26829 => "0011000010100101",
26830 => "0011000010100111",
26831 => "0011000010101010",
26832 => "0011000010101100",
26833 => "0011000010101111",
26834 => "0011000010110001",
26835 => "0011000010110100",
26836 => "0011000010110110",
26837 => "0011000010111001",
26838 => "0011000010111011",
26839 => "0011000010111110",
26840 => "0011000011000000",
26841 => "0011000011000011",
26842 => "0011000011000101",
26843 => "0011000011000111",
26844 => "0011000011001010",
26845 => "0011000011001100",
26846 => "0011000011001111",
26847 => "0011000011010001",
26848 => "0011000011010100",
26849 => "0011000011010110",
26850 => "0011000011011001",
26851 => "0011000011011011",
26852 => "0011000011011110",
26853 => "0011000011100000",
26854 => "0011000011100011",
26855 => "0011000011100101",
26856 => "0011000011101000",
26857 => "0011000011101010",
26858 => "0011000011101101",
26859 => "0011000011101111",
26860 => "0011000011110001",
26861 => "0011000011110100",
26862 => "0011000011110110",
26863 => "0011000011111001",
26864 => "0011000011111011",
26865 => "0011000011111110",
26866 => "0011000100000000",
26867 => "0011000100000011",
26868 => "0011000100000101",
26869 => "0011000100001000",
26870 => "0011000100001010",
26871 => "0011000100001101",
26872 => "0011000100001111",
26873 => "0011000100010010",
26874 => "0011000100010100",
26875 => "0011000100010111",
26876 => "0011000100011001",
26877 => "0011000100011100",
26878 => "0011000100011110",
26879 => "0011000100100001",
26880 => "0011000100100011",
26881 => "0011000100100110",
26882 => "0011000100101000",
26883 => "0011000100101010",
26884 => "0011000100101101",
26885 => "0011000100101111",
26886 => "0011000100110010",
26887 => "0011000100110100",
26888 => "0011000100110111",
26889 => "0011000100111001",
26890 => "0011000100111100",
26891 => "0011000100111110",
26892 => "0011000101000001",
26893 => "0011000101000011",
26894 => "0011000101000110",
26895 => "0011000101001000",
26896 => "0011000101001011",
26897 => "0011000101001101",
26898 => "0011000101010000",
26899 => "0011000101010010",
26900 => "0011000101010101",
26901 => "0011000101010111",
26902 => "0011000101011010",
26903 => "0011000101011100",
26904 => "0011000101011111",
26905 => "0011000101100001",
26906 => "0011000101100100",
26907 => "0011000101100110",
26908 => "0011000101101001",
26909 => "0011000101101011",
26910 => "0011000101101110",
26911 => "0011000101110000",
26912 => "0011000101110011",
26913 => "0011000101110101",
26914 => "0011000101111000",
26915 => "0011000101111010",
26916 => "0011000101111101",
26917 => "0011000101111111",
26918 => "0011000110000010",
26919 => "0011000110000100",
26920 => "0011000110000111",
26921 => "0011000110001001",
26922 => "0011000110001100",
26923 => "0011000110001110",
26924 => "0011000110010001",
26925 => "0011000110010011",
26926 => "0011000110010110",
26927 => "0011000110011000",
26928 => "0011000110011011",
26929 => "0011000110011101",
26930 => "0011000110100000",
26931 => "0011000110100010",
26932 => "0011000110100101",
26933 => "0011000110100111",
26934 => "0011000110101010",
26935 => "0011000110101100",
26936 => "0011000110101111",
26937 => "0011000110110001",
26938 => "0011000110110100",
26939 => "0011000110110110",
26940 => "0011000110111001",
26941 => "0011000110111011",
26942 => "0011000110111110",
26943 => "0011000111000000",
26944 => "0011000111000011",
26945 => "0011000111000101",
26946 => "0011000111001000",
26947 => "0011000111001010",
26948 => "0011000111001101",
26949 => "0011000111001111",
26950 => "0011000111010010",
26951 => "0011000111010100",
26952 => "0011000111010111",
26953 => "0011000111011001",
26954 => "0011000111011100",
26955 => "0011000111011110",
26956 => "0011000111100001",
26957 => "0011000111100011",
26958 => "0011000111100110",
26959 => "0011000111101000",
26960 => "0011000111101011",
26961 => "0011000111101101",
26962 => "0011000111110000",
26963 => "0011000111110010",
26964 => "0011000111110101",
26965 => "0011000111110111",
26966 => "0011000111111010",
26967 => "0011000111111100",
26968 => "0011000111111111",
26969 => "0011001000000001",
26970 => "0011001000000100",
26971 => "0011001000000110",
26972 => "0011001000001001",
26973 => "0011001000001011",
26974 => "0011001000001110",
26975 => "0011001000010000",
26976 => "0011001000010011",
26977 => "0011001000010110",
26978 => "0011001000011000",
26979 => "0011001000011011",
26980 => "0011001000011101",
26981 => "0011001000100000",
26982 => "0011001000100010",
26983 => "0011001000100101",
26984 => "0011001000100111",
26985 => "0011001000101010",
26986 => "0011001000101100",
26987 => "0011001000101111",
26988 => "0011001000110001",
26989 => "0011001000110100",
26990 => "0011001000110110",
26991 => "0011001000111001",
26992 => "0011001000111011",
26993 => "0011001000111110",
26994 => "0011001001000000",
26995 => "0011001001000011",
26996 => "0011001001000101",
26997 => "0011001001001000",
26998 => "0011001001001010",
26999 => "0011001001001101",
27000 => "0011001001010000",
27001 => "0011001001010010",
27002 => "0011001001010101",
27003 => "0011001001010111",
27004 => "0011001001011010",
27005 => "0011001001011100",
27006 => "0011001001011111",
27007 => "0011001001100001",
27008 => "0011001001100100",
27009 => "0011001001100110",
27010 => "0011001001101001",
27011 => "0011001001101011",
27012 => "0011001001101110",
27013 => "0011001001110000",
27014 => "0011001001110011",
27015 => "0011001001110101",
27016 => "0011001001111000",
27017 => "0011001001111011",
27018 => "0011001001111101",
27019 => "0011001010000000",
27020 => "0011001010000010",
27021 => "0011001010000101",
27022 => "0011001010000111",
27023 => "0011001010001010",
27024 => "0011001010001100",
27025 => "0011001010001111",
27026 => "0011001010010001",
27027 => "0011001010010100",
27028 => "0011001010010110",
27029 => "0011001010011001",
27030 => "0011001010011011",
27031 => "0011001010011110",
27032 => "0011001010100001",
27033 => "0011001010100011",
27034 => "0011001010100110",
27035 => "0011001010101000",
27036 => "0011001010101011",
27037 => "0011001010101101",
27038 => "0011001010110000",
27039 => "0011001010110010",
27040 => "0011001010110101",
27041 => "0011001010110111",
27042 => "0011001010111010",
27043 => "0011001010111101",
27044 => "0011001010111111",
27045 => "0011001011000010",
27046 => "0011001011000100",
27047 => "0011001011000111",
27048 => "0011001011001001",
27049 => "0011001011001100",
27050 => "0011001011001110",
27051 => "0011001011010001",
27052 => "0011001011010011",
27053 => "0011001011010110",
27054 => "0011001011011001",
27055 => "0011001011011011",
27056 => "0011001011011110",
27057 => "0011001011100000",
27058 => "0011001011100011",
27059 => "0011001011100101",
27060 => "0011001011101000",
27061 => "0011001011101010",
27062 => "0011001011101101",
27063 => "0011001011101111",
27064 => "0011001011110010",
27065 => "0011001011110101",
27066 => "0011001011110111",
27067 => "0011001011111010",
27068 => "0011001011111100",
27069 => "0011001011111111",
27070 => "0011001100000001",
27071 => "0011001100000100",
27072 => "0011001100000110",
27073 => "0011001100001001",
27074 => "0011001100001100",
27075 => "0011001100001110",
27076 => "0011001100010001",
27077 => "0011001100010011",
27078 => "0011001100010110",
27079 => "0011001100011000",
27080 => "0011001100011011",
27081 => "0011001100011101",
27082 => "0011001100100000",
27083 => "0011001100100011",
27084 => "0011001100100101",
27085 => "0011001100101000",
27086 => "0011001100101010",
27087 => "0011001100101101",
27088 => "0011001100101111",
27089 => "0011001100110010",
27090 => "0011001100110100",
27091 => "0011001100110111",
27092 => "0011001100111010",
27093 => "0011001100111100",
27094 => "0011001100111111",
27095 => "0011001101000001",
27096 => "0011001101000100",
27097 => "0011001101000110",
27098 => "0011001101001001",
27099 => "0011001101001011",
27100 => "0011001101001110",
27101 => "0011001101010001",
27102 => "0011001101010011",
27103 => "0011001101010110",
27104 => "0011001101011000",
27105 => "0011001101011011",
27106 => "0011001101011101",
27107 => "0011001101100000",
27108 => "0011001101100011",
27109 => "0011001101100101",
27110 => "0011001101101000",
27111 => "0011001101101010",
27112 => "0011001101101101",
27113 => "0011001101101111",
27114 => "0011001101110010",
27115 => "0011001101110101",
27116 => "0011001101110111",
27117 => "0011001101111010",
27118 => "0011001101111100",
27119 => "0011001101111111",
27120 => "0011001110000001",
27121 => "0011001110000100",
27122 => "0011001110000111",
27123 => "0011001110001001",
27124 => "0011001110001100",
27125 => "0011001110001110",
27126 => "0011001110010001",
27127 => "0011001110010011",
27128 => "0011001110010110",
27129 => "0011001110011001",
27130 => "0011001110011011",
27131 => "0011001110011110",
27132 => "0011001110100000",
27133 => "0011001110100011",
27134 => "0011001110100101",
27135 => "0011001110101000",
27136 => "0011001110101011",
27137 => "0011001110101101",
27138 => "0011001110110000",
27139 => "0011001110110010",
27140 => "0011001110110101",
27141 => "0011001110110111",
27142 => "0011001110111010",
27143 => "0011001110111101",
27144 => "0011001110111111",
27145 => "0011001111000010",
27146 => "0011001111000100",
27147 => "0011001111000111",
27148 => "0011001111001010",
27149 => "0011001111001100",
27150 => "0011001111001111",
27151 => "0011001111010001",
27152 => "0011001111010100",
27153 => "0011001111010110",
27154 => "0011001111011001",
27155 => "0011001111011100",
27156 => "0011001111011110",
27157 => "0011001111100001",
27158 => "0011001111100011",
27159 => "0011001111100110",
27160 => "0011001111101001",
27161 => "0011001111101011",
27162 => "0011001111101110",
27163 => "0011001111110000",
27164 => "0011001111110011",
27165 => "0011001111110110",
27166 => "0011001111111000",
27167 => "0011001111111011",
27168 => "0011001111111101",
27169 => "0011010000000000",
27170 => "0011010000000010",
27171 => "0011010000000101",
27172 => "0011010000001000",
27173 => "0011010000001010",
27174 => "0011010000001101",
27175 => "0011010000001111",
27176 => "0011010000010010",
27177 => "0011010000010101",
27178 => "0011010000010111",
27179 => "0011010000011010",
27180 => "0011010000011100",
27181 => "0011010000011111",
27182 => "0011010000100010",
27183 => "0011010000100100",
27184 => "0011010000100111",
27185 => "0011010000101001",
27186 => "0011010000101100",
27187 => "0011010000101111",
27188 => "0011010000110001",
27189 => "0011010000110100",
27190 => "0011010000110110",
27191 => "0011010000111001",
27192 => "0011010000111100",
27193 => "0011010000111110",
27194 => "0011010001000001",
27195 => "0011010001000011",
27196 => "0011010001000110",
27197 => "0011010001001001",
27198 => "0011010001001011",
27199 => "0011010001001110",
27200 => "0011010001010000",
27201 => "0011010001010011",
27202 => "0011010001010110",
27203 => "0011010001011000",
27204 => "0011010001011011",
27205 => "0011010001011101",
27206 => "0011010001100000",
27207 => "0011010001100011",
27208 => "0011010001100101",
27209 => "0011010001101000",
27210 => "0011010001101010",
27211 => "0011010001101101",
27212 => "0011010001110000",
27213 => "0011010001110010",
27214 => "0011010001110101",
27215 => "0011010001110111",
27216 => "0011010001111010",
27217 => "0011010001111101",
27218 => "0011010001111111",
27219 => "0011010010000010",
27220 => "0011010010000100",
27221 => "0011010010000111",
27222 => "0011010010001010",
27223 => "0011010010001100",
27224 => "0011010010001111",
27225 => "0011010010010001",
27226 => "0011010010010100",
27227 => "0011010010010111",
27228 => "0011010010011001",
27229 => "0011010010011100",
27230 => "0011010010011111",
27231 => "0011010010100001",
27232 => "0011010010100100",
27233 => "0011010010100110",
27234 => "0011010010101001",
27235 => "0011010010101100",
27236 => "0011010010101110",
27237 => "0011010010110001",
27238 => "0011010010110011",
27239 => "0011010010110110",
27240 => "0011010010111001",
27241 => "0011010010111011",
27242 => "0011010010111110",
27243 => "0011010011000001",
27244 => "0011010011000011",
27245 => "0011010011000110",
27246 => "0011010011001000",
27247 => "0011010011001011",
27248 => "0011010011001110",
27249 => "0011010011010000",
27250 => "0011010011010011",
27251 => "0011010011010101",
27252 => "0011010011011000",
27253 => "0011010011011011",
27254 => "0011010011011101",
27255 => "0011010011100000",
27256 => "0011010011100011",
27257 => "0011010011100101",
27258 => "0011010011101000",
27259 => "0011010011101010",
27260 => "0011010011101101",
27261 => "0011010011110000",
27262 => "0011010011110010",
27263 => "0011010011110101",
27264 => "0011010011111000",
27265 => "0011010011111010",
27266 => "0011010011111101",
27267 => "0011010011111111",
27268 => "0011010100000010",
27269 => "0011010100000101",
27270 => "0011010100000111",
27271 => "0011010100001010",
27272 => "0011010100001101",
27273 => "0011010100001111",
27274 => "0011010100010010",
27275 => "0011010100010101",
27276 => "0011010100010111",
27277 => "0011010100011010",
27278 => "0011010100011100",
27279 => "0011010100011111",
27280 => "0011010100100010",
27281 => "0011010100100100",
27282 => "0011010100100111",
27283 => "0011010100101010",
27284 => "0011010100101100",
27285 => "0011010100101111",
27286 => "0011010100110001",
27287 => "0011010100110100",
27288 => "0011010100110111",
27289 => "0011010100111001",
27290 => "0011010100111100",
27291 => "0011010100111111",
27292 => "0011010101000001",
27293 => "0011010101000100",
27294 => "0011010101000111",
27295 => "0011010101001001",
27296 => "0011010101001100",
27297 => "0011010101001110",
27298 => "0011010101010001",
27299 => "0011010101010100",
27300 => "0011010101010110",
27301 => "0011010101011001",
27302 => "0011010101011100",
27303 => "0011010101011110",
27304 => "0011010101100001",
27305 => "0011010101100100",
27306 => "0011010101100110",
27307 => "0011010101101001",
27308 => "0011010101101011",
27309 => "0011010101101110",
27310 => "0011010101110001",
27311 => "0011010101110011",
27312 => "0011010101110110",
27313 => "0011010101111001",
27314 => "0011010101111011",
27315 => "0011010101111110",
27316 => "0011010110000001",
27317 => "0011010110000011",
27318 => "0011010110000110",
27319 => "0011010110001001",
27320 => "0011010110001011",
27321 => "0011010110001110",
27322 => "0011010110010001",
27323 => "0011010110010011",
27324 => "0011010110010110",
27325 => "0011010110011000",
27326 => "0011010110011011",
27327 => "0011010110011110",
27328 => "0011010110100000",
27329 => "0011010110100011",
27330 => "0011010110100110",
27331 => "0011010110101000",
27332 => "0011010110101011",
27333 => "0011010110101110",
27334 => "0011010110110000",
27335 => "0011010110110011",
27336 => "0011010110110110",
27337 => "0011010110111000",
27338 => "0011010110111011",
27339 => "0011010110111110",
27340 => "0011010111000000",
27341 => "0011010111000011",
27342 => "0011010111000110",
27343 => "0011010111001000",
27344 => "0011010111001011",
27345 => "0011010111001110",
27346 => "0011010111010000",
27347 => "0011010111010011",
27348 => "0011010111010101",
27349 => "0011010111011000",
27350 => "0011010111011011",
27351 => "0011010111011101",
27352 => "0011010111100000",
27353 => "0011010111100011",
27354 => "0011010111100101",
27355 => "0011010111101000",
27356 => "0011010111101011",
27357 => "0011010111101101",
27358 => "0011010111110000",
27359 => "0011010111110011",
27360 => "0011010111110101",
27361 => "0011010111111000",
27362 => "0011010111111011",
27363 => "0011010111111101",
27364 => "0011011000000000",
27365 => "0011011000000011",
27366 => "0011011000000101",
27367 => "0011011000001000",
27368 => "0011011000001011",
27369 => "0011011000001101",
27370 => "0011011000010000",
27371 => "0011011000010011",
27372 => "0011011000010101",
27373 => "0011011000011000",
27374 => "0011011000011011",
27375 => "0011011000011101",
27376 => "0011011000100000",
27377 => "0011011000100011",
27378 => "0011011000100101",
27379 => "0011011000101000",
27380 => "0011011000101011",
27381 => "0011011000101101",
27382 => "0011011000110000",
27383 => "0011011000110011",
27384 => "0011011000110101",
27385 => "0011011000111000",
27386 => "0011011000111011",
27387 => "0011011000111101",
27388 => "0011011001000000",
27389 => "0011011001000011",
27390 => "0011011001000101",
27391 => "0011011001001000",
27392 => "0011011001001011",
27393 => "0011011001001101",
27394 => "0011011001010000",
27395 => "0011011001010011",
27396 => "0011011001010101",
27397 => "0011011001011000",
27398 => "0011011001011011",
27399 => "0011011001011101",
27400 => "0011011001100000",
27401 => "0011011001100011",
27402 => "0011011001100110",
27403 => "0011011001101000",
27404 => "0011011001101011",
27405 => "0011011001101110",
27406 => "0011011001110000",
27407 => "0011011001110011",
27408 => "0011011001110110",
27409 => "0011011001111000",
27410 => "0011011001111011",
27411 => "0011011001111110",
27412 => "0011011010000000",
27413 => "0011011010000011",
27414 => "0011011010000110",
27415 => "0011011010001000",
27416 => "0011011010001011",
27417 => "0011011010001110",
27418 => "0011011010010000",
27419 => "0011011010010011",
27420 => "0011011010010110",
27421 => "0011011010011000",
27422 => "0011011010011011",
27423 => "0011011010011110",
27424 => "0011011010100001",
27425 => "0011011010100011",
27426 => "0011011010100110",
27427 => "0011011010101001",
27428 => "0011011010101011",
27429 => "0011011010101110",
27430 => "0011011010110001",
27431 => "0011011010110011",
27432 => "0011011010110110",
27433 => "0011011010111001",
27434 => "0011011010111011",
27435 => "0011011010111110",
27436 => "0011011011000001",
27437 => "0011011011000011",
27438 => "0011011011000110",
27439 => "0011011011001001",
27440 => "0011011011001100",
27441 => "0011011011001110",
27442 => "0011011011010001",
27443 => "0011011011010100",
27444 => "0011011011010110",
27445 => "0011011011011001",
27446 => "0011011011011100",
27447 => "0011011011011110",
27448 => "0011011011100001",
27449 => "0011011011100100",
27450 => "0011011011100110",
27451 => "0011011011101001",
27452 => "0011011011101100",
27453 => "0011011011101111",
27454 => "0011011011110001",
27455 => "0011011011110100",
27456 => "0011011011110111",
27457 => "0011011011111001",
27458 => "0011011011111100",
27459 => "0011011011111111",
27460 => "0011011100000001",
27461 => "0011011100000100",
27462 => "0011011100000111",
27463 => "0011011100001010",
27464 => "0011011100001100",
27465 => "0011011100001111",
27466 => "0011011100010010",
27467 => "0011011100010100",
27468 => "0011011100010111",
27469 => "0011011100011010",
27470 => "0011011100011100",
27471 => "0011011100011111",
27472 => "0011011100100010",
27473 => "0011011100100101",
27474 => "0011011100100111",
27475 => "0011011100101010",
27476 => "0011011100101101",
27477 => "0011011100101111",
27478 => "0011011100110010",
27479 => "0011011100110101",
27480 => "0011011100111000",
27481 => "0011011100111010",
27482 => "0011011100111101",
27483 => "0011011101000000",
27484 => "0011011101000010",
27485 => "0011011101000101",
27486 => "0011011101001000",
27487 => "0011011101001010",
27488 => "0011011101001101",
27489 => "0011011101010000",
27490 => "0011011101010011",
27491 => "0011011101010101",
27492 => "0011011101011000",
27493 => "0011011101011011",
27494 => "0011011101011101",
27495 => "0011011101100000",
27496 => "0011011101100011",
27497 => "0011011101100110",
27498 => "0011011101101000",
27499 => "0011011101101011",
27500 => "0011011101101110",
27501 => "0011011101110000",
27502 => "0011011101110011",
27503 => "0011011101110110",
27504 => "0011011101111001",
27505 => "0011011101111011",
27506 => "0011011101111110",
27507 => "0011011110000001",
27508 => "0011011110000011",
27509 => "0011011110000110",
27510 => "0011011110001001",
27511 => "0011011110001100",
27512 => "0011011110001110",
27513 => "0011011110010001",
27514 => "0011011110010100",
27515 => "0011011110010110",
27516 => "0011011110011001",
27517 => "0011011110011100",
27518 => "0011011110011111",
27519 => "0011011110100001",
27520 => "0011011110100100",
27521 => "0011011110100111",
27522 => "0011011110101010",
27523 => "0011011110101100",
27524 => "0011011110101111",
27525 => "0011011110110010",
27526 => "0011011110110100",
27527 => "0011011110110111",
27528 => "0011011110111010",
27529 => "0011011110111101",
27530 => "0011011110111111",
27531 => "0011011111000010",
27532 => "0011011111000101",
27533 => "0011011111000111",
27534 => "0011011111001010",
27535 => "0011011111001101",
27536 => "0011011111010000",
27537 => "0011011111010010",
27538 => "0011011111010101",
27539 => "0011011111011000",
27540 => "0011011111011011",
27541 => "0011011111011101",
27542 => "0011011111100000",
27543 => "0011011111100011",
27544 => "0011011111100110",
27545 => "0011011111101000",
27546 => "0011011111101011",
27547 => "0011011111101110",
27548 => "0011011111110000",
27549 => "0011011111110011",
27550 => "0011011111110110",
27551 => "0011011111111001",
27552 => "0011011111111011",
27553 => "0011011111111110",
27554 => "0011100000000001",
27555 => "0011100000000100",
27556 => "0011100000000110",
27557 => "0011100000001001",
27558 => "0011100000001100",
27559 => "0011100000001111",
27560 => "0011100000010001",
27561 => "0011100000010100",
27562 => "0011100000010111",
27563 => "0011100000011001",
27564 => "0011100000011100",
27565 => "0011100000011111",
27566 => "0011100000100010",
27567 => "0011100000100100",
27568 => "0011100000100111",
27569 => "0011100000101010",
27570 => "0011100000101101",
27571 => "0011100000101111",
27572 => "0011100000110010",
27573 => "0011100000110101",
27574 => "0011100000111000",
27575 => "0011100000111010",
27576 => "0011100000111101",
27577 => "0011100001000000",
27578 => "0011100001000011",
27579 => "0011100001000101",
27580 => "0011100001001000",
27581 => "0011100001001011",
27582 => "0011100001001110",
27583 => "0011100001010000",
27584 => "0011100001010011",
27585 => "0011100001010110",
27586 => "0011100001011001",
27587 => "0011100001011011",
27588 => "0011100001011110",
27589 => "0011100001100001",
27590 => "0011100001100100",
27591 => "0011100001100110",
27592 => "0011100001101001",
27593 => "0011100001101100",
27594 => "0011100001101111",
27595 => "0011100001110001",
27596 => "0011100001110100",
27597 => "0011100001110111",
27598 => "0011100001111010",
27599 => "0011100001111100",
27600 => "0011100001111111",
27601 => "0011100010000010",
27602 => "0011100010000101",
27603 => "0011100010000111",
27604 => "0011100010001010",
27605 => "0011100010001101",
27606 => "0011100010010000",
27607 => "0011100010010010",
27608 => "0011100010010101",
27609 => "0011100010011000",
27610 => "0011100010011011",
27611 => "0011100010011101",
27612 => "0011100010100000",
27613 => "0011100010100011",
27614 => "0011100010100110",
27615 => "0011100010101000",
27616 => "0011100010101011",
27617 => "0011100010101110",
27618 => "0011100010110001",
27619 => "0011100010110011",
27620 => "0011100010110110",
27621 => "0011100010111001",
27622 => "0011100010111100",
27623 => "0011100010111110",
27624 => "0011100011000001",
27625 => "0011100011000100",
27626 => "0011100011000111",
27627 => "0011100011001001",
27628 => "0011100011001100",
27629 => "0011100011001111",
27630 => "0011100011010010",
27631 => "0011100011010101",
27632 => "0011100011010111",
27633 => "0011100011011010",
27634 => "0011100011011101",
27635 => "0011100011100000",
27636 => "0011100011100010",
27637 => "0011100011100101",
27638 => "0011100011101000",
27639 => "0011100011101011",
27640 => "0011100011101101",
27641 => "0011100011110000",
27642 => "0011100011110011",
27643 => "0011100011110110",
27644 => "0011100011111000",
27645 => "0011100011111011",
27646 => "0011100011111110",
27647 => "0011100100000001",
27648 => "0011100100000100",
27649 => "0011100100000110",
27650 => "0011100100001001",
27651 => "0011100100001100",
27652 => "0011100100001111",
27653 => "0011100100010001",
27654 => "0011100100010100",
27655 => "0011100100010111",
27656 => "0011100100011010",
27657 => "0011100100011100",
27658 => "0011100100011111",
27659 => "0011100100100010",
27660 => "0011100100100101",
27661 => "0011100100101000",
27662 => "0011100100101010",
27663 => "0011100100101101",
27664 => "0011100100110000",
27665 => "0011100100110011",
27666 => "0011100100110101",
27667 => "0011100100111000",
27668 => "0011100100111011",
27669 => "0011100100111110",
27670 => "0011100101000001",
27671 => "0011100101000011",
27672 => "0011100101000110",
27673 => "0011100101001001",
27674 => "0011100101001100",
27675 => "0011100101001110",
27676 => "0011100101010001",
27677 => "0011100101010100",
27678 => "0011100101010111",
27679 => "0011100101011010",
27680 => "0011100101011100",
27681 => "0011100101011111",
27682 => "0011100101100010",
27683 => "0011100101100101",
27684 => "0011100101101000",
27685 => "0011100101101010",
27686 => "0011100101101101",
27687 => "0011100101110000",
27688 => "0011100101110011",
27689 => "0011100101110101",
27690 => "0011100101111000",
27691 => "0011100101111011",
27692 => "0011100101111110",
27693 => "0011100110000001",
27694 => "0011100110000011",
27695 => "0011100110000110",
27696 => "0011100110001001",
27697 => "0011100110001100",
27698 => "0011100110001111",
27699 => "0011100110010001",
27700 => "0011100110010100",
27701 => "0011100110010111",
27702 => "0011100110011010",
27703 => "0011100110011100",
27704 => "0011100110011111",
27705 => "0011100110100010",
27706 => "0011100110100101",
27707 => "0011100110101000",
27708 => "0011100110101010",
27709 => "0011100110101101",
27710 => "0011100110110000",
27711 => "0011100110110011",
27712 => "0011100110110110",
27713 => "0011100110111000",
27714 => "0011100110111011",
27715 => "0011100110111110",
27716 => "0011100111000001",
27717 => "0011100111000100",
27718 => "0011100111000110",
27719 => "0011100111001001",
27720 => "0011100111001100",
27721 => "0011100111001111",
27722 => "0011100111010010",
27723 => "0011100111010100",
27724 => "0011100111010111",
27725 => "0011100111011010",
27726 => "0011100111011101",
27727 => "0011100111100000",
27728 => "0011100111100010",
27729 => "0011100111100101",
27730 => "0011100111101000",
27731 => "0011100111101011",
27732 => "0011100111101110",
27733 => "0011100111110000",
27734 => "0011100111110011",
27735 => "0011100111110110",
27736 => "0011100111111001",
27737 => "0011100111111100",
27738 => "0011100111111110",
27739 => "0011101000000001",
27740 => "0011101000000100",
27741 => "0011101000000111",
27742 => "0011101000001010",
27743 => "0011101000001100",
27744 => "0011101000001111",
27745 => "0011101000010010",
27746 => "0011101000010101",
27747 => "0011101000011000",
27748 => "0011101000011010",
27749 => "0011101000011101",
27750 => "0011101000100000",
27751 => "0011101000100011",
27752 => "0011101000100110",
27753 => "0011101000101000",
27754 => "0011101000101011",
27755 => "0011101000101110",
27756 => "0011101000110001",
27757 => "0011101000110100",
27758 => "0011101000110110",
27759 => "0011101000111001",
27760 => "0011101000111100",
27761 => "0011101000111111",
27762 => "0011101001000010",
27763 => "0011101001000101",
27764 => "0011101001000111",
27765 => "0011101001001010",
27766 => "0011101001001101",
27767 => "0011101001010000",
27768 => "0011101001010011",
27769 => "0011101001010101",
27770 => "0011101001011000",
27771 => "0011101001011011",
27772 => "0011101001011110",
27773 => "0011101001100001",
27774 => "0011101001100100",
27775 => "0011101001100110",
27776 => "0011101001101001",
27777 => "0011101001101100",
27778 => "0011101001101111",
27779 => "0011101001110010",
27780 => "0011101001110100",
27781 => "0011101001110111",
27782 => "0011101001111010",
27783 => "0011101001111101",
27784 => "0011101010000000",
27785 => "0011101010000011",
27786 => "0011101010000101",
27787 => "0011101010001000",
27788 => "0011101010001011",
27789 => "0011101010001110",
27790 => "0011101010010001",
27791 => "0011101010010011",
27792 => "0011101010010110",
27793 => "0011101010011001",
27794 => "0011101010011100",
27795 => "0011101010011111",
27796 => "0011101010100010",
27797 => "0011101010100100",
27798 => "0011101010100111",
27799 => "0011101010101010",
27800 => "0011101010101101",
27801 => "0011101010110000",
27802 => "0011101010110011",
27803 => "0011101010110101",
27804 => "0011101010111000",
27805 => "0011101010111011",
27806 => "0011101010111110",
27807 => "0011101011000001",
27808 => "0011101011000100",
27809 => "0011101011000110",
27810 => "0011101011001001",
27811 => "0011101011001100",
27812 => "0011101011001111",
27813 => "0011101011010010",
27814 => "0011101011010101",
27815 => "0011101011010111",
27816 => "0011101011011010",
27817 => "0011101011011101",
27818 => "0011101011100000",
27819 => "0011101011100011",
27820 => "0011101011100110",
27821 => "0011101011101000",
27822 => "0011101011101011",
27823 => "0011101011101110",
27824 => "0011101011110001",
27825 => "0011101011110100",
27826 => "0011101011110111",
27827 => "0011101011111001",
27828 => "0011101011111100",
27829 => "0011101011111111",
27830 => "0011101100000010",
27831 => "0011101100000101",
27832 => "0011101100001000",
27833 => "0011101100001010",
27834 => "0011101100001101",
27835 => "0011101100010000",
27836 => "0011101100010011",
27837 => "0011101100010110",
27838 => "0011101100011001",
27839 => "0011101100011011",
27840 => "0011101100011110",
27841 => "0011101100100001",
27842 => "0011101100100100",
27843 => "0011101100100111",
27844 => "0011101100101010",
27845 => "0011101100101100",
27846 => "0011101100101111",
27847 => "0011101100110010",
27848 => "0011101100110101",
27849 => "0011101100111000",
27850 => "0011101100111011",
27851 => "0011101100111110",
27852 => "0011101101000000",
27853 => "0011101101000011",
27854 => "0011101101000110",
27855 => "0011101101001001",
27856 => "0011101101001100",
27857 => "0011101101001111",
27858 => "0011101101010001",
27859 => "0011101101010100",
27860 => "0011101101010111",
27861 => "0011101101011010",
27862 => "0011101101011101",
27863 => "0011101101100000",
27864 => "0011101101100011",
27865 => "0011101101100101",
27866 => "0011101101101000",
27867 => "0011101101101011",
27868 => "0011101101101110",
27869 => "0011101101110001",
27870 => "0011101101110100",
27871 => "0011101101110111",
27872 => "0011101101111001",
27873 => "0011101101111100",
27874 => "0011101101111111",
27875 => "0011101110000010",
27876 => "0011101110000101",
27877 => "0011101110001000",
27878 => "0011101110001011",
27879 => "0011101110001101",
27880 => "0011101110010000",
27881 => "0011101110010011",
27882 => "0011101110010110",
27883 => "0011101110011001",
27884 => "0011101110011100",
27885 => "0011101110011111",
27886 => "0011101110100001",
27887 => "0011101110100100",
27888 => "0011101110100111",
27889 => "0011101110101010",
27890 => "0011101110101101",
27891 => "0011101110110000",
27892 => "0011101110110011",
27893 => "0011101110110101",
27894 => "0011101110111000",
27895 => "0011101110111011",
27896 => "0011101110111110",
27897 => "0011101111000001",
27898 => "0011101111000100",
27899 => "0011101111000111",
27900 => "0011101111001001",
27901 => "0011101111001100",
27902 => "0011101111001111",
27903 => "0011101111010010",
27904 => "0011101111010101",
27905 => "0011101111011000",
27906 => "0011101111011011",
27907 => "0011101111011101",
27908 => "0011101111100000",
27909 => "0011101111100011",
27910 => "0011101111100110",
27911 => "0011101111101001",
27912 => "0011101111101100",
27913 => "0011101111101111",
27914 => "0011101111110010",
27915 => "0011101111110100",
27916 => "0011101111110111",
27917 => "0011101111111010",
27918 => "0011101111111101",
27919 => "0011110000000000",
27920 => "0011110000000011",
27921 => "0011110000000110",
27922 => "0011110000001001",
27923 => "0011110000001011",
27924 => "0011110000001110",
27925 => "0011110000010001",
27926 => "0011110000010100",
27927 => "0011110000010111",
27928 => "0011110000011010",
27929 => "0011110000011101",
27930 => "0011110000100000",
27931 => "0011110000100010",
27932 => "0011110000100101",
27933 => "0011110000101000",
27934 => "0011110000101011",
27935 => "0011110000101110",
27936 => "0011110000110001",
27937 => "0011110000110100",
27938 => "0011110000110111",
27939 => "0011110000111001",
27940 => "0011110000111100",
27941 => "0011110000111111",
27942 => "0011110001000010",
27943 => "0011110001000101",
27944 => "0011110001001000",
27945 => "0011110001001011",
27946 => "0011110001001110",
27947 => "0011110001010000",
27948 => "0011110001010011",
27949 => "0011110001010110",
27950 => "0011110001011001",
27951 => "0011110001011100",
27952 => "0011110001011111",
27953 => "0011110001100010",
27954 => "0011110001100101",
27955 => "0011110001101000",
27956 => "0011110001101010",
27957 => "0011110001101101",
27958 => "0011110001110000",
27959 => "0011110001110011",
27960 => "0011110001110110",
27961 => "0011110001111001",
27962 => "0011110001111100",
27963 => "0011110001111111",
27964 => "0011110010000010",
27965 => "0011110010000100",
27966 => "0011110010000111",
27967 => "0011110010001010",
27968 => "0011110010001101",
27969 => "0011110010010000",
27970 => "0011110010010011",
27971 => "0011110010010110",
27972 => "0011110010011001",
27973 => "0011110010011100",
27974 => "0011110010011110",
27975 => "0011110010100001",
27976 => "0011110010100100",
27977 => "0011110010100111",
27978 => "0011110010101010",
27979 => "0011110010101101",
27980 => "0011110010110000",
27981 => "0011110010110011",
27982 => "0011110010110110",
27983 => "0011110010111000",
27984 => "0011110010111011",
27985 => "0011110010111110",
27986 => "0011110011000001",
27987 => "0011110011000100",
27988 => "0011110011000111",
27989 => "0011110011001010",
27990 => "0011110011001101",
27991 => "0011110011010000",
27992 => "0011110011010011",
27993 => "0011110011010101",
27994 => "0011110011011000",
27995 => "0011110011011011",
27996 => "0011110011011110",
27997 => "0011110011100001",
27998 => "0011110011100100",
27999 => "0011110011100111",
28000 => "0011110011101010",
28001 => "0011110011101101",
28002 => "0011110011110000",
28003 => "0011110011110010",
28004 => "0011110011110101",
28005 => "0011110011111000",
28006 => "0011110011111011",
28007 => "0011110011111110",
28008 => "0011110100000001",
28009 => "0011110100000100",
28010 => "0011110100000111",
28011 => "0011110100001010",
28012 => "0011110100001101",
28013 => "0011110100001111",
28014 => "0011110100010010",
28015 => "0011110100010101",
28016 => "0011110100011000",
28017 => "0011110100011011",
28018 => "0011110100011110",
28019 => "0011110100100001",
28020 => "0011110100100100",
28021 => "0011110100100111",
28022 => "0011110100101010",
28023 => "0011110100101101",
28024 => "0011110100101111",
28025 => "0011110100110010",
28026 => "0011110100110101",
28027 => "0011110100111000",
28028 => "0011110100111011",
28029 => "0011110100111110",
28030 => "0011110101000001",
28031 => "0011110101000100",
28032 => "0011110101000111",
28033 => "0011110101001010",
28034 => "0011110101001101",
28035 => "0011110101001111",
28036 => "0011110101010010",
28037 => "0011110101010101",
28038 => "0011110101011000",
28039 => "0011110101011011",
28040 => "0011110101011110",
28041 => "0011110101100001",
28042 => "0011110101100100",
28043 => "0011110101100111",
28044 => "0011110101101010",
28045 => "0011110101101101",
28046 => "0011110101110000",
28047 => "0011110101110010",
28048 => "0011110101110101",
28049 => "0011110101111000",
28050 => "0011110101111011",
28051 => "0011110101111110",
28052 => "0011110110000001",
28053 => "0011110110000100",
28054 => "0011110110000111",
28055 => "0011110110001010",
28056 => "0011110110001101",
28057 => "0011110110010000",
28058 => "0011110110010011",
28059 => "0011110110010110",
28060 => "0011110110011000",
28061 => "0011110110011011",
28062 => "0011110110011110",
28063 => "0011110110100001",
28064 => "0011110110100100",
28065 => "0011110110100111",
28066 => "0011110110101010",
28067 => "0011110110101101",
28068 => "0011110110110000",
28069 => "0011110110110011",
28070 => "0011110110110110",
28071 => "0011110110111001",
28072 => "0011110110111100",
28073 => "0011110110111110",
28074 => "0011110111000001",
28075 => "0011110111000100",
28076 => "0011110111000111",
28077 => "0011110111001010",
28078 => "0011110111001101",
28079 => "0011110111010000",
28080 => "0011110111010011",
28081 => "0011110111010110",
28082 => "0011110111011001",
28083 => "0011110111011100",
28084 => "0011110111011111",
28085 => "0011110111100010",
28086 => "0011110111100101",
28087 => "0011110111101000",
28088 => "0011110111101010",
28089 => "0011110111101101",
28090 => "0011110111110000",
28091 => "0011110111110011",
28092 => "0011110111110110",
28093 => "0011110111111001",
28094 => "0011110111111100",
28095 => "0011110111111111",
28096 => "0011111000000010",
28097 => "0011111000000101",
28098 => "0011111000001000",
28099 => "0011111000001011",
28100 => "0011111000001110",
28101 => "0011111000010001",
28102 => "0011111000010100",
28103 => "0011111000010111",
28104 => "0011111000011001",
28105 => "0011111000011100",
28106 => "0011111000011111",
28107 => "0011111000100010",
28108 => "0011111000100101",
28109 => "0011111000101000",
28110 => "0011111000101011",
28111 => "0011111000101110",
28112 => "0011111000110001",
28113 => "0011111000110100",
28114 => "0011111000110111",
28115 => "0011111000111010",
28116 => "0011111000111101",
28117 => "0011111001000000",
28118 => "0011111001000011",
28119 => "0011111001000110",
28120 => "0011111001001001",
28121 => "0011111001001011",
28122 => "0011111001001110",
28123 => "0011111001010001",
28124 => "0011111001010100",
28125 => "0011111001010111",
28126 => "0011111001011010",
28127 => "0011111001011101",
28128 => "0011111001100000",
28129 => "0011111001100011",
28130 => "0011111001100110",
28131 => "0011111001101001",
28132 => "0011111001101100",
28133 => "0011111001101111",
28134 => "0011111001110010",
28135 => "0011111001110101",
28136 => "0011111001111000",
28137 => "0011111001111011",
28138 => "0011111001111110",
28139 => "0011111010000001",
28140 => "0011111010000100",
28141 => "0011111010000110",
28142 => "0011111010001001",
28143 => "0011111010001100",
28144 => "0011111010001111",
28145 => "0011111010010010",
28146 => "0011111010010101",
28147 => "0011111010011000",
28148 => "0011111010011011",
28149 => "0011111010011110",
28150 => "0011111010100001",
28151 => "0011111010100100",
28152 => "0011111010100111",
28153 => "0011111010101010",
28154 => "0011111010101101",
28155 => "0011111010110000",
28156 => "0011111010110011",
28157 => "0011111010110110",
28158 => "0011111010111001",
28159 => "0011111010111100",
28160 => "0011111010111111",
28161 => "0011111011000010",
28162 => "0011111011000101",
28163 => "0011111011001000",
28164 => "0011111011001011",
28165 => "0011111011001101",
28166 => "0011111011010000",
28167 => "0011111011010011",
28168 => "0011111011010110",
28169 => "0011111011011001",
28170 => "0011111011011100",
28171 => "0011111011011111",
28172 => "0011111011100010",
28173 => "0011111011100101",
28174 => "0011111011101000",
28175 => "0011111011101011",
28176 => "0011111011101110",
28177 => "0011111011110001",
28178 => "0011111011110100",
28179 => "0011111011110111",
28180 => "0011111011111010",
28181 => "0011111011111101",
28182 => "0011111100000000",
28183 => "0011111100000011",
28184 => "0011111100000110",
28185 => "0011111100001001",
28186 => "0011111100001100",
28187 => "0011111100001111",
28188 => "0011111100010010",
28189 => "0011111100010101",
28190 => "0011111100011000",
28191 => "0011111100011011",
28192 => "0011111100011110",
28193 => "0011111100100001",
28194 => "0011111100100100",
28195 => "0011111100100111",
28196 => "0011111100101001",
28197 => "0011111100101100",
28198 => "0011111100101111",
28199 => "0011111100110010",
28200 => "0011111100110101",
28201 => "0011111100111000",
28202 => "0011111100111011",
28203 => "0011111100111110",
28204 => "0011111101000001",
28205 => "0011111101000100",
28206 => "0011111101000111",
28207 => "0011111101001010",
28208 => "0011111101001101",
28209 => "0011111101010000",
28210 => "0011111101010011",
28211 => "0011111101010110",
28212 => "0011111101011001",
28213 => "0011111101011100",
28214 => "0011111101011111",
28215 => "0011111101100010",
28216 => "0011111101100101",
28217 => "0011111101101000",
28218 => "0011111101101011",
28219 => "0011111101101110",
28220 => "0011111101110001",
28221 => "0011111101110100",
28222 => "0011111101110111",
28223 => "0011111101111010",
28224 => "0011111101111101",
28225 => "0011111110000000",
28226 => "0011111110000011",
28227 => "0011111110000110",
28228 => "0011111110001001",
28229 => "0011111110001100",
28230 => "0011111110001111",
28231 => "0011111110010010",
28232 => "0011111110010101",
28233 => "0011111110011000",
28234 => "0011111110011011",
28235 => "0011111110011110",
28236 => "0011111110100001",
28237 => "0011111110100100",
28238 => "0011111110100111",
28239 => "0011111110101010",
28240 => "0011111110101101",
28241 => "0011111110110000",
28242 => "0011111110110011",
28243 => "0011111110110110",
28244 => "0011111110111001",
28245 => "0011111110111100",
28246 => "0011111110111111",
28247 => "0011111111000010",
28248 => "0011111111000101",
28249 => "0011111111001000",
28250 => "0011111111001011",
28251 => "0011111111001110",
28252 => "0011111111010001",
28253 => "0011111111010100",
28254 => "0011111111010111",
28255 => "0011111111011010",
28256 => "0011111111011101",
28257 => "0011111111100000",
28258 => "0011111111100011",
28259 => "0011111111100110",
28260 => "0011111111101001",
28261 => "0011111111101100",
28262 => "0011111111101111",
28263 => "0011111111110010",
28264 => "0011111111110101",
28265 => "0011111111111000",
28266 => "0011111111111011",
28267 => "0011111111111110",
28268 => "0100000000000001",
28269 => "0100000000000100",
28270 => "0100000000000111",
28271 => "0100000000001010",
28272 => "0100000000001101",
28273 => "0100000000010000",
28274 => "0100000000010011",
28275 => "0100000000010110",
28276 => "0100000000011001",
28277 => "0100000000011100",
28278 => "0100000000011111",
28279 => "0100000000100010",
28280 => "0100000000100101",
28281 => "0100000000101000",
28282 => "0100000000101011",
28283 => "0100000000101110",
28284 => "0100000000110001",
28285 => "0100000000110100",
28286 => "0100000000110111",
28287 => "0100000000111010",
28288 => "0100000000111101",
28289 => "0100000001000000",
28290 => "0100000001000011",
28291 => "0100000001000110",
28292 => "0100000001001001",
28293 => "0100000001001100",
28294 => "0100000001001111",
28295 => "0100000001010010",
28296 => "0100000001010101",
28297 => "0100000001011000",
28298 => "0100000001011011",
28299 => "0100000001011110",
28300 => "0100000001100001",
28301 => "0100000001100100",
28302 => "0100000001100111",
28303 => "0100000001101010",
28304 => "0100000001101101",
28305 => "0100000001110000",
28306 => "0100000001110011",
28307 => "0100000001110110",
28308 => "0100000001111001",
28309 => "0100000001111100",
28310 => "0100000001111111",
28311 => "0100000010000010",
28312 => "0100000010000101",
28313 => "0100000010001000",
28314 => "0100000010001011",
28315 => "0100000010001110",
28316 => "0100000010010001",
28317 => "0100000010010100",
28318 => "0100000010010111",
28319 => "0100000010011010",
28320 => "0100000010011101",
28321 => "0100000010100000",
28322 => "0100000010100011",
28323 => "0100000010100110",
28324 => "0100000010101001",
28325 => "0100000010101100",
28326 => "0100000010101111",
28327 => "0100000010110010",
28328 => "0100000010110101",
28329 => "0100000010111000",
28330 => "0100000010111011",
28331 => "0100000010111110",
28332 => "0100000011000001",
28333 => "0100000011000100",
28334 => "0100000011000111",
28335 => "0100000011001010",
28336 => "0100000011001101",
28337 => "0100000011010000",
28338 => "0100000011010011",
28339 => "0100000011010110",
28340 => "0100000011011010",
28341 => "0100000011011101",
28342 => "0100000011100000",
28343 => "0100000011100011",
28344 => "0100000011100110",
28345 => "0100000011101001",
28346 => "0100000011101100",
28347 => "0100000011101111",
28348 => "0100000011110010",
28349 => "0100000011110101",
28350 => "0100000011111000",
28351 => "0100000011111011",
28352 => "0100000011111110",
28353 => "0100000100000001",
28354 => "0100000100000100",
28355 => "0100000100000111",
28356 => "0100000100001010",
28357 => "0100000100001101",
28358 => "0100000100010000",
28359 => "0100000100010011",
28360 => "0100000100010110",
28361 => "0100000100011001",
28362 => "0100000100011100",
28363 => "0100000100011111",
28364 => "0100000100100010",
28365 => "0100000100100101",
28366 => "0100000100101000",
28367 => "0100000100101011",
28368 => "0100000100101110",
28369 => "0100000100110001",
28370 => "0100000100110100",
28371 => "0100000100110111",
28372 => "0100000100111011",
28373 => "0100000100111110",
28374 => "0100000101000001",
28375 => "0100000101000100",
28376 => "0100000101000111",
28377 => "0100000101001010",
28378 => "0100000101001101",
28379 => "0100000101010000",
28380 => "0100000101010011",
28381 => "0100000101010110",
28382 => "0100000101011001",
28383 => "0100000101011100",
28384 => "0100000101011111",
28385 => "0100000101100010",
28386 => "0100000101100101",
28387 => "0100000101101000",
28388 => "0100000101101011",
28389 => "0100000101101110",
28390 => "0100000101110001",
28391 => "0100000101110100",
28392 => "0100000101110111",
28393 => "0100000101111010",
28394 => "0100000101111101",
28395 => "0100000110000001",
28396 => "0100000110000100",
28397 => "0100000110000111",
28398 => "0100000110001010",
28399 => "0100000110001101",
28400 => "0100000110010000",
28401 => "0100000110010011",
28402 => "0100000110010110",
28403 => "0100000110011001",
28404 => "0100000110011100",
28405 => "0100000110011111",
28406 => "0100000110100010",
28407 => "0100000110100101",
28408 => "0100000110101000",
28409 => "0100000110101011",
28410 => "0100000110101110",
28411 => "0100000110110001",
28412 => "0100000110110100",
28413 => "0100000110110111",
28414 => "0100000110111010",
28415 => "0100000110111110",
28416 => "0100000111000001",
28417 => "0100000111000100",
28418 => "0100000111000111",
28419 => "0100000111001010",
28420 => "0100000111001101",
28421 => "0100000111010000",
28422 => "0100000111010011",
28423 => "0100000111010110",
28424 => "0100000111011001",
28425 => "0100000111011100",
28426 => "0100000111011111",
28427 => "0100000111100010",
28428 => "0100000111100101",
28429 => "0100000111101000",
28430 => "0100000111101011",
28431 => "0100000111101110",
28432 => "0100000111110001",
28433 => "0100000111110101",
28434 => "0100000111111000",
28435 => "0100000111111011",
28436 => "0100000111111110",
28437 => "0100001000000001",
28438 => "0100001000000100",
28439 => "0100001000000111",
28440 => "0100001000001010",
28441 => "0100001000001101",
28442 => "0100001000010000",
28443 => "0100001000010011",
28444 => "0100001000010110",
28445 => "0100001000011001",
28446 => "0100001000011100",
28447 => "0100001000011111",
28448 => "0100001000100010",
28449 => "0100001000100110",
28450 => "0100001000101001",
28451 => "0100001000101100",
28452 => "0100001000101111",
28453 => "0100001000110010",
28454 => "0100001000110101",
28455 => "0100001000111000",
28456 => "0100001000111011",
28457 => "0100001000111110",
28458 => "0100001001000001",
28459 => "0100001001000100",
28460 => "0100001001000111",
28461 => "0100001001001010",
28462 => "0100001001001101",
28463 => "0100001001010001",
28464 => "0100001001010100",
28465 => "0100001001010111",
28466 => "0100001001011010",
28467 => "0100001001011101",
28468 => "0100001001100000",
28469 => "0100001001100011",
28470 => "0100001001100110",
28471 => "0100001001101001",
28472 => "0100001001101100",
28473 => "0100001001101111",
28474 => "0100001001110010",
28475 => "0100001001110101",
28476 => "0100001001111000",
28477 => "0100001001111100",
28478 => "0100001001111111",
28479 => "0100001010000010",
28480 => "0100001010000101",
28481 => "0100001010001000",
28482 => "0100001010001011",
28483 => "0100001010001110",
28484 => "0100001010010001",
28485 => "0100001010010100",
28486 => "0100001010010111",
28487 => "0100001010011010",
28488 => "0100001010011101",
28489 => "0100001010100000",
28490 => "0100001010100100",
28491 => "0100001010100111",
28492 => "0100001010101010",
28493 => "0100001010101101",
28494 => "0100001010110000",
28495 => "0100001010110011",
28496 => "0100001010110110",
28497 => "0100001010111001",
28498 => "0100001010111100",
28499 => "0100001010111111",
28500 => "0100001011000010",
28501 => "0100001011000101",
28502 => "0100001011001001",
28503 => "0100001011001100",
28504 => "0100001011001111",
28505 => "0100001011010010",
28506 => "0100001011010101",
28507 => "0100001011011000",
28508 => "0100001011011011",
28509 => "0100001011011110",
28510 => "0100001011100001",
28511 => "0100001011100100",
28512 => "0100001011100111",
28513 => "0100001011101011",
28514 => "0100001011101110",
28515 => "0100001011110001",
28516 => "0100001011110100",
28517 => "0100001011110111",
28518 => "0100001011111010",
28519 => "0100001011111101",
28520 => "0100001100000000",
28521 => "0100001100000011",
28522 => "0100001100000110",
28523 => "0100001100001001",
28524 => "0100001100001101",
28525 => "0100001100010000",
28526 => "0100001100010011",
28527 => "0100001100010110",
28528 => "0100001100011001",
28529 => "0100001100011100",
28530 => "0100001100011111",
28531 => "0100001100100010",
28532 => "0100001100100101",
28533 => "0100001100101000",
28534 => "0100001100101011",
28535 => "0100001100101111",
28536 => "0100001100110010",
28537 => "0100001100110101",
28538 => "0100001100111000",
28539 => "0100001100111011",
28540 => "0100001100111110",
28541 => "0100001101000001",
28542 => "0100001101000100",
28543 => "0100001101000111",
28544 => "0100001101001010",
28545 => "0100001101001110",
28546 => "0100001101010001",
28547 => "0100001101010100",
28548 => "0100001101010111",
28549 => "0100001101011010",
28550 => "0100001101011101",
28551 => "0100001101100000",
28552 => "0100001101100011",
28553 => "0100001101100110",
28554 => "0100001101101001",
28555 => "0100001101101101",
28556 => "0100001101110000",
28557 => "0100001101110011",
28558 => "0100001101110110",
28559 => "0100001101111001",
28560 => "0100001101111100",
28561 => "0100001101111111",
28562 => "0100001110000010",
28563 => "0100001110000101",
28564 => "0100001110001001",
28565 => "0100001110001100",
28566 => "0100001110001111",
28567 => "0100001110010010",
28568 => "0100001110010101",
28569 => "0100001110011000",
28570 => "0100001110011011",
28571 => "0100001110011110",
28572 => "0100001110100001",
28573 => "0100001110100101",
28574 => "0100001110101000",
28575 => "0100001110101011",
28576 => "0100001110101110",
28577 => "0100001110110001",
28578 => "0100001110110100",
28579 => "0100001110110111",
28580 => "0100001110111010",
28581 => "0100001110111101",
28582 => "0100001111000001",
28583 => "0100001111000100",
28584 => "0100001111000111",
28585 => "0100001111001010",
28586 => "0100001111001101",
28587 => "0100001111010000",
28588 => "0100001111010011",
28589 => "0100001111010110",
28590 => "0100001111011001",
28591 => "0100001111011101",
28592 => "0100001111100000",
28593 => "0100001111100011",
28594 => "0100001111100110",
28595 => "0100001111101001",
28596 => "0100001111101100",
28597 => "0100001111101111",
28598 => "0100001111110010",
28599 => "0100001111110110",
28600 => "0100001111111001",
28601 => "0100001111111100",
28602 => "0100001111111111",
28603 => "0100010000000010",
28604 => "0100010000000101",
28605 => "0100010000001000",
28606 => "0100010000001011",
28607 => "0100010000001110",
28608 => "0100010000010010",
28609 => "0100010000010101",
28610 => "0100010000011000",
28611 => "0100010000011011",
28612 => "0100010000011110",
28613 => "0100010000100001",
28614 => "0100010000100100",
28615 => "0100010000100111",
28616 => "0100010000101011",
28617 => "0100010000101110",
28618 => "0100010000110001",
28619 => "0100010000110100",
28620 => "0100010000110111",
28621 => "0100010000111010",
28622 => "0100010000111101",
28623 => "0100010001000000",
28624 => "0100010001000100",
28625 => "0100010001000111",
28626 => "0100010001001010",
28627 => "0100010001001101",
28628 => "0100010001010000",
28629 => "0100010001010011",
28630 => "0100010001010110",
28631 => "0100010001011010",
28632 => "0100010001011101",
28633 => "0100010001100000",
28634 => "0100010001100011",
28635 => "0100010001100110",
28636 => "0100010001101001",
28637 => "0100010001101100",
28638 => "0100010001101111",
28639 => "0100010001110011",
28640 => "0100010001110110",
28641 => "0100010001111001",
28642 => "0100010001111100",
28643 => "0100010001111111",
28644 => "0100010010000010",
28645 => "0100010010000101",
28646 => "0100010010001001",
28647 => "0100010010001100",
28648 => "0100010010001111",
28649 => "0100010010010010",
28650 => "0100010010010101",
28651 => "0100010010011000",
28652 => "0100010010011011",
28653 => "0100010010011111",
28654 => "0100010010100010",
28655 => "0100010010100101",
28656 => "0100010010101000",
28657 => "0100010010101011",
28658 => "0100010010101110",
28659 => "0100010010110001",
28660 => "0100010010110100",
28661 => "0100010010111000",
28662 => "0100010010111011",
28663 => "0100010010111110",
28664 => "0100010011000001",
28665 => "0100010011000100",
28666 => "0100010011000111",
28667 => "0100010011001010",
28668 => "0100010011001110",
28669 => "0100010011010001",
28670 => "0100010011010100",
28671 => "0100010011010111",
28672 => "0100010011011010",
28673 => "0100010011011101",
28674 => "0100010011100001",
28675 => "0100010011100100",
28676 => "0100010011100111",
28677 => "0100010011101010",
28678 => "0100010011101101",
28679 => "0100010011110000",
28680 => "0100010011110011",
28681 => "0100010011110111",
28682 => "0100010011111010",
28683 => "0100010011111101",
28684 => "0100010100000000",
28685 => "0100010100000011",
28686 => "0100010100000110",
28687 => "0100010100001001",
28688 => "0100010100001101",
28689 => "0100010100010000",
28690 => "0100010100010011",
28691 => "0100010100010110",
28692 => "0100010100011001",
28693 => "0100010100011100",
28694 => "0100010100100000",
28695 => "0100010100100011",
28696 => "0100010100100110",
28697 => "0100010100101001",
28698 => "0100010100101100",
28699 => "0100010100101111",
28700 => "0100010100110010",
28701 => "0100010100110110",
28702 => "0100010100111001",
28703 => "0100010100111100",
28704 => "0100010100111111",
28705 => "0100010101000010",
28706 => "0100010101000101",
28707 => "0100010101001001",
28708 => "0100010101001100",
28709 => "0100010101001111",
28710 => "0100010101010010",
28711 => "0100010101010101",
28712 => "0100010101011000",
28713 => "0100010101011100",
28714 => "0100010101011111",
28715 => "0100010101100010",
28716 => "0100010101100101",
28717 => "0100010101101000",
28718 => "0100010101101011",
28719 => "0100010101101110",
28720 => "0100010101110010",
28721 => "0100010101110101",
28722 => "0100010101111000",
28723 => "0100010101111011",
28724 => "0100010101111110",
28725 => "0100010110000001",
28726 => "0100010110000101",
28727 => "0100010110001000",
28728 => "0100010110001011",
28729 => "0100010110001110",
28730 => "0100010110010001",
28731 => "0100010110010100",
28732 => "0100010110011000",
28733 => "0100010110011011",
28734 => "0100010110011110",
28735 => "0100010110100001",
28736 => "0100010110100100",
28737 => "0100010110100111",
28738 => "0100010110101011",
28739 => "0100010110101110",
28740 => "0100010110110001",
28741 => "0100010110110100",
28742 => "0100010110110111",
28743 => "0100010110111010",
28744 => "0100010110111110",
28745 => "0100010111000001",
28746 => "0100010111000100",
28747 => "0100010111000111",
28748 => "0100010111001010",
28749 => "0100010111001110",
28750 => "0100010111010001",
28751 => "0100010111010100",
28752 => "0100010111010111",
28753 => "0100010111011010",
28754 => "0100010111011101",
28755 => "0100010111100001",
28756 => "0100010111100100",
28757 => "0100010111100111",
28758 => "0100010111101010",
28759 => "0100010111101101",
28760 => "0100010111110000",
28761 => "0100010111110100",
28762 => "0100010111110111",
28763 => "0100010111111010",
28764 => "0100010111111101",
28765 => "0100011000000000",
28766 => "0100011000000100",
28767 => "0100011000000111",
28768 => "0100011000001010",
28769 => "0100011000001101",
28770 => "0100011000010000",
28771 => "0100011000010011",
28772 => "0100011000010111",
28773 => "0100011000011010",
28774 => "0100011000011101",
28775 => "0100011000100000",
28776 => "0100011000100011",
28777 => "0100011000100111",
28778 => "0100011000101010",
28779 => "0100011000101101",
28780 => "0100011000110000",
28781 => "0100011000110011",
28782 => "0100011000110110",
28783 => "0100011000111010",
28784 => "0100011000111101",
28785 => "0100011001000000",
28786 => "0100011001000011",
28787 => "0100011001000110",
28788 => "0100011001001010",
28789 => "0100011001001101",
28790 => "0100011001010000",
28791 => "0100011001010011",
28792 => "0100011001010110",
28793 => "0100011001011001",
28794 => "0100011001011101",
28795 => "0100011001100000",
28796 => "0100011001100011",
28797 => "0100011001100110",
28798 => "0100011001101001",
28799 => "0100011001101101",
28800 => "0100011001110000",
28801 => "0100011001110011",
28802 => "0100011001110110",
28803 => "0100011001111001",
28804 => "0100011001111101",
28805 => "0100011010000000",
28806 => "0100011010000011",
28807 => "0100011010000110",
28808 => "0100011010001001",
28809 => "0100011010001101",
28810 => "0100011010010000",
28811 => "0100011010010011",
28812 => "0100011010010110",
28813 => "0100011010011001",
28814 => "0100011010011101",
28815 => "0100011010100000",
28816 => "0100011010100011",
28817 => "0100011010100110",
28818 => "0100011010101001",
28819 => "0100011010101100",
28820 => "0100011010110000",
28821 => "0100011010110011",
28822 => "0100011010110110",
28823 => "0100011010111001",
28824 => "0100011010111100",
28825 => "0100011011000000",
28826 => "0100011011000011",
28827 => "0100011011000110",
28828 => "0100011011001001",
28829 => "0100011011001100",
28830 => "0100011011010000",
28831 => "0100011011010011",
28832 => "0100011011010110",
28833 => "0100011011011001",
28834 => "0100011011011101",
28835 => "0100011011100000",
28836 => "0100011011100011",
28837 => "0100011011100110",
28838 => "0100011011101001",
28839 => "0100011011101101",
28840 => "0100011011110000",
28841 => "0100011011110011",
28842 => "0100011011110110",
28843 => "0100011011111001",
28844 => "0100011011111101",
28845 => "0100011100000000",
28846 => "0100011100000011",
28847 => "0100011100000110",
28848 => "0100011100001001",
28849 => "0100011100001101",
28850 => "0100011100010000",
28851 => "0100011100010011",
28852 => "0100011100010110",
28853 => "0100011100011001",
28854 => "0100011100011101",
28855 => "0100011100100000",
28856 => "0100011100100011",
28857 => "0100011100100110",
28858 => "0100011100101001",
28859 => "0100011100101101",
28860 => "0100011100110000",
28861 => "0100011100110011",
28862 => "0100011100110110",
28863 => "0100011100111010",
28864 => "0100011100111101",
28865 => "0100011101000000",
28866 => "0100011101000011",
28867 => "0100011101000110",
28868 => "0100011101001010",
28869 => "0100011101001101",
28870 => "0100011101010000",
28871 => "0100011101010011",
28872 => "0100011101010110",
28873 => "0100011101011010",
28874 => "0100011101011101",
28875 => "0100011101100000",
28876 => "0100011101100011",
28877 => "0100011101100111",
28878 => "0100011101101010",
28879 => "0100011101101101",
28880 => "0100011101110000",
28881 => "0100011101110011",
28882 => "0100011101110111",
28883 => "0100011101111010",
28884 => "0100011101111101",
28885 => "0100011110000000",
28886 => "0100011110000100",
28887 => "0100011110000111",
28888 => "0100011110001010",
28889 => "0100011110001101",
28890 => "0100011110010000",
28891 => "0100011110010100",
28892 => "0100011110010111",
28893 => "0100011110011010",
28894 => "0100011110011101",
28895 => "0100011110100001",
28896 => "0100011110100100",
28897 => "0100011110100111",
28898 => "0100011110101010",
28899 => "0100011110101101",
28900 => "0100011110110001",
28901 => "0100011110110100",
28902 => "0100011110110111",
28903 => "0100011110111010",
28904 => "0100011110111110",
28905 => "0100011111000001",
28906 => "0100011111000100",
28907 => "0100011111000111",
28908 => "0100011111001010",
28909 => "0100011111001110",
28910 => "0100011111010001",
28911 => "0100011111010100",
28912 => "0100011111010111",
28913 => "0100011111011011",
28914 => "0100011111011110",
28915 => "0100011111100001",
28916 => "0100011111100100",
28917 => "0100011111101000",
28918 => "0100011111101011",
28919 => "0100011111101110",
28920 => "0100011111110001",
28921 => "0100011111110100",
28922 => "0100011111111000",
28923 => "0100011111111011",
28924 => "0100011111111110",
28925 => "0100100000000001",
28926 => "0100100000000101",
28927 => "0100100000001000",
28928 => "0100100000001011",
28929 => "0100100000001110",
28930 => "0100100000010010",
28931 => "0100100000010101",
28932 => "0100100000011000",
28933 => "0100100000011011",
28934 => "0100100000011111",
28935 => "0100100000100010",
28936 => "0100100000100101",
28937 => "0100100000101000",
28938 => "0100100000101100",
28939 => "0100100000101111",
28940 => "0100100000110010",
28941 => "0100100000110101",
28942 => "0100100000111000",
28943 => "0100100000111100",
28944 => "0100100000111111",
28945 => "0100100001000010",
28946 => "0100100001000101",
28947 => "0100100001001001",
28948 => "0100100001001100",
28949 => "0100100001001111",
28950 => "0100100001010010",
28951 => "0100100001010110",
28952 => "0100100001011001",
28953 => "0100100001011100",
28954 => "0100100001011111",
28955 => "0100100001100011",
28956 => "0100100001100110",
28957 => "0100100001101001",
28958 => "0100100001101100",
28959 => "0100100001110000",
28960 => "0100100001110011",
28961 => "0100100001110110",
28962 => "0100100001111001",
28963 => "0100100001111101",
28964 => "0100100010000000",
28965 => "0100100010000011",
28966 => "0100100010000110",
28967 => "0100100010001010",
28968 => "0100100010001101",
28969 => "0100100010010000",
28970 => "0100100010010011",
28971 => "0100100010010111",
28972 => "0100100010011010",
28973 => "0100100010011101",
28974 => "0100100010100000",
28975 => "0100100010100100",
28976 => "0100100010100111",
28977 => "0100100010101010",
28978 => "0100100010101101",
28979 => "0100100010110001",
28980 => "0100100010110100",
28981 => "0100100010110111",
28982 => "0100100010111010",
28983 => "0100100010111110",
28984 => "0100100011000001",
28985 => "0100100011000100",
28986 => "0100100011000111",
28987 => "0100100011001011",
28988 => "0100100011001110",
28989 => "0100100011010001",
28990 => "0100100011010100",
28991 => "0100100011011000",
28992 => "0100100011011011",
28993 => "0100100011011110",
28994 => "0100100011100001",
28995 => "0100100011100101",
28996 => "0100100011101000",
28997 => "0100100011101011",
28998 => "0100100011101110",
28999 => "0100100011110010",
29000 => "0100100011110101",
29001 => "0100100011111000",
29002 => "0100100011111100",
29003 => "0100100011111111",
29004 => "0100100100000010",
29005 => "0100100100000101",
29006 => "0100100100001001",
29007 => "0100100100001100",
29008 => "0100100100001111",
29009 => "0100100100010010",
29010 => "0100100100010110",
29011 => "0100100100011001",
29012 => "0100100100011100",
29013 => "0100100100011111",
29014 => "0100100100100011",
29015 => "0100100100100110",
29016 => "0100100100101001",
29017 => "0100100100101100",
29018 => "0100100100110000",
29019 => "0100100100110011",
29020 => "0100100100110110",
29021 => "0100100100111010",
29022 => "0100100100111101",
29023 => "0100100101000000",
29024 => "0100100101000011",
29025 => "0100100101000111",
29026 => "0100100101001010",
29027 => "0100100101001101",
29028 => "0100100101010000",
29029 => "0100100101010100",
29030 => "0100100101010111",
29031 => "0100100101011010",
29032 => "0100100101011101",
29033 => "0100100101100001",
29034 => "0100100101100100",
29035 => "0100100101100111",
29036 => "0100100101101011",
29037 => "0100100101101110",
29038 => "0100100101110001",
29039 => "0100100101110100",
29040 => "0100100101111000",
29041 => "0100100101111011",
29042 => "0100100101111110",
29043 => "0100100110000010",
29044 => "0100100110000101",
29045 => "0100100110001000",
29046 => "0100100110001011",
29047 => "0100100110001111",
29048 => "0100100110010010",
29049 => "0100100110010101",
29050 => "0100100110011000",
29051 => "0100100110011100",
29052 => "0100100110011111",
29053 => "0100100110100010",
29054 => "0100100110100110",
29055 => "0100100110101001",
29056 => "0100100110101100",
29057 => "0100100110101111",
29058 => "0100100110110011",
29059 => "0100100110110110",
29060 => "0100100110111001",
29061 => "0100100110111101",
29062 => "0100100111000000",
29063 => "0100100111000011",
29064 => "0100100111000110",
29065 => "0100100111001010",
29066 => "0100100111001101",
29067 => "0100100111010000",
29068 => "0100100111010011",
29069 => "0100100111010111",
29070 => "0100100111011010",
29071 => "0100100111011101",
29072 => "0100100111100001",
29073 => "0100100111100100",
29074 => "0100100111100111",
29075 => "0100100111101010",
29076 => "0100100111101110",
29077 => "0100100111110001",
29078 => "0100100111110100",
29079 => "0100100111111000",
29080 => "0100100111111011",
29081 => "0100100111111110",
29082 => "0100101000000001",
29083 => "0100101000000101",
29084 => "0100101000001000",
29085 => "0100101000001011",
29086 => "0100101000001111",
29087 => "0100101000010010",
29088 => "0100101000010101",
29089 => "0100101000011001",
29090 => "0100101000011100",
29091 => "0100101000011111",
29092 => "0100101000100010",
29093 => "0100101000100110",
29094 => "0100101000101001",
29095 => "0100101000101100",
29096 => "0100101000110000",
29097 => "0100101000110011",
29098 => "0100101000110110",
29099 => "0100101000111001",
29100 => "0100101000111101",
29101 => "0100101001000000",
29102 => "0100101001000011",
29103 => "0100101001000111",
29104 => "0100101001001010",
29105 => "0100101001001101",
29106 => "0100101001010001",
29107 => "0100101001010100",
29108 => "0100101001010111",
29109 => "0100101001011010",
29110 => "0100101001011110",
29111 => "0100101001100001",
29112 => "0100101001100100",
29113 => "0100101001101000",
29114 => "0100101001101011",
29115 => "0100101001101110",
29116 => "0100101001110001",
29117 => "0100101001110101",
29118 => "0100101001111000",
29119 => "0100101001111011",
29120 => "0100101001111111",
29121 => "0100101010000010",
29122 => "0100101010000101",
29123 => "0100101010001001",
29124 => "0100101010001100",
29125 => "0100101010001111",
29126 => "0100101010010011",
29127 => "0100101010010110",
29128 => "0100101010011001",
29129 => "0100101010011100",
29130 => "0100101010100000",
29131 => "0100101010100011",
29132 => "0100101010100110",
29133 => "0100101010101010",
29134 => "0100101010101101",
29135 => "0100101010110000",
29136 => "0100101010110100",
29137 => "0100101010110111",
29138 => "0100101010111010",
29139 => "0100101010111101",
29140 => "0100101011000001",
29141 => "0100101011000100",
29142 => "0100101011000111",
29143 => "0100101011001011",
29144 => "0100101011001110",
29145 => "0100101011010001",
29146 => "0100101011010101",
29147 => "0100101011011000",
29148 => "0100101011011011",
29149 => "0100101011011111",
29150 => "0100101011100010",
29151 => "0100101011100101",
29152 => "0100101011101000",
29153 => "0100101011101100",
29154 => "0100101011101111",
29155 => "0100101011110010",
29156 => "0100101011110110",
29157 => "0100101011111001",
29158 => "0100101011111100",
29159 => "0100101100000000",
29160 => "0100101100000011",
29161 => "0100101100000110",
29162 => "0100101100001010",
29163 => "0100101100001101",
29164 => "0100101100010000",
29165 => "0100101100010100",
29166 => "0100101100010111",
29167 => "0100101100011010",
29168 => "0100101100011110",
29169 => "0100101100100001",
29170 => "0100101100100100",
29171 => "0100101100100111",
29172 => "0100101100101011",
29173 => "0100101100101110",
29174 => "0100101100110001",
29175 => "0100101100110101",
29176 => "0100101100111000",
29177 => "0100101100111011",
29178 => "0100101100111111",
29179 => "0100101101000010",
29180 => "0100101101000101",
29181 => "0100101101001001",
29182 => "0100101101001100",
29183 => "0100101101001111",
29184 => "0100101101010011",
29185 => "0100101101010110",
29186 => "0100101101011001",
29187 => "0100101101011101",
29188 => "0100101101100000",
29189 => "0100101101100011",
29190 => "0100101101100111",
29191 => "0100101101101010",
29192 => "0100101101101101",
29193 => "0100101101110001",
29194 => "0100101101110100",
29195 => "0100101101110111",
29196 => "0100101101111011",
29197 => "0100101101111110",
29198 => "0100101110000001",
29199 => "0100101110000101",
29200 => "0100101110001000",
29201 => "0100101110001011",
29202 => "0100101110001111",
29203 => "0100101110010010",
29204 => "0100101110010101",
29205 => "0100101110011001",
29206 => "0100101110011100",
29207 => "0100101110011111",
29208 => "0100101110100010",
29209 => "0100101110100110",
29210 => "0100101110101001",
29211 => "0100101110101100",
29212 => "0100101110110000",
29213 => "0100101110110011",
29214 => "0100101110110110",
29215 => "0100101110111010",
29216 => "0100101110111101",
29217 => "0100101111000000",
29218 => "0100101111000100",
29219 => "0100101111000111",
29220 => "0100101111001010",
29221 => "0100101111001110",
29222 => "0100101111010001",
29223 => "0100101111010100",
29224 => "0100101111011000",
29225 => "0100101111011011",
29226 => "0100101111011110",
29227 => "0100101111100010",
29228 => "0100101111100101",
29229 => "0100101111101001",
29230 => "0100101111101100",
29231 => "0100101111101111",
29232 => "0100101111110011",
29233 => "0100101111110110",
29234 => "0100101111111001",
29235 => "0100101111111101",
29236 => "0100110000000000",
29237 => "0100110000000011",
29238 => "0100110000000111",
29239 => "0100110000001010",
29240 => "0100110000001101",
29241 => "0100110000010001",
29242 => "0100110000010100",
29243 => "0100110000010111",
29244 => "0100110000011011",
29245 => "0100110000011110",
29246 => "0100110000100001",
29247 => "0100110000100101",
29248 => "0100110000101000",
29249 => "0100110000101011",
29250 => "0100110000101111",
29251 => "0100110000110010",
29252 => "0100110000110101",
29253 => "0100110000111001",
29254 => "0100110000111100",
29255 => "0100110000111111",
29256 => "0100110001000011",
29257 => "0100110001000110",
29258 => "0100110001001001",
29259 => "0100110001001101",
29260 => "0100110001010000",
29261 => "0100110001010011",
29262 => "0100110001010111",
29263 => "0100110001011010",
29264 => "0100110001011110",
29265 => "0100110001100001",
29266 => "0100110001100100",
29267 => "0100110001101000",
29268 => "0100110001101011",
29269 => "0100110001101110",
29270 => "0100110001110010",
29271 => "0100110001110101",
29272 => "0100110001111000",
29273 => "0100110001111100",
29274 => "0100110001111111",
29275 => "0100110010000010",
29276 => "0100110010000110",
29277 => "0100110010001001",
29278 => "0100110010001100",
29279 => "0100110010010000",
29280 => "0100110010010011",
29281 => "0100110010010111",
29282 => "0100110010011010",
29283 => "0100110010011101",
29284 => "0100110010100001",
29285 => "0100110010100100",
29286 => "0100110010100111",
29287 => "0100110010101011",
29288 => "0100110010101110",
29289 => "0100110010110001",
29290 => "0100110010110101",
29291 => "0100110010111000",
29292 => "0100110010111011",
29293 => "0100110010111111",
29294 => "0100110011000010",
29295 => "0100110011000110",
29296 => "0100110011001001",
29297 => "0100110011001100",
29298 => "0100110011010000",
29299 => "0100110011010011",
29300 => "0100110011010110",
29301 => "0100110011011010",
29302 => "0100110011011101",
29303 => "0100110011100000",
29304 => "0100110011100100",
29305 => "0100110011100111",
29306 => "0100110011101010",
29307 => "0100110011101110",
29308 => "0100110011110001",
29309 => "0100110011110101",
29310 => "0100110011111000",
29311 => "0100110011111011",
29312 => "0100110011111111",
29313 => "0100110100000010",
29314 => "0100110100000101",
29315 => "0100110100001001",
29316 => "0100110100001100",
29317 => "0100110100001111",
29318 => "0100110100010011",
29319 => "0100110100010110",
29320 => "0100110100011010",
29321 => "0100110100011101",
29322 => "0100110100100000",
29323 => "0100110100100100",
29324 => "0100110100100111",
29325 => "0100110100101010",
29326 => "0100110100101110",
29327 => "0100110100110001",
29328 => "0100110100110101",
29329 => "0100110100111000",
29330 => "0100110100111011",
29331 => "0100110100111111",
29332 => "0100110101000010",
29333 => "0100110101000101",
29334 => "0100110101001001",
29335 => "0100110101001100",
29336 => "0100110101010000",
29337 => "0100110101010011",
29338 => "0100110101010110",
29339 => "0100110101011010",
29340 => "0100110101011101",
29341 => "0100110101100000",
29342 => "0100110101100100",
29343 => "0100110101100111",
29344 => "0100110101101011",
29345 => "0100110101101110",
29346 => "0100110101110001",
29347 => "0100110101110101",
29348 => "0100110101111000",
29349 => "0100110101111011",
29350 => "0100110101111111",
29351 => "0100110110000010",
29352 => "0100110110000110",
29353 => "0100110110001001",
29354 => "0100110110001100",
29355 => "0100110110010000",
29356 => "0100110110010011",
29357 => "0100110110010110",
29358 => "0100110110011010",
29359 => "0100110110011101",
29360 => "0100110110100001",
29361 => "0100110110100100",
29362 => "0100110110100111",
29363 => "0100110110101011",
29364 => "0100110110101110",
29365 => "0100110110110001",
29366 => "0100110110110101",
29367 => "0100110110111000",
29368 => "0100110110111100",
29369 => "0100110110111111",
29370 => "0100110111000010",
29371 => "0100110111000110",
29372 => "0100110111001001",
29373 => "0100110111001101",
29374 => "0100110111010000",
29375 => "0100110111010011",
29376 => "0100110111010111",
29377 => "0100110111011010",
29378 => "0100110111011101",
29379 => "0100110111100001",
29380 => "0100110111100100",
29381 => "0100110111101000",
29382 => "0100110111101011",
29383 => "0100110111101110",
29384 => "0100110111110010",
29385 => "0100110111110101",
29386 => "0100110111111001",
29387 => "0100110111111100",
29388 => "0100110111111111",
29389 => "0100111000000011",
29390 => "0100111000000110",
29391 => "0100111000001010",
29392 => "0100111000001101",
29393 => "0100111000010000",
29394 => "0100111000010100",
29395 => "0100111000010111",
29396 => "0100111000011010",
29397 => "0100111000011110",
29398 => "0100111000100001",
29399 => "0100111000100101",
29400 => "0100111000101000",
29401 => "0100111000101011",
29402 => "0100111000101111",
29403 => "0100111000110010",
29404 => "0100111000110110",
29405 => "0100111000111001",
29406 => "0100111000111100",
29407 => "0100111001000000",
29408 => "0100111001000011",
29409 => "0100111001000111",
29410 => "0100111001001010",
29411 => "0100111001001101",
29412 => "0100111001010001",
29413 => "0100111001010100",
29414 => "0100111001011000",
29415 => "0100111001011011",
29416 => "0100111001011110",
29417 => "0100111001100010",
29418 => "0100111001100101",
29419 => "0100111001101001",
29420 => "0100111001101100",
29421 => "0100111001101111",
29422 => "0100111001110011",
29423 => "0100111001110110",
29424 => "0100111001111010",
29425 => "0100111001111101",
29426 => "0100111010000000",
29427 => "0100111010000100",
29428 => "0100111010000111",
29429 => "0100111010001011",
29430 => "0100111010001110",
29431 => "0100111010010001",
29432 => "0100111010010101",
29433 => "0100111010011000",
29434 => "0100111010011100",
29435 => "0100111010011111",
29436 => "0100111010100010",
29437 => "0100111010100110",
29438 => "0100111010101001",
29439 => "0100111010101101",
29440 => "0100111010110000",
29441 => "0100111010110011",
29442 => "0100111010110111",
29443 => "0100111010111010",
29444 => "0100111010111110",
29445 => "0100111011000001",
29446 => "0100111011000100",
29447 => "0100111011001000",
29448 => "0100111011001011",
29449 => "0100111011001111",
29450 => "0100111011010010",
29451 => "0100111011010110",
29452 => "0100111011011001",
29453 => "0100111011011100",
29454 => "0100111011100000",
29455 => "0100111011100011",
29456 => "0100111011100111",
29457 => "0100111011101010",
29458 => "0100111011101101",
29459 => "0100111011110001",
29460 => "0100111011110100",
29461 => "0100111011111000",
29462 => "0100111011111011",
29463 => "0100111011111110",
29464 => "0100111100000010",
29465 => "0100111100000101",
29466 => "0100111100001001",
29467 => "0100111100001100",
29468 => "0100111100010000",
29469 => "0100111100010011",
29470 => "0100111100010110",
29471 => "0100111100011010",
29472 => "0100111100011101",
29473 => "0100111100100001",
29474 => "0100111100100100",
29475 => "0100111100100111",
29476 => "0100111100101011",
29477 => "0100111100101110",
29478 => "0100111100110010",
29479 => "0100111100110101",
29480 => "0100111100111001",
29481 => "0100111100111100",
29482 => "0100111100111111",
29483 => "0100111101000011",
29484 => "0100111101000110",
29485 => "0100111101001010",
29486 => "0100111101001101",
29487 => "0100111101010000",
29488 => "0100111101010100",
29489 => "0100111101010111",
29490 => "0100111101011011",
29491 => "0100111101011110",
29492 => "0100111101100010",
29493 => "0100111101100101",
29494 => "0100111101101000",
29495 => "0100111101101100",
29496 => "0100111101101111",
29497 => "0100111101110011",
29498 => "0100111101110110",
29499 => "0100111101111010",
29500 => "0100111101111101",
29501 => "0100111110000000",
29502 => "0100111110000100",
29503 => "0100111110000111",
29504 => "0100111110001011",
29505 => "0100111110001110",
29506 => "0100111110010010",
29507 => "0100111110010101",
29508 => "0100111110011000",
29509 => "0100111110011100",
29510 => "0100111110011111",
29511 => "0100111110100011",
29512 => "0100111110100110",
29513 => "0100111110101010",
29514 => "0100111110101101",
29515 => "0100111110110000",
29516 => "0100111110110100",
29517 => "0100111110110111",
29518 => "0100111110111011",
29519 => "0100111110111110",
29520 => "0100111111000010",
29521 => "0100111111000101",
29522 => "0100111111001000",
29523 => "0100111111001100",
29524 => "0100111111001111",
29525 => "0100111111010011",
29526 => "0100111111010110",
29527 => "0100111111011010",
29528 => "0100111111011101",
29529 => "0100111111100000",
29530 => "0100111111100100",
29531 => "0100111111100111",
29532 => "0100111111101011",
29533 => "0100111111101110",
29534 => "0100111111110010",
29535 => "0100111111110101",
29536 => "0100111111111001",
29537 => "0100111111111100",
29538 => "0100111111111111",
29539 => "0101000000000011",
29540 => "0101000000000110",
29541 => "0101000000001010",
29542 => "0101000000001101",
29543 => "0101000000010001",
29544 => "0101000000010100",
29545 => "0101000000010111",
29546 => "0101000000011011",
29547 => "0101000000011110",
29548 => "0101000000100010",
29549 => "0101000000100101",
29550 => "0101000000101001",
29551 => "0101000000101100",
29552 => "0101000000110000",
29553 => "0101000000110011",
29554 => "0101000000110110",
29555 => "0101000000111010",
29556 => "0101000000111101",
29557 => "0101000001000001",
29558 => "0101000001000100",
29559 => "0101000001001000",
29560 => "0101000001001011",
29561 => "0101000001001111",
29562 => "0101000001010010",
29563 => "0101000001010101",
29564 => "0101000001011001",
29565 => "0101000001011100",
29566 => "0101000001100000",
29567 => "0101000001100011",
29568 => "0101000001100111",
29569 => "0101000001101010",
29570 => "0101000001101110",
29571 => "0101000001110001",
29572 => "0101000001110100",
29573 => "0101000001111000",
29574 => "0101000001111011",
29575 => "0101000001111111",
29576 => "0101000010000010",
29577 => "0101000010000110",
29578 => "0101000010001001",
29579 => "0101000010001101",
29580 => "0101000010010000",
29581 => "0101000010010100",
29582 => "0101000010010111",
29583 => "0101000010011010",
29584 => "0101000010011110",
29585 => "0101000010100001",
29586 => "0101000010100101",
29587 => "0101000010101000",
29588 => "0101000010101100",
29589 => "0101000010101111",
29590 => "0101000010110011",
29591 => "0101000010110110",
29592 => "0101000010111001",
29593 => "0101000010111101",
29594 => "0101000011000000",
29595 => "0101000011000100",
29596 => "0101000011000111",
29597 => "0101000011001011",
29598 => "0101000011001110",
29599 => "0101000011010010",
29600 => "0101000011010101",
29601 => "0101000011011001",
29602 => "0101000011011100",
29603 => "0101000011100000",
29604 => "0101000011100011",
29605 => "0101000011100110",
29606 => "0101000011101010",
29607 => "0101000011101101",
29608 => "0101000011110001",
29609 => "0101000011110100",
29610 => "0101000011111000",
29611 => "0101000011111011",
29612 => "0101000011111111",
29613 => "0101000100000010",
29614 => "0101000100000110",
29615 => "0101000100001001",
29616 => "0101000100001100",
29617 => "0101000100010000",
29618 => "0101000100010011",
29619 => "0101000100010111",
29620 => "0101000100011010",
29621 => "0101000100011110",
29622 => "0101000100100001",
29623 => "0101000100100101",
29624 => "0101000100101000",
29625 => "0101000100101100",
29626 => "0101000100101111",
29627 => "0101000100110011",
29628 => "0101000100110110",
29629 => "0101000100111010",
29630 => "0101000100111101",
29631 => "0101000101000000",
29632 => "0101000101000100",
29633 => "0101000101000111",
29634 => "0101000101001011",
29635 => "0101000101001110",
29636 => "0101000101010010",
29637 => "0101000101010101",
29638 => "0101000101011001",
29639 => "0101000101011100",
29640 => "0101000101100000",
29641 => "0101000101100011",
29642 => "0101000101100111",
29643 => "0101000101101010",
29644 => "0101000101101110",
29645 => "0101000101110001",
29646 => "0101000101110100",
29647 => "0101000101111000",
29648 => "0101000101111011",
29649 => "0101000101111111",
29650 => "0101000110000010",
29651 => "0101000110000110",
29652 => "0101000110001001",
29653 => "0101000110001101",
29654 => "0101000110010000",
29655 => "0101000110010100",
29656 => "0101000110010111",
29657 => "0101000110011011",
29658 => "0101000110011110",
29659 => "0101000110100010",
29660 => "0101000110100101",
29661 => "0101000110101001",
29662 => "0101000110101100",
29663 => "0101000110110000",
29664 => "0101000110110011",
29665 => "0101000110110110",
29666 => "0101000110111010",
29667 => "0101000110111101",
29668 => "0101000111000001",
29669 => "0101000111000100",
29670 => "0101000111001000",
29671 => "0101000111001011",
29672 => "0101000111001111",
29673 => "0101000111010010",
29674 => "0101000111010110",
29675 => "0101000111011001",
29676 => "0101000111011101",
29677 => "0101000111100000",
29678 => "0101000111100100",
29679 => "0101000111100111",
29680 => "0101000111101011",
29681 => "0101000111101110",
29682 => "0101000111110010",
29683 => "0101000111110101",
29684 => "0101000111111001",
29685 => "0101000111111100",
29686 => "0101001000000000",
29687 => "0101001000000011",
29688 => "0101001000000111",
29689 => "0101001000001010",
29690 => "0101001000001110",
29691 => "0101001000010001",
29692 => "0101001000010100",
29693 => "0101001000011000",
29694 => "0101001000011011",
29695 => "0101001000011111",
29696 => "0101001000100010",
29697 => "0101001000100110",
29698 => "0101001000101001",
29699 => "0101001000101101",
29700 => "0101001000110000",
29701 => "0101001000110100",
29702 => "0101001000110111",
29703 => "0101001000111011",
29704 => "0101001000111110",
29705 => "0101001001000010",
29706 => "0101001001000101",
29707 => "0101001001001001",
29708 => "0101001001001100",
29709 => "0101001001010000",
29710 => "0101001001010011",
29711 => "0101001001010111",
29712 => "0101001001011010",
29713 => "0101001001011110",
29714 => "0101001001100001",
29715 => "0101001001100101",
29716 => "0101001001101000",
29717 => "0101001001101100",
29718 => "0101001001101111",
29719 => "0101001001110011",
29720 => "0101001001110110",
29721 => "0101001001111010",
29722 => "0101001001111101",
29723 => "0101001010000001",
29724 => "0101001010000100",
29725 => "0101001010001000",
29726 => "0101001010001011",
29727 => "0101001010001111",
29728 => "0101001010010010",
29729 => "0101001010010110",
29730 => "0101001010011001",
29731 => "0101001010011101",
29732 => "0101001010100000",
29733 => "0101001010100100",
29734 => "0101001010100111",
29735 => "0101001010101011",
29736 => "0101001010101110",
29737 => "0101001010110010",
29738 => "0101001010110101",
29739 => "0101001010111001",
29740 => "0101001010111100",
29741 => "0101001011000000",
29742 => "0101001011000011",
29743 => "0101001011000111",
29744 => "0101001011001010",
29745 => "0101001011001110",
29746 => "0101001011010001",
29747 => "0101001011010101",
29748 => "0101001011011000",
29749 => "0101001011011100",
29750 => "0101001011011111",
29751 => "0101001011100011",
29752 => "0101001011100110",
29753 => "0101001011101010",
29754 => "0101001011101101",
29755 => "0101001011110001",
29756 => "0101001011110100",
29757 => "0101001011111000",
29758 => "0101001011111011",
29759 => "0101001011111111",
29760 => "0101001100000010",
29761 => "0101001100000110",
29762 => "0101001100001001",
29763 => "0101001100001101",
29764 => "0101001100010000",
29765 => "0101001100010100",
29766 => "0101001100010111",
29767 => "0101001100011011",
29768 => "0101001100011110",
29769 => "0101001100100010",
29770 => "0101001100100101",
29771 => "0101001100101001",
29772 => "0101001100101100",
29773 => "0101001100110000",
29774 => "0101001100110011",
29775 => "0101001100110111",
29776 => "0101001100111010",
29777 => "0101001100111110",
29778 => "0101001101000001",
29779 => "0101001101000101",
29780 => "0101001101001000",
29781 => "0101001101001100",
29782 => "0101001101001111",
29783 => "0101001101010011",
29784 => "0101001101010110",
29785 => "0101001101011010",
29786 => "0101001101011101",
29787 => "0101001101100001",
29788 => "0101001101100100",
29789 => "0101001101101000",
29790 => "0101001101101011",
29791 => "0101001101101111",
29792 => "0101001101110011",
29793 => "0101001101110110",
29794 => "0101001101111010",
29795 => "0101001101111101",
29796 => "0101001110000001",
29797 => "0101001110000100",
29798 => "0101001110001000",
29799 => "0101001110001011",
29800 => "0101001110001111",
29801 => "0101001110010010",
29802 => "0101001110010110",
29803 => "0101001110011001",
29804 => "0101001110011101",
29805 => "0101001110100000",
29806 => "0101001110100100",
29807 => "0101001110100111",
29808 => "0101001110101011",
29809 => "0101001110101110",
29810 => "0101001110110010",
29811 => "0101001110110101",
29812 => "0101001110111001",
29813 => "0101001110111100",
29814 => "0101001111000000",
29815 => "0101001111000011",
29816 => "0101001111000111",
29817 => "0101001111001011",
29818 => "0101001111001110",
29819 => "0101001111010010",
29820 => "0101001111010101",
29821 => "0101001111011001",
29822 => "0101001111011100",
29823 => "0101001111100000",
29824 => "0101001111100011",
29825 => "0101001111100111",
29826 => "0101001111101010",
29827 => "0101001111101110",
29828 => "0101001111110001",
29829 => "0101001111110101",
29830 => "0101001111111000",
29831 => "0101001111111100",
29832 => "0101001111111111",
29833 => "0101010000000011",
29834 => "0101010000000110",
29835 => "0101010000001010",
29836 => "0101010000001101",
29837 => "0101010000010001",
29838 => "0101010000010101",
29839 => "0101010000011000",
29840 => "0101010000011100",
29841 => "0101010000011111",
29842 => "0101010000100011",
29843 => "0101010000100110",
29844 => "0101010000101010",
29845 => "0101010000101101",
29846 => "0101010000110001",
29847 => "0101010000110100",
29848 => "0101010000111000",
29849 => "0101010000111011",
29850 => "0101010000111111",
29851 => "0101010001000010",
29852 => "0101010001000110",
29853 => "0101010001001010",
29854 => "0101010001001101",
29855 => "0101010001010001",
29856 => "0101010001010100",
29857 => "0101010001011000",
29858 => "0101010001011011",
29859 => "0101010001011111",
29860 => "0101010001100010",
29861 => "0101010001100110",
29862 => "0101010001101001",
29863 => "0101010001101101",
29864 => "0101010001110000",
29865 => "0101010001110100",
29866 => "0101010001110111",
29867 => "0101010001111011",
29868 => "0101010001111111",
29869 => "0101010010000010",
29870 => "0101010010000110",
29871 => "0101010010001001",
29872 => "0101010010001101",
29873 => "0101010010010000",
29874 => "0101010010010100",
29875 => "0101010010010111",
29876 => "0101010010011011",
29877 => "0101010010011110",
29878 => "0101010010100010",
29879 => "0101010010100101",
29880 => "0101010010101001",
29881 => "0101010010101101",
29882 => "0101010010110000",
29883 => "0101010010110100",
29884 => "0101010010110111",
29885 => "0101010010111011",
29886 => "0101010010111110",
29887 => "0101010011000010",
29888 => "0101010011000101",
29889 => "0101010011001001",
29890 => "0101010011001100",
29891 => "0101010011010000",
29892 => "0101010011010100",
29893 => "0101010011010111",
29894 => "0101010011011011",
29895 => "0101010011011110",
29896 => "0101010011100010",
29897 => "0101010011100101",
29898 => "0101010011101001",
29899 => "0101010011101100",
29900 => "0101010011110000",
29901 => "0101010011110011",
29902 => "0101010011110111",
29903 => "0101010011111011",
29904 => "0101010011111110",
29905 => "0101010100000010",
29906 => "0101010100000101",
29907 => "0101010100001001",
29908 => "0101010100001100",
29909 => "0101010100010000",
29910 => "0101010100010011",
29911 => "0101010100010111",
29912 => "0101010100011011",
29913 => "0101010100011110",
29914 => "0101010100100010",
29915 => "0101010100100101",
29916 => "0101010100101001",
29917 => "0101010100101100",
29918 => "0101010100110000",
29919 => "0101010100110011",
29920 => "0101010100110111",
29921 => "0101010100111010",
29922 => "0101010100111110",
29923 => "0101010101000010",
29924 => "0101010101000101",
29925 => "0101010101001001",
29926 => "0101010101001100",
29927 => "0101010101010000",
29928 => "0101010101010011",
29929 => "0101010101010111",
29930 => "0101010101011010",
29931 => "0101010101011110",
29932 => "0101010101100010",
29933 => "0101010101100101",
29934 => "0101010101101001",
29935 => "0101010101101100",
29936 => "0101010101110000",
29937 => "0101010101110011",
29938 => "0101010101110111",
29939 => "0101010101111010",
29940 => "0101010101111110",
29941 => "0101010110000010",
29942 => "0101010110000101",
29943 => "0101010110001001",
29944 => "0101010110001100",
29945 => "0101010110010000",
29946 => "0101010110010011",
29947 => "0101010110010111",
29948 => "0101010110011011",
29949 => "0101010110011110",
29950 => "0101010110100010",
29951 => "0101010110100101",
29952 => "0101010110101001",
29953 => "0101010110101100",
29954 => "0101010110110000",
29955 => "0101010110110011",
29956 => "0101010110110111",
29957 => "0101010110111011",
29958 => "0101010110111110",
29959 => "0101010111000010",
29960 => "0101010111000101",
29961 => "0101010111001001",
29962 => "0101010111001100",
29963 => "0101010111010000",
29964 => "0101010111010100",
29965 => "0101010111010111",
29966 => "0101010111011011",
29967 => "0101010111011110",
29968 => "0101010111100010",
29969 => "0101010111100101",
29970 => "0101010111101001",
29971 => "0101010111101101",
29972 => "0101010111110000",
29973 => "0101010111110100",
29974 => "0101010111110111",
29975 => "0101010111111011",
29976 => "0101010111111110",
29977 => "0101011000000010",
29978 => "0101011000000110",
29979 => "0101011000001001",
29980 => "0101011000001101",
29981 => "0101011000010000",
29982 => "0101011000010100",
29983 => "0101011000010111",
29984 => "0101011000011011",
29985 => "0101011000011110",
29986 => "0101011000100010",
29987 => "0101011000100110",
29988 => "0101011000101001",
29989 => "0101011000101101",
29990 => "0101011000110000",
29991 => "0101011000110100",
29992 => "0101011000111000",
29993 => "0101011000111011",
29994 => "0101011000111111",
29995 => "0101011001000010",
29996 => "0101011001000110",
29997 => "0101011001001001",
29998 => "0101011001001101",
29999 => "0101011001010001",
30000 => "0101011001010100",
30001 => "0101011001011000",
30002 => "0101011001011011",
30003 => "0101011001011111",
30004 => "0101011001100010",
30005 => "0101011001100110",
30006 => "0101011001101010",
30007 => "0101011001101101",
30008 => "0101011001110001",
30009 => "0101011001110100",
30010 => "0101011001111000",
30011 => "0101011001111011",
30012 => "0101011001111111",
30013 => "0101011010000011",
30014 => "0101011010000110",
30015 => "0101011010001010",
30016 => "0101011010001101",
30017 => "0101011010010001",
30018 => "0101011010010101",
30019 => "0101011010011000",
30020 => "0101011010011100",
30021 => "0101011010011111",
30022 => "0101011010100011",
30023 => "0101011010100110",
30024 => "0101011010101010",
30025 => "0101011010101110",
30026 => "0101011010110001",
30027 => "0101011010110101",
30028 => "0101011010111000",
30029 => "0101011010111100",
30030 => "0101011011000000",
30031 => "0101011011000011",
30032 => "0101011011000111",
30033 => "0101011011001010",
30034 => "0101011011001110",
30035 => "0101011011010001",
30036 => "0101011011010101",
30037 => "0101011011011001",
30038 => "0101011011011100",
30039 => "0101011011100000",
30040 => "0101011011100011",
30041 => "0101011011100111",
30042 => "0101011011101011",
30043 => "0101011011101110",
30044 => "0101011011110010",
30045 => "0101011011110101",
30046 => "0101011011111001",
30047 => "0101011011111100",
30048 => "0101011100000000",
30049 => "0101011100000100",
30050 => "0101011100000111",
30051 => "0101011100001011",
30052 => "0101011100001110",
30053 => "0101011100010010",
30054 => "0101011100010110",
30055 => "0101011100011001",
30056 => "0101011100011101",
30057 => "0101011100100000",
30058 => "0101011100100100",
30059 => "0101011100101000",
30060 => "0101011100101011",
30061 => "0101011100101111",
30062 => "0101011100110010",
30063 => "0101011100110110",
30064 => "0101011100111010",
30065 => "0101011100111101",
30066 => "0101011101000001",
30067 => "0101011101000100",
30068 => "0101011101001000",
30069 => "0101011101001100",
30070 => "0101011101001111",
30071 => "0101011101010011",
30072 => "0101011101010110",
30073 => "0101011101011010",
30074 => "0101011101011110",
30075 => "0101011101100001",
30076 => "0101011101100101",
30077 => "0101011101101000",
30078 => "0101011101101100",
30079 => "0101011101110000",
30080 => "0101011101110011",
30081 => "0101011101110111",
30082 => "0101011101111010",
30083 => "0101011101111110",
30084 => "0101011110000001",
30085 => "0101011110000101",
30086 => "0101011110001001",
30087 => "0101011110001100",
30088 => "0101011110010000",
30089 => "0101011110010100",
30090 => "0101011110010111",
30091 => "0101011110011011",
30092 => "0101011110011110",
30093 => "0101011110100010",
30094 => "0101011110100110",
30095 => "0101011110101001",
30096 => "0101011110101101",
30097 => "0101011110110000",
30098 => "0101011110110100",
30099 => "0101011110111000",
30100 => "0101011110111011",
30101 => "0101011110111111",
30102 => "0101011111000010",
30103 => "0101011111000110",
30104 => "0101011111001010",
30105 => "0101011111001101",
30106 => "0101011111010001",
30107 => "0101011111010100",
30108 => "0101011111011000",
30109 => "0101011111011100",
30110 => "0101011111011111",
30111 => "0101011111100011",
30112 => "0101011111100110",
30113 => "0101011111101010",
30114 => "0101011111101110",
30115 => "0101011111110001",
30116 => "0101011111110101",
30117 => "0101011111111000",
30118 => "0101011111111100",
30119 => "0101100000000000",
30120 => "0101100000000011",
30121 => "0101100000000111",
30122 => "0101100000001010",
30123 => "0101100000001110",
30124 => "0101100000010010",
30125 => "0101100000010101",
30126 => "0101100000011001",
30127 => "0101100000011101",
30128 => "0101100000100000",
30129 => "0101100000100100",
30130 => "0101100000100111",
30131 => "0101100000101011",
30132 => "0101100000101111",
30133 => "0101100000110010",
30134 => "0101100000110110",
30135 => "0101100000111001",
30136 => "0101100000111101",
30137 => "0101100001000001",
30138 => "0101100001000100",
30139 => "0101100001001000",
30140 => "0101100001001100",
30141 => "0101100001001111",
30142 => "0101100001010011",
30143 => "0101100001010110",
30144 => "0101100001011010",
30145 => "0101100001011110",
30146 => "0101100001100001",
30147 => "0101100001100101",
30148 => "0101100001101000",
30149 => "0101100001101100",
30150 => "0101100001110000",
30151 => "0101100001110011",
30152 => "0101100001110111",
30153 => "0101100001111011",
30154 => "0101100001111110",
30155 => "0101100010000010",
30156 => "0101100010000101",
30157 => "0101100010001001",
30158 => "0101100010001101",
30159 => "0101100010010000",
30160 => "0101100010010100",
30161 => "0101100010010111",
30162 => "0101100010011011",
30163 => "0101100010011111",
30164 => "0101100010100010",
30165 => "0101100010100110",
30166 => "0101100010101010",
30167 => "0101100010101101",
30168 => "0101100010110001",
30169 => "0101100010110100",
30170 => "0101100010111000",
30171 => "0101100010111100",
30172 => "0101100010111111",
30173 => "0101100011000011",
30174 => "0101100011000111",
30175 => "0101100011001010",
30176 => "0101100011001110",
30177 => "0101100011010001",
30178 => "0101100011010101",
30179 => "0101100011011001",
30180 => "0101100011011100",
30181 => "0101100011100000",
30182 => "0101100011100100",
30183 => "0101100011100111",
30184 => "0101100011101011",
30185 => "0101100011101110",
30186 => "0101100011110010",
30187 => "0101100011110110",
30188 => "0101100011111001",
30189 => "0101100011111101",
30190 => "0101100100000001",
30191 => "0101100100000100",
30192 => "0101100100001000",
30193 => "0101100100001100",
30194 => "0101100100001111",
30195 => "0101100100010011",
30196 => "0101100100010110",
30197 => "0101100100011010",
30198 => "0101100100011110",
30199 => "0101100100100001",
30200 => "0101100100100101",
30201 => "0101100100101001",
30202 => "0101100100101100",
30203 => "0101100100110000",
30204 => "0101100100110011",
30205 => "0101100100110111",
30206 => "0101100100111011",
30207 => "0101100100111110",
30208 => "0101100101000010",
30209 => "0101100101000110",
30210 => "0101100101001001",
30211 => "0101100101001101",
30212 => "0101100101010001",
30213 => "0101100101010100",
30214 => "0101100101011000",
30215 => "0101100101011011",
30216 => "0101100101011111",
30217 => "0101100101100011",
30218 => "0101100101100110",
30219 => "0101100101101010",
30220 => "0101100101101110",
30221 => "0101100101110001",
30222 => "0101100101110101",
30223 => "0101100101111001",
30224 => "0101100101111100",
30225 => "0101100110000000",
30226 => "0101100110000011",
30227 => "0101100110000111",
30228 => "0101100110001011",
30229 => "0101100110001110",
30230 => "0101100110010010",
30231 => "0101100110010110",
30232 => "0101100110011001",
30233 => "0101100110011101",
30234 => "0101100110100001",
30235 => "0101100110100100",
30236 => "0101100110101000",
30237 => "0101100110101011",
30238 => "0101100110101111",
30239 => "0101100110110011",
30240 => "0101100110110110",
30241 => "0101100110111010",
30242 => "0101100110111110",
30243 => "0101100111000001",
30244 => "0101100111000101",
30245 => "0101100111001001",
30246 => "0101100111001100",
30247 => "0101100111010000",
30248 => "0101100111010100",
30249 => "0101100111010111",
30250 => "0101100111011011",
30251 => "0101100111011110",
30252 => "0101100111100010",
30253 => "0101100111100110",
30254 => "0101100111101001",
30255 => "0101100111101101",
30256 => "0101100111110001",
30257 => "0101100111110100",
30258 => "0101100111111000",
30259 => "0101100111111100",
30260 => "0101100111111111",
30261 => "0101101000000011",
30262 => "0101101000000111",
30263 => "0101101000001010",
30264 => "0101101000001110",
30265 => "0101101000010010",
30266 => "0101101000010101",
30267 => "0101101000011001",
30268 => "0101101000011100",
30269 => "0101101000100000",
30270 => "0101101000100100",
30271 => "0101101000100111",
30272 => "0101101000101011",
30273 => "0101101000101111",
30274 => "0101101000110010",
30275 => "0101101000110110",
30276 => "0101101000111010",
30277 => "0101101000111101",
30278 => "0101101001000001",
30279 => "0101101001000101",
30280 => "0101101001001000",
30281 => "0101101001001100",
30282 => "0101101001010000",
30283 => "0101101001010011",
30284 => "0101101001010111",
30285 => "0101101001011011",
30286 => "0101101001011110",
30287 => "0101101001100010",
30288 => "0101101001100110",
30289 => "0101101001101001",
30290 => "0101101001101101",
30291 => "0101101001110000",
30292 => "0101101001110100",
30293 => "0101101001111000",
30294 => "0101101001111011",
30295 => "0101101001111111",
30296 => "0101101010000011",
30297 => "0101101010000110",
30298 => "0101101010001010",
30299 => "0101101010001110",
30300 => "0101101010010001",
30301 => "0101101010010101",
30302 => "0101101010011001",
30303 => "0101101010011100",
30304 => "0101101010100000",
30305 => "0101101010100100",
30306 => "0101101010100111",
30307 => "0101101010101011",
30308 => "0101101010101111",
30309 => "0101101010110010",
30310 => "0101101010110110",
30311 => "0101101010111010",
30312 => "0101101010111101",
30313 => "0101101011000001",
30314 => "0101101011000101",
30315 => "0101101011001000",
30316 => "0101101011001100",
30317 => "0101101011010000",
30318 => "0101101011010011",
30319 => "0101101011010111",
30320 => "0101101011011011",
30321 => "0101101011011110",
30322 => "0101101011100010",
30323 => "0101101011100110",
30324 => "0101101011101001",
30325 => "0101101011101101",
30326 => "0101101011110001",
30327 => "0101101011110100",
30328 => "0101101011111000",
30329 => "0101101011111100",
30330 => "0101101011111111",
30331 => "0101101100000011",
30332 => "0101101100000111",
30333 => "0101101100001010",
30334 => "0101101100001110",
30335 => "0101101100010010",
30336 => "0101101100010101",
30337 => "0101101100011001",
30338 => "0101101100011101",
30339 => "0101101100100000",
30340 => "0101101100100100",
30341 => "0101101100101000",
30342 => "0101101100101011",
30343 => "0101101100101111",
30344 => "0101101100110011",
30345 => "0101101100110110",
30346 => "0101101100111010",
30347 => "0101101100111110",
30348 => "0101101101000001",
30349 => "0101101101000101",
30350 => "0101101101001001",
30351 => "0101101101001100",
30352 => "0101101101010000",
30353 => "0101101101010100",
30354 => "0101101101010111",
30355 => "0101101101011011",
30356 => "0101101101011111",
30357 => "0101101101100010",
30358 => "0101101101100110",
30359 => "0101101101101010",
30360 => "0101101101101101",
30361 => "0101101101110001",
30362 => "0101101101110101",
30363 => "0101101101111000",
30364 => "0101101101111100",
30365 => "0101101110000000",
30366 => "0101101110000011",
30367 => "0101101110000111",
30368 => "0101101110001011",
30369 => "0101101110001110",
30370 => "0101101110010010",
30371 => "0101101110010110",
30372 => "0101101110011001",
30373 => "0101101110011101",
30374 => "0101101110100001",
30375 => "0101101110100100",
30376 => "0101101110101000",
30377 => "0101101110101100",
30378 => "0101101110110000",
30379 => "0101101110110011",
30380 => "0101101110110111",
30381 => "0101101110111011",
30382 => "0101101110111110",
30383 => "0101101111000010",
30384 => "0101101111000110",
30385 => "0101101111001001",
30386 => "0101101111001101",
30387 => "0101101111010001",
30388 => "0101101111010100",
30389 => "0101101111011000",
30390 => "0101101111011100",
30391 => "0101101111011111",
30392 => "0101101111100011",
30393 => "0101101111100111",
30394 => "0101101111101010",
30395 => "0101101111101110",
30396 => "0101101111110010",
30397 => "0101101111110101",
30398 => "0101101111111001",
30399 => "0101101111111101",
30400 => "0101110000000000",
30401 => "0101110000000100",
30402 => "0101110000001000",
30403 => "0101110000001100",
30404 => "0101110000001111",
30405 => "0101110000010011",
30406 => "0101110000010111",
30407 => "0101110000011010",
30408 => "0101110000011110",
30409 => "0101110000100010",
30410 => "0101110000100101",
30411 => "0101110000101001",
30412 => "0101110000101101",
30413 => "0101110000110000",
30414 => "0101110000110100",
30415 => "0101110000111000",
30416 => "0101110000111011",
30417 => "0101110000111111",
30418 => "0101110001000011",
30419 => "0101110001000111",
30420 => "0101110001001010",
30421 => "0101110001001110",
30422 => "0101110001010010",
30423 => "0101110001010101",
30424 => "0101110001011001",
30425 => "0101110001011101",
30426 => "0101110001100000",
30427 => "0101110001100100",
30428 => "0101110001101000",
30429 => "0101110001101011",
30430 => "0101110001101111",
30431 => "0101110001110011",
30432 => "0101110001110111",
30433 => "0101110001111010",
30434 => "0101110001111110",
30435 => "0101110010000010",
30436 => "0101110010000101",
30437 => "0101110010001001",
30438 => "0101110010001101",
30439 => "0101110010010000",
30440 => "0101110010010100",
30441 => "0101110010011000",
30442 => "0101110010011011",
30443 => "0101110010011111",
30444 => "0101110010100011",
30445 => "0101110010100111",
30446 => "0101110010101010",
30447 => "0101110010101110",
30448 => "0101110010110010",
30449 => "0101110010110101",
30450 => "0101110010111001",
30451 => "0101110010111101",
30452 => "0101110011000000",
30453 => "0101110011000100",
30454 => "0101110011001000",
30455 => "0101110011001011",
30456 => "0101110011001111",
30457 => "0101110011010011",
30458 => "0101110011010111",
30459 => "0101110011011010",
30460 => "0101110011011110",
30461 => "0101110011100010",
30462 => "0101110011100101",
30463 => "0101110011101001",
30464 => "0101110011101101",
30465 => "0101110011110000",
30466 => "0101110011110100",
30467 => "0101110011111000",
30468 => "0101110011111100",
30469 => "0101110011111111",
30470 => "0101110100000011",
30471 => "0101110100000111",
30472 => "0101110100001010",
30473 => "0101110100001110",
30474 => "0101110100010010",
30475 => "0101110100010101",
30476 => "0101110100011001",
30477 => "0101110100011101",
30478 => "0101110100100001",
30479 => "0101110100100100",
30480 => "0101110100101000",
30481 => "0101110100101100",
30482 => "0101110100101111",
30483 => "0101110100110011",
30484 => "0101110100110111",
30485 => "0101110100111011",
30486 => "0101110100111110",
30487 => "0101110101000010",
30488 => "0101110101000110",
30489 => "0101110101001001",
30490 => "0101110101001101",
30491 => "0101110101010001",
30492 => "0101110101010100",
30493 => "0101110101011000",
30494 => "0101110101011100",
30495 => "0101110101100000",
30496 => "0101110101100011",
30497 => "0101110101100111",
30498 => "0101110101101011",
30499 => "0101110101101110",
30500 => "0101110101110010",
30501 => "0101110101110110",
30502 => "0101110101111010",
30503 => "0101110101111101",
30504 => "0101110110000001",
30505 => "0101110110000101",
30506 => "0101110110001000",
30507 => "0101110110001100",
30508 => "0101110110010000",
30509 => "0101110110010100",
30510 => "0101110110010111",
30511 => "0101110110011011",
30512 => "0101110110011111",
30513 => "0101110110100010",
30514 => "0101110110100110",
30515 => "0101110110101010",
30516 => "0101110110101101",
30517 => "0101110110110001",
30518 => "0101110110110101",
30519 => "0101110110111001",
30520 => "0101110110111100",
30521 => "0101110111000000",
30522 => "0101110111000100",
30523 => "0101110111000111",
30524 => "0101110111001011",
30525 => "0101110111001111",
30526 => "0101110111010011",
30527 => "0101110111010110",
30528 => "0101110111011010",
30529 => "0101110111011110",
30530 => "0101110111100001",
30531 => "0101110111100101",
30532 => "0101110111101001",
30533 => "0101110111101101",
30534 => "0101110111110000",
30535 => "0101110111110100",
30536 => "0101110111111000",
30537 => "0101110111111100",
30538 => "0101110111111111",
30539 => "0101111000000011",
30540 => "0101111000000111",
30541 => "0101111000001010",
30542 => "0101111000001110",
30543 => "0101111000010010",
30544 => "0101111000010110",
30545 => "0101111000011001",
30546 => "0101111000011101",
30547 => "0101111000100001",
30548 => "0101111000100100",
30549 => "0101111000101000",
30550 => "0101111000101100",
30551 => "0101111000110000",
30552 => "0101111000110011",
30553 => "0101111000110111",
30554 => "0101111000111011",
30555 => "0101111000111110",
30556 => "0101111001000010",
30557 => "0101111001000110",
30558 => "0101111001001010",
30559 => "0101111001001101",
30560 => "0101111001010001",
30561 => "0101111001010101",
30562 => "0101111001011001",
30563 => "0101111001011100",
30564 => "0101111001100000",
30565 => "0101111001100100",
30566 => "0101111001100111",
30567 => "0101111001101011",
30568 => "0101111001101111",
30569 => "0101111001110011",
30570 => "0101111001110110",
30571 => "0101111001111010",
30572 => "0101111001111110",
30573 => "0101111010000001",
30574 => "0101111010000101",
30575 => "0101111010001001",
30576 => "0101111010001101",
30577 => "0101111010010000",
30578 => "0101111010010100",
30579 => "0101111010011000",
30580 => "0101111010011100",
30581 => "0101111010011111",
30582 => "0101111010100011",
30583 => "0101111010100111",
30584 => "0101111010101010",
30585 => "0101111010101110",
30586 => "0101111010110010",
30587 => "0101111010110110",
30588 => "0101111010111001",
30589 => "0101111010111101",
30590 => "0101111011000001",
30591 => "0101111011000101",
30592 => "0101111011001000",
30593 => "0101111011001100",
30594 => "0101111011010000",
30595 => "0101111011010100",
30596 => "0101111011010111",
30597 => "0101111011011011",
30598 => "0101111011011111",
30599 => "0101111011100010",
30600 => "0101111011100110",
30601 => "0101111011101010",
30602 => "0101111011101110",
30603 => "0101111011110001",
30604 => "0101111011110101",
30605 => "0101111011111001",
30606 => "0101111011111101",
30607 => "0101111100000000",
30608 => "0101111100000100",
30609 => "0101111100001000",
30610 => "0101111100001100",
30611 => "0101111100001111",
30612 => "0101111100010011",
30613 => "0101111100010111",
30614 => "0101111100011010",
30615 => "0101111100011110",
30616 => "0101111100100010",
30617 => "0101111100100110",
30618 => "0101111100101001",
30619 => "0101111100101101",
30620 => "0101111100110001",
30621 => "0101111100110101",
30622 => "0101111100111000",
30623 => "0101111100111100",
30624 => "0101111101000000",
30625 => "0101111101000100",
30626 => "0101111101000111",
30627 => "0101111101001011",
30628 => "0101111101001111",
30629 => "0101111101010011",
30630 => "0101111101010110",
30631 => "0101111101011010",
30632 => "0101111101011110",
30633 => "0101111101100001",
30634 => "0101111101100101",
30635 => "0101111101101001",
30636 => "0101111101101101",
30637 => "0101111101110000",
30638 => "0101111101110100",
30639 => "0101111101111000",
30640 => "0101111101111100",
30641 => "0101111101111111",
30642 => "0101111110000011",
30643 => "0101111110000111",
30644 => "0101111110001011",
30645 => "0101111110001110",
30646 => "0101111110010010",
30647 => "0101111110010110",
30648 => "0101111110011010",
30649 => "0101111110011101",
30650 => "0101111110100001",
30651 => "0101111110100101",
30652 => "0101111110101001",
30653 => "0101111110101100",
30654 => "0101111110110000",
30655 => "0101111110110100",
30656 => "0101111110111000",
30657 => "0101111110111011",
30658 => "0101111110111111",
30659 => "0101111111000011",
30660 => "0101111111000111",
30661 => "0101111111001010",
30662 => "0101111111001110",
30663 => "0101111111010010",
30664 => "0101111111010110",
30665 => "0101111111011001",
30666 => "0101111111011101",
30667 => "0101111111100001",
30668 => "0101111111100101",
30669 => "0101111111101000",
30670 => "0101111111101100",
30671 => "0101111111110000",
30672 => "0101111111110100",
30673 => "0101111111110111",
30674 => "0101111111111011",
30675 => "0101111111111111",
30676 => "0110000000000011",
30677 => "0110000000000110",
30678 => "0110000000001010",
30679 => "0110000000001110",
30680 => "0110000000010010",
30681 => "0110000000010101",
30682 => "0110000000011001",
30683 => "0110000000011101",
30684 => "0110000000100001",
30685 => "0110000000100100",
30686 => "0110000000101000",
30687 => "0110000000101100",
30688 => "0110000000110000",
30689 => "0110000000110011",
30690 => "0110000000110111",
30691 => "0110000000111011",
30692 => "0110000000111111",
30693 => "0110000001000010",
30694 => "0110000001000110",
30695 => "0110000001001010",
30696 => "0110000001001110",
30697 => "0110000001010001",
30698 => "0110000001010101",
30699 => "0110000001011001",
30700 => "0110000001011101",
30701 => "0110000001100000",
30702 => "0110000001100100",
30703 => "0110000001101000",
30704 => "0110000001101100",
30705 => "0110000001101111",
30706 => "0110000001110011",
30707 => "0110000001110111",
30708 => "0110000001111011",
30709 => "0110000001111110",
30710 => "0110000010000010",
30711 => "0110000010000110",
30712 => "0110000010001010",
30713 => "0110000010001101",
30714 => "0110000010010001",
30715 => "0110000010010101",
30716 => "0110000010011001",
30717 => "0110000010011100",
30718 => "0110000010100000",
30719 => "0110000010100100",
30720 => "0110000010101000",
30721 => "0110000010101100",
30722 => "0110000010101111",
30723 => "0110000010110011",
30724 => "0110000010110111",
30725 => "0110000010111011",
30726 => "0110000010111110",
30727 => "0110000011000010",
30728 => "0110000011000110",
30729 => "0110000011001010",
30730 => "0110000011001101",
30731 => "0110000011010001",
30732 => "0110000011010101",
30733 => "0110000011011001",
30734 => "0110000011011100",
30735 => "0110000011100000",
30736 => "0110000011100100",
30737 => "0110000011101000",
30738 => "0110000011101011",
30739 => "0110000011101111",
30740 => "0110000011110011",
30741 => "0110000011110111",
30742 => "0110000011111011",
30743 => "0110000011111110",
30744 => "0110000100000010",
30745 => "0110000100000110",
30746 => "0110000100001010",
30747 => "0110000100001101",
30748 => "0110000100010001",
30749 => "0110000100010101",
30750 => "0110000100011001",
30751 => "0110000100011100",
30752 => "0110000100100000",
30753 => "0110000100100100",
30754 => "0110000100101000",
30755 => "0110000100101100",
30756 => "0110000100101111",
30757 => "0110000100110011",
30758 => "0110000100110111",
30759 => "0110000100111011",
30760 => "0110000100111110",
30761 => "0110000101000010",
30762 => "0110000101000110",
30763 => "0110000101001010",
30764 => "0110000101001101",
30765 => "0110000101010001",
30766 => "0110000101010101",
30767 => "0110000101011001",
30768 => "0110000101011101",
30769 => "0110000101100000",
30770 => "0110000101100100",
30771 => "0110000101101000",
30772 => "0110000101101100",
30773 => "0110000101101111",
30774 => "0110000101110011",
30775 => "0110000101110111",
30776 => "0110000101111011",
30777 => "0110000101111110",
30778 => "0110000110000010",
30779 => "0110000110000110",
30780 => "0110000110001010",
30781 => "0110000110001110",
30782 => "0110000110010001",
30783 => "0110000110010101",
30784 => "0110000110011001",
30785 => "0110000110011101",
30786 => "0110000110100000",
30787 => "0110000110100100",
30788 => "0110000110101000",
30789 => "0110000110101100",
30790 => "0110000110110000",
30791 => "0110000110110011",
30792 => "0110000110110111",
30793 => "0110000110111011",
30794 => "0110000110111111",
30795 => "0110000111000010",
30796 => "0110000111000110",
30797 => "0110000111001010",
30798 => "0110000111001110",
30799 => "0110000111010010",
30800 => "0110000111010101",
30801 => "0110000111011001",
30802 => "0110000111011101",
30803 => "0110000111100001",
30804 => "0110000111100100",
30805 => "0110000111101000",
30806 => "0110000111101100",
30807 => "0110000111110000",
30808 => "0110000111110100",
30809 => "0110000111110111",
30810 => "0110000111111011",
30811 => "0110000111111111",
30812 => "0110001000000011",
30813 => "0110001000000110",
30814 => "0110001000001010",
30815 => "0110001000001110",
30816 => "0110001000010010",
30817 => "0110001000010110",
30818 => "0110001000011001",
30819 => "0110001000011101",
30820 => "0110001000100001",
30821 => "0110001000100101",
30822 => "0110001000101000",
30823 => "0110001000101100",
30824 => "0110001000110000",
30825 => "0110001000110100",
30826 => "0110001000111000",
30827 => "0110001000111011",
30828 => "0110001000111111",
30829 => "0110001001000011",
30830 => "0110001001000111",
30831 => "0110001001001011",
30832 => "0110001001001110",
30833 => "0110001001010010",
30834 => "0110001001010110",
30835 => "0110001001011010",
30836 => "0110001001011101",
30837 => "0110001001100001",
30838 => "0110001001100101",
30839 => "0110001001101001",
30840 => "0110001001101101",
30841 => "0110001001110000",
30842 => "0110001001110100",
30843 => "0110001001111000",
30844 => "0110001001111100",
30845 => "0110001010000000",
30846 => "0110001010000011",
30847 => "0110001010000111",
30848 => "0110001010001011",
30849 => "0110001010001111",
30850 => "0110001010010010",
30851 => "0110001010010110",
30852 => "0110001010011010",
30853 => "0110001010011110",
30854 => "0110001010100010",
30855 => "0110001010100101",
30856 => "0110001010101001",
30857 => "0110001010101101",
30858 => "0110001010110001",
30859 => "0110001010110101",
30860 => "0110001010111000",
30861 => "0110001010111100",
30862 => "0110001011000000",
30863 => "0110001011000100",
30864 => "0110001011001000",
30865 => "0110001011001011",
30866 => "0110001011001111",
30867 => "0110001011010011",
30868 => "0110001011010111",
30869 => "0110001011011010",
30870 => "0110001011011110",
30871 => "0110001011100010",
30872 => "0110001011100110",
30873 => "0110001011101010",
30874 => "0110001011101101",
30875 => "0110001011110001",
30876 => "0110001011110101",
30877 => "0110001011111001",
30878 => "0110001011111101",
30879 => "0110001100000000",
30880 => "0110001100000100",
30881 => "0110001100001000",
30882 => "0110001100001100",
30883 => "0110001100010000",
30884 => "0110001100010011",
30885 => "0110001100010111",
30886 => "0110001100011011",
30887 => "0110001100011111",
30888 => "0110001100100011",
30889 => "0110001100100110",
30890 => "0110001100101010",
30891 => "0110001100101110",
30892 => "0110001100110010",
30893 => "0110001100110110",
30894 => "0110001100111001",
30895 => "0110001100111101",
30896 => "0110001101000001",
30897 => "0110001101000101",
30898 => "0110001101001001",
30899 => "0110001101001100",
30900 => "0110001101010000",
30901 => "0110001101010100",
30902 => "0110001101011000",
30903 => "0110001101011100",
30904 => "0110001101011111",
30905 => "0110001101100011",
30906 => "0110001101100111",
30907 => "0110001101101011",
30908 => "0110001101101111",
30909 => "0110001101110010",
30910 => "0110001101110110",
30911 => "0110001101111010",
30912 => "0110001101111110",
30913 => "0110001110000010",
30914 => "0110001110000101",
30915 => "0110001110001001",
30916 => "0110001110001101",
30917 => "0110001110010001",
30918 => "0110001110010101",
30919 => "0110001110011000",
30920 => "0110001110011100",
30921 => "0110001110100000",
30922 => "0110001110100100",
30923 => "0110001110101000",
30924 => "0110001110101011",
30925 => "0110001110101111",
30926 => "0110001110110011",
30927 => "0110001110110111",
30928 => "0110001110111011",
30929 => "0110001110111110",
30930 => "0110001111000010",
30931 => "0110001111000110",
30932 => "0110001111001010",
30933 => "0110001111001110",
30934 => "0110001111010001",
30935 => "0110001111010101",
30936 => "0110001111011001",
30937 => "0110001111011101",
30938 => "0110001111100001",
30939 => "0110001111100100",
30940 => "0110001111101000",
30941 => "0110001111101100",
30942 => "0110001111110000",
30943 => "0110001111110100",
30944 => "0110001111111000",
30945 => "0110001111111011",
30946 => "0110001111111111",
30947 => "0110010000000011",
30948 => "0110010000000111",
30949 => "0110010000001011",
30950 => "0110010000001110",
30951 => "0110010000010010",
30952 => "0110010000010110",
30953 => "0110010000011010",
30954 => "0110010000011110",
30955 => "0110010000100001",
30956 => "0110010000100101",
30957 => "0110010000101001",
30958 => "0110010000101101",
30959 => "0110010000110001",
30960 => "0110010000110100",
30961 => "0110010000111000",
30962 => "0110010000111100",
30963 => "0110010001000000",
30964 => "0110010001000100",
30965 => "0110010001001000",
30966 => "0110010001001011",
30967 => "0110010001001111",
30968 => "0110010001010011",
30969 => "0110010001010111",
30970 => "0110010001011011",
30971 => "0110010001011110",
30972 => "0110010001100010",
30973 => "0110010001100110",
30974 => "0110010001101010",
30975 => "0110010001101110",
30976 => "0110010001110001",
30977 => "0110010001110101",
30978 => "0110010001111001",
30979 => "0110010001111101",
30980 => "0110010010000001",
30981 => "0110010010000101",
30982 => "0110010010001000",
30983 => "0110010010001100",
30984 => "0110010010010000",
30985 => "0110010010010100",
30986 => "0110010010011000",
30987 => "0110010010011011",
30988 => "0110010010011111",
30989 => "0110010010100011",
30990 => "0110010010100111",
30991 => "0110010010101011",
30992 => "0110010010101111",
30993 => "0110010010110010",
30994 => "0110010010110110",
30995 => "0110010010111010",
30996 => "0110010010111110",
30997 => "0110010011000010",
30998 => "0110010011000101",
30999 => "0110010011001001",
31000 => "0110010011001101",
31001 => "0110010011010001",
31002 => "0110010011010101",
31003 => "0110010011011001",
31004 => "0110010011011100",
31005 => "0110010011100000",
31006 => "0110010011100100",
31007 => "0110010011101000",
31008 => "0110010011101100",
31009 => "0110010011101111",
31010 => "0110010011110011",
31011 => "0110010011110111",
31012 => "0110010011111011",
31013 => "0110010011111111",
31014 => "0110010100000011",
31015 => "0110010100000110",
31016 => "0110010100001010",
31017 => "0110010100001110",
31018 => "0110010100010010",
31019 => "0110010100010110",
31020 => "0110010100011010",
31021 => "0110010100011101",
31022 => "0110010100100001",
31023 => "0110010100100101",
31024 => "0110010100101001",
31025 => "0110010100101101",
31026 => "0110010100110000",
31027 => "0110010100110100",
31028 => "0110010100111000",
31029 => "0110010100111100",
31030 => "0110010101000000",
31031 => "0110010101000100",
31032 => "0110010101000111",
31033 => "0110010101001011",
31034 => "0110010101001111",
31035 => "0110010101010011",
31036 => "0110010101010111",
31037 => "0110010101011011",
31038 => "0110010101011110",
31039 => "0110010101100010",
31040 => "0110010101100110",
31041 => "0110010101101010",
31042 => "0110010101101110",
31043 => "0110010101110010",
31044 => "0110010101110101",
31045 => "0110010101111001",
31046 => "0110010101111101",
31047 => "0110010110000001",
31048 => "0110010110000101",
31049 => "0110010110001000",
31050 => "0110010110001100",
31051 => "0110010110010000",
31052 => "0110010110010100",
31053 => "0110010110011000",
31054 => "0110010110011100",
31055 => "0110010110011111",
31056 => "0110010110100011",
31057 => "0110010110100111",
31058 => "0110010110101011",
31059 => "0110010110101111",
31060 => "0110010110110011",
31061 => "0110010110110110",
31062 => "0110010110111010",
31063 => "0110010110111110",
31064 => "0110010111000010",
31065 => "0110010111000110",
31066 => "0110010111001010",
31067 => "0110010111001101",
31068 => "0110010111010001",
31069 => "0110010111010101",
31070 => "0110010111011001",
31071 => "0110010111011101",
31072 => "0110010111100001",
31073 => "0110010111100100",
31074 => "0110010111101000",
31075 => "0110010111101100",
31076 => "0110010111110000",
31077 => "0110010111110100",
31078 => "0110010111111000",
31079 => "0110010111111011",
31080 => "0110010111111111",
31081 => "0110011000000011",
31082 => "0110011000000111",
31083 => "0110011000001011",
31084 => "0110011000001111",
31085 => "0110011000010010",
31086 => "0110011000010110",
31087 => "0110011000011010",
31088 => "0110011000011110",
31089 => "0110011000100010",
31090 => "0110011000100110",
31091 => "0110011000101001",
31092 => "0110011000101101",
31093 => "0110011000110001",
31094 => "0110011000110101",
31095 => "0110011000111001",
31096 => "0110011000111101",
31097 => "0110011001000001",
31098 => "0110011001000100",
31099 => "0110011001001000",
31100 => "0110011001001100",
31101 => "0110011001010000",
31102 => "0110011001010100",
31103 => "0110011001011000",
31104 => "0110011001011011",
31105 => "0110011001011111",
31106 => "0110011001100011",
31107 => "0110011001100111",
31108 => "0110011001101011",
31109 => "0110011001101111",
31110 => "0110011001110010",
31111 => "0110011001110110",
31112 => "0110011001111010",
31113 => "0110011001111110",
31114 => "0110011010000010",
31115 => "0110011010000110",
31116 => "0110011010001001",
31117 => "0110011010001101",
31118 => "0110011010010001",
31119 => "0110011010010101",
31120 => "0110011010011001",
31121 => "0110011010011101",
31122 => "0110011010100001",
31123 => "0110011010100100",
31124 => "0110011010101000",
31125 => "0110011010101100",
31126 => "0110011010110000",
31127 => "0110011010110100",
31128 => "0110011010111000",
31129 => "0110011010111011",
31130 => "0110011010111111",
31131 => "0110011011000011",
31132 => "0110011011000111",
31133 => "0110011011001011",
31134 => "0110011011001111",
31135 => "0110011011010010",
31136 => "0110011011010110",
31137 => "0110011011011010",
31138 => "0110011011011110",
31139 => "0110011011100010",
31140 => "0110011011100110",
31141 => "0110011011101010",
31142 => "0110011011101101",
31143 => "0110011011110001",
31144 => "0110011011110101",
31145 => "0110011011111001",
31146 => "0110011011111101",
31147 => "0110011100000001",
31148 => "0110011100000100",
31149 => "0110011100001000",
31150 => "0110011100001100",
31151 => "0110011100010000",
31152 => "0110011100010100",
31153 => "0110011100011000",
31154 => "0110011100011100",
31155 => "0110011100011111",
31156 => "0110011100100011",
31157 => "0110011100100111",
31158 => "0110011100101011",
31159 => "0110011100101111",
31160 => "0110011100110011",
31161 => "0110011100110111",
31162 => "0110011100111010",
31163 => "0110011100111110",
31164 => "0110011101000010",
31165 => "0110011101000110",
31166 => "0110011101001010",
31167 => "0110011101001110",
31168 => "0110011101010001",
31169 => "0110011101010101",
31170 => "0110011101011001",
31171 => "0110011101011101",
31172 => "0110011101100001",
31173 => "0110011101100101",
31174 => "0110011101101001",
31175 => "0110011101101100",
31176 => "0110011101110000",
31177 => "0110011101110100",
31178 => "0110011101111000",
31179 => "0110011101111100",
31180 => "0110011110000000",
31181 => "0110011110000100",
31182 => "0110011110000111",
31183 => "0110011110001011",
31184 => "0110011110001111",
31185 => "0110011110010011",
31186 => "0110011110010111",
31187 => "0110011110011011",
31188 => "0110011110011111",
31189 => "0110011110100010",
31190 => "0110011110100110",
31191 => "0110011110101010",
31192 => "0110011110101110",
31193 => "0110011110110010",
31194 => "0110011110110110",
31195 => "0110011110111010",
31196 => "0110011110111101",
31197 => "0110011111000001",
31198 => "0110011111000101",
31199 => "0110011111001001",
31200 => "0110011111001101",
31201 => "0110011111010001",
31202 => "0110011111010101",
31203 => "0110011111011000",
31204 => "0110011111011100",
31205 => "0110011111100000",
31206 => "0110011111100100",
31207 => "0110011111101000",
31208 => "0110011111101100",
31209 => "0110011111110000",
31210 => "0110011111110011",
31211 => "0110011111110111",
31212 => "0110011111111011",
31213 => "0110011111111111",
31214 => "0110100000000011",
31215 => "0110100000000111",
31216 => "0110100000001011",
31217 => "0110100000001110",
31218 => "0110100000010010",
31219 => "0110100000010110",
31220 => "0110100000011010",
31221 => "0110100000011110",
31222 => "0110100000100010",
31223 => "0110100000100110",
31224 => "0110100000101001",
31225 => "0110100000101101",
31226 => "0110100000110001",
31227 => "0110100000110101",
31228 => "0110100000111001",
31229 => "0110100000111101",
31230 => "0110100001000001",
31231 => "0110100001000100",
31232 => "0110100001001000",
31233 => "0110100001001100",
31234 => "0110100001010000",
31235 => "0110100001010100",
31236 => "0110100001011000",
31237 => "0110100001011100",
31238 => "0110100001100000",
31239 => "0110100001100011",
31240 => "0110100001100111",
31241 => "0110100001101011",
31242 => "0110100001101111",
31243 => "0110100001110011",
31244 => "0110100001110111",
31245 => "0110100001111011",
31246 => "0110100001111110",
31247 => "0110100010000010",
31248 => "0110100010000110",
31249 => "0110100010001010",
31250 => "0110100010001110",
31251 => "0110100010010010",
31252 => "0110100010010110",
31253 => "0110100010011001",
31254 => "0110100010011101",
31255 => "0110100010100001",
31256 => "0110100010100101",
31257 => "0110100010101001",
31258 => "0110100010101101",
31259 => "0110100010110001",
31260 => "0110100010110101",
31261 => "0110100010111000",
31262 => "0110100010111100",
31263 => "0110100011000000",
31264 => "0110100011000100",
31265 => "0110100011001000",
31266 => "0110100011001100",
31267 => "0110100011010000",
31268 => "0110100011010100",
31269 => "0110100011010111",
31270 => "0110100011011011",
31271 => "0110100011011111",
31272 => "0110100011100011",
31273 => "0110100011100111",
31274 => "0110100011101011",
31275 => "0110100011101111",
31276 => "0110100011110010",
31277 => "0110100011110110",
31278 => "0110100011111010",
31279 => "0110100011111110",
31280 => "0110100100000010",
31281 => "0110100100000110",
31282 => "0110100100001010",
31283 => "0110100100001110",
31284 => "0110100100010001",
31285 => "0110100100010101",
31286 => "0110100100011001",
31287 => "0110100100011101",
31288 => "0110100100100001",
31289 => "0110100100100101",
31290 => "0110100100101001",
31291 => "0110100100101101",
31292 => "0110100100110000",
31293 => "0110100100110100",
31294 => "0110100100111000",
31295 => "0110100100111100",
31296 => "0110100101000000",
31297 => "0110100101000100",
31298 => "0110100101001000",
31299 => "0110100101001100",
31300 => "0110100101001111",
31301 => "0110100101010011",
31302 => "0110100101010111",
31303 => "0110100101011011",
31304 => "0110100101011111",
31305 => "0110100101100011",
31306 => "0110100101100111",
31307 => "0110100101101011",
31308 => "0110100101101110",
31309 => "0110100101110010",
31310 => "0110100101110110",
31311 => "0110100101111010",
31312 => "0110100101111110",
31313 => "0110100110000010",
31314 => "0110100110000110",
31315 => "0110100110001010",
31316 => "0110100110001101",
31317 => "0110100110010001",
31318 => "0110100110010101",
31319 => "0110100110011001",
31320 => "0110100110011101",
31321 => "0110100110100001",
31322 => "0110100110100101",
31323 => "0110100110101001",
31324 => "0110100110101100",
31325 => "0110100110110000",
31326 => "0110100110110100",
31327 => "0110100110111000",
31328 => "0110100110111100",
31329 => "0110100111000000",
31330 => "0110100111000100",
31331 => "0110100111001000",
31332 => "0110100111001011",
31333 => "0110100111001111",
31334 => "0110100111010011",
31335 => "0110100111010111",
31336 => "0110100111011011",
31337 => "0110100111011111",
31338 => "0110100111100011",
31339 => "0110100111100111",
31340 => "0110100111101011",
31341 => "0110100111101110",
31342 => "0110100111110010",
31343 => "0110100111110110",
31344 => "0110100111111010",
31345 => "0110100111111110",
31346 => "0110101000000010",
31347 => "0110101000000110",
31348 => "0110101000001010",
31349 => "0110101000001101",
31350 => "0110101000010001",
31351 => "0110101000010101",
31352 => "0110101000011001",
31353 => "0110101000011101",
31354 => "0110101000100001",
31355 => "0110101000100101",
31356 => "0110101000101001",
31357 => "0110101000101101",
31358 => "0110101000110000",
31359 => "0110101000110100",
31360 => "0110101000111000",
31361 => "0110101000111100",
31362 => "0110101001000000",
31363 => "0110101001000100",
31364 => "0110101001001000",
31365 => "0110101001001100",
31366 => "0110101001001111",
31367 => "0110101001010011",
31368 => "0110101001010111",
31369 => "0110101001011011",
31370 => "0110101001011111",
31371 => "0110101001100011",
31372 => "0110101001100111",
31373 => "0110101001101011",
31374 => "0110101001101111",
31375 => "0110101001110010",
31376 => "0110101001110110",
31377 => "0110101001111010",
31378 => "0110101001111110",
31379 => "0110101010000010",
31380 => "0110101010000110",
31381 => "0110101010001010",
31382 => "0110101010001110",
31383 => "0110101010010010",
31384 => "0110101010010101",
31385 => "0110101010011001",
31386 => "0110101010011101",
31387 => "0110101010100001",
31388 => "0110101010100101",
31389 => "0110101010101001",
31390 => "0110101010101101",
31391 => "0110101010110001",
31392 => "0110101010110101",
31393 => "0110101010111000",
31394 => "0110101010111100",
31395 => "0110101011000000",
31396 => "0110101011000100",
31397 => "0110101011001000",
31398 => "0110101011001100",
31399 => "0110101011010000",
31400 => "0110101011010100",
31401 => "0110101011011000",
31402 => "0110101011011011",
31403 => "0110101011011111",
31404 => "0110101011100011",
31405 => "0110101011100111",
31406 => "0110101011101011",
31407 => "0110101011101111",
31408 => "0110101011110011",
31409 => "0110101011110111",
31410 => "0110101011111011",
31411 => "0110101011111110",
31412 => "0110101100000010",
31413 => "0110101100000110",
31414 => "0110101100001010",
31415 => "0110101100001110",
31416 => "0110101100010010",
31417 => "0110101100010110",
31418 => "0110101100011010",
31419 => "0110101100011110",
31420 => "0110101100100010",
31421 => "0110101100100101",
31422 => "0110101100101001",
31423 => "0110101100101101",
31424 => "0110101100110001",
31425 => "0110101100110101",
31426 => "0110101100111001",
31427 => "0110101100111101",
31428 => "0110101101000001",
31429 => "0110101101000101",
31430 => "0110101101001000",
31431 => "0110101101001100",
31432 => "0110101101010000",
31433 => "0110101101010100",
31434 => "0110101101011000",
31435 => "0110101101011100",
31436 => "0110101101100000",
31437 => "0110101101100100",
31438 => "0110101101101000",
31439 => "0110101101101100",
31440 => "0110101101101111",
31441 => "0110101101110011",
31442 => "0110101101110111",
31443 => "0110101101111011",
31444 => "0110101101111111",
31445 => "0110101110000011",
31446 => "0110101110000111",
31447 => "0110101110001011",
31448 => "0110101110001111",
31449 => "0110101110010010",
31450 => "0110101110010110",
31451 => "0110101110011010",
31452 => "0110101110011110",
31453 => "0110101110100010",
31454 => "0110101110100110",
31455 => "0110101110101010",
31456 => "0110101110101110",
31457 => "0110101110110010",
31458 => "0110101110110110",
31459 => "0110101110111001",
31460 => "0110101110111101",
31461 => "0110101111000001",
31462 => "0110101111000101",
31463 => "0110101111001001",
31464 => "0110101111001101",
31465 => "0110101111010001",
31466 => "0110101111010101",
31467 => "0110101111011001",
31468 => "0110101111011101",
31469 => "0110101111100000",
31470 => "0110101111100100",
31471 => "0110101111101000",
31472 => "0110101111101100",
31473 => "0110101111110000",
31474 => "0110101111110100",
31475 => "0110101111111000",
31476 => "0110101111111100",
31477 => "0110110000000000",
31478 => "0110110000000100",
31479 => "0110110000001000",
31480 => "0110110000001011",
31481 => "0110110000001111",
31482 => "0110110000010011",
31483 => "0110110000010111",
31484 => "0110110000011011",
31485 => "0110110000011111",
31486 => "0110110000100011",
31487 => "0110110000100111",
31488 => "0110110000101011",
31489 => "0110110000101111",
31490 => "0110110000110010",
31491 => "0110110000110110",
31492 => "0110110000111010",
31493 => "0110110000111110",
31494 => "0110110001000010",
31495 => "0110110001000110",
31496 => "0110110001001010",
31497 => "0110110001001110",
31498 => "0110110001010010",
31499 => "0110110001010110",
31500 => "0110110001011001",
31501 => "0110110001011101",
31502 => "0110110001100001",
31503 => "0110110001100101",
31504 => "0110110001101001",
31505 => "0110110001101101",
31506 => "0110110001110001",
31507 => "0110110001110101",
31508 => "0110110001111001",
31509 => "0110110001111101",
31510 => "0110110010000001",
31511 => "0110110010000100",
31512 => "0110110010001000",
31513 => "0110110010001100",
31514 => "0110110010010000",
31515 => "0110110010010100",
31516 => "0110110010011000",
31517 => "0110110010011100",
31518 => "0110110010100000",
31519 => "0110110010100100",
31520 => "0110110010101000",
31521 => "0110110010101100",
31522 => "0110110010101111",
31523 => "0110110010110011",
31524 => "0110110010110111",
31525 => "0110110010111011",
31526 => "0110110010111111",
31527 => "0110110011000011",
31528 => "0110110011000111",
31529 => "0110110011001011",
31530 => "0110110011001111",
31531 => "0110110011010011",
31532 => "0110110011010111",
31533 => "0110110011011010",
31534 => "0110110011011110",
31535 => "0110110011100010",
31536 => "0110110011100110",
31537 => "0110110011101010",
31538 => "0110110011101110",
31539 => "0110110011110010",
31540 => "0110110011110110",
31541 => "0110110011111010",
31542 => "0110110011111110",
31543 => "0110110100000010",
31544 => "0110110100000101",
31545 => "0110110100001001",
31546 => "0110110100001101",
31547 => "0110110100010001",
31548 => "0110110100010101",
31549 => "0110110100011001",
31550 => "0110110100011101",
31551 => "0110110100100001",
31552 => "0110110100100101",
31553 => "0110110100101001",
31554 => "0110110100101101",
31555 => "0110110100110001",
31556 => "0110110100110100",
31557 => "0110110100111000",
31558 => "0110110100111100",
31559 => "0110110101000000",
31560 => "0110110101000100",
31561 => "0110110101001000",
31562 => "0110110101001100",
31563 => "0110110101010000",
31564 => "0110110101010100",
31565 => "0110110101011000",
31566 => "0110110101011100",
31567 => "0110110101100000",
31568 => "0110110101100011",
31569 => "0110110101100111",
31570 => "0110110101101011",
31571 => "0110110101101111",
31572 => "0110110101110011",
31573 => "0110110101110111",
31574 => "0110110101111011",
31575 => "0110110101111111",
31576 => "0110110110000011",
31577 => "0110110110000111",
31578 => "0110110110001011",
31579 => "0110110110001111",
31580 => "0110110110010010",
31581 => "0110110110010110",
31582 => "0110110110011010",
31583 => "0110110110011110",
31584 => "0110110110100010",
31585 => "0110110110100110",
31586 => "0110110110101010",
31587 => "0110110110101110",
31588 => "0110110110110010",
31589 => "0110110110110110",
31590 => "0110110110111010",
31591 => "0110110110111110",
31592 => "0110110111000001",
31593 => "0110110111000101",
31594 => "0110110111001001",
31595 => "0110110111001101",
31596 => "0110110111010001",
31597 => "0110110111010101",
31598 => "0110110111011001",
31599 => "0110110111011101",
31600 => "0110110111100001",
31601 => "0110110111100101",
31602 => "0110110111101001",
31603 => "0110110111101101",
31604 => "0110110111110000",
31605 => "0110110111110100",
31606 => "0110110111111000",
31607 => "0110110111111100",
31608 => "0110111000000000",
31609 => "0110111000000100",
31610 => "0110111000001000",
31611 => "0110111000001100",
31612 => "0110111000010000",
31613 => "0110111000010100",
31614 => "0110111000011000",
31615 => "0110111000011100",
31616 => "0110111000100000",
31617 => "0110111000100011",
31618 => "0110111000100111",
31619 => "0110111000101011",
31620 => "0110111000101111",
31621 => "0110111000110011",
31622 => "0110111000110111",
31623 => "0110111000111011",
31624 => "0110111000111111",
31625 => "0110111001000011",
31626 => "0110111001000111",
31627 => "0110111001001011",
31628 => "0110111001001111",
31629 => "0110111001010011",
31630 => "0110111001010110",
31631 => "0110111001011010",
31632 => "0110111001011110",
31633 => "0110111001100010",
31634 => "0110111001100110",
31635 => "0110111001101010",
31636 => "0110111001101110",
31637 => "0110111001110010",
31638 => "0110111001110110",
31639 => "0110111001111010",
31640 => "0110111001111110",
31641 => "0110111010000010",
31642 => "0110111010000110",
31643 => "0110111010001001",
31644 => "0110111010001101",
31645 => "0110111010010001",
31646 => "0110111010010101",
31647 => "0110111010011001",
31648 => "0110111010011101",
31649 => "0110111010100001",
31650 => "0110111010100101",
31651 => "0110111010101001",
31652 => "0110111010101101",
31653 => "0110111010110001",
31654 => "0110111010110101",
31655 => "0110111010111001",
31656 => "0110111010111101",
31657 => "0110111011000000",
31658 => "0110111011000100",
31659 => "0110111011001000",
31660 => "0110111011001100",
31661 => "0110111011010000",
31662 => "0110111011010100",
31663 => "0110111011011000",
31664 => "0110111011011100",
31665 => "0110111011100000",
31666 => "0110111011100100",
31667 => "0110111011101000",
31668 => "0110111011101100",
31669 => "0110111011110000",
31670 => "0110111011110100",
31671 => "0110111011110111",
31672 => "0110111011111011",
31673 => "0110111011111111",
31674 => "0110111100000011",
31675 => "0110111100000111",
31676 => "0110111100001011",
31677 => "0110111100001111",
31678 => "0110111100010011",
31679 => "0110111100010111",
31680 => "0110111100011011",
31681 => "0110111100011111",
31682 => "0110111100100011",
31683 => "0110111100100111",
31684 => "0110111100101011",
31685 => "0110111100101110",
31686 => "0110111100110010",
31687 => "0110111100110110",
31688 => "0110111100111010",
31689 => "0110111100111110",
31690 => "0110111101000010",
31691 => "0110111101000110",
31692 => "0110111101001010",
31693 => "0110111101001110",
31694 => "0110111101010010",
31695 => "0110111101010110",
31696 => "0110111101011010",
31697 => "0110111101011110",
31698 => "0110111101100010",
31699 => "0110111101100110",
31700 => "0110111101101001",
31701 => "0110111101101101",
31702 => "0110111101110001",
31703 => "0110111101110101",
31704 => "0110111101111001",
31705 => "0110111101111101",
31706 => "0110111110000001",
31707 => "0110111110000101",
31708 => "0110111110001001",
31709 => "0110111110001101",
31710 => "0110111110010001",
31711 => "0110111110010101",
31712 => "0110111110011001",
31713 => "0110111110011101",
31714 => "0110111110100001",
31715 => "0110111110100100",
31716 => "0110111110101000",
31717 => "0110111110101100",
31718 => "0110111110110000",
31719 => "0110111110110100",
31720 => "0110111110111000",
31721 => "0110111110111100",
31722 => "0110111111000000",
31723 => "0110111111000100",
31724 => "0110111111001000",
31725 => "0110111111001100",
31726 => "0110111111010000",
31727 => "0110111111010100",
31728 => "0110111111011000",
31729 => "0110111111011100",
31730 => "0110111111011111",
31731 => "0110111111100011",
31732 => "0110111111100111",
31733 => "0110111111101011",
31734 => "0110111111101111",
31735 => "0110111111110011",
31736 => "0110111111110111",
31737 => "0110111111111011",
31738 => "0110111111111111",
31739 => "0111000000000011",
31740 => "0111000000000111",
31741 => "0111000000001011",
31742 => "0111000000001111",
31743 => "0111000000010011",
31744 => "0111000000010111",
31745 => "0111000000011011",
31746 => "0111000000011110",
31747 => "0111000000100010",
31748 => "0111000000100110",
31749 => "0111000000101010",
31750 => "0111000000101110",
31751 => "0111000000110010",
31752 => "0111000000110110",
31753 => "0111000000111010",
31754 => "0111000000111110",
31755 => "0111000001000010",
31756 => "0111000001000110",
31757 => "0111000001001010",
31758 => "0111000001001110",
31759 => "0111000001010010",
31760 => "0111000001010110",
31761 => "0111000001011010",
31762 => "0111000001011110",
31763 => "0111000001100001",
31764 => "0111000001100101",
31765 => "0111000001101001",
31766 => "0111000001101101",
31767 => "0111000001110001",
31768 => "0111000001110101",
31769 => "0111000001111001",
31770 => "0111000001111101",
31771 => "0111000010000001",
31772 => "0111000010000101",
31773 => "0111000010001001",
31774 => "0111000010001101",
31775 => "0111000010010001",
31776 => "0111000010010101",
31777 => "0111000010011001",
31778 => "0111000010011101",
31779 => "0111000010100001",
31780 => "0111000010100100",
31781 => "0111000010101000",
31782 => "0111000010101100",
31783 => "0111000010110000",
31784 => "0111000010110100",
31785 => "0111000010111000",
31786 => "0111000010111100",
31787 => "0111000011000000",
31788 => "0111000011000100",
31789 => "0111000011001000",
31790 => "0111000011001100",
31791 => "0111000011010000",
31792 => "0111000011010100",
31793 => "0111000011011000",
31794 => "0111000011011100",
31795 => "0111000011100000",
31796 => "0111000011100100",
31797 => "0111000011101000",
31798 => "0111000011101011",
31799 => "0111000011101111",
31800 => "0111000011110011",
31801 => "0111000011110111",
31802 => "0111000011111011",
31803 => "0111000011111111",
31804 => "0111000100000011",
31805 => "0111000100000111",
31806 => "0111000100001011",
31807 => "0111000100001111",
31808 => "0111000100010011",
31809 => "0111000100010111",
31810 => "0111000100011011",
31811 => "0111000100011111",
31812 => "0111000100100011",
31813 => "0111000100100111",
31814 => "0111000100101011",
31815 => "0111000100101111",
31816 => "0111000100110010",
31817 => "0111000100110110",
31818 => "0111000100111010",
31819 => "0111000100111110",
31820 => "0111000101000010",
31821 => "0111000101000110",
31822 => "0111000101001010",
31823 => "0111000101001110",
31824 => "0111000101010010",
31825 => "0111000101010110",
31826 => "0111000101011010",
31827 => "0111000101011110",
31828 => "0111000101100010",
31829 => "0111000101100110",
31830 => "0111000101101010",
31831 => "0111000101101110",
31832 => "0111000101110010",
31833 => "0111000101110110",
31834 => "0111000101111010",
31835 => "0111000101111101",
31836 => "0111000110000001",
31837 => "0111000110000101",
31838 => "0111000110001001",
31839 => "0111000110001101",
31840 => "0111000110010001",
31841 => "0111000110010101",
31842 => "0111000110011001",
31843 => "0111000110011101",
31844 => "0111000110100001",
31845 => "0111000110100101",
31846 => "0111000110101001",
31847 => "0111000110101101",
31848 => "0111000110110001",
31849 => "0111000110110101",
31850 => "0111000110111001",
31851 => "0111000110111101",
31852 => "0111000111000001",
31853 => "0111000111000101",
31854 => "0111000111001001",
31855 => "0111000111001100",
31856 => "0111000111010000",
31857 => "0111000111010100",
31858 => "0111000111011000",
31859 => "0111000111011100",
31860 => "0111000111100000",
31861 => "0111000111100100",
31862 => "0111000111101000",
31863 => "0111000111101100",
31864 => "0111000111110000",
31865 => "0111000111110100",
31866 => "0111000111111000",
31867 => "0111000111111100",
31868 => "0111001000000000",
31869 => "0111001000000100",
31870 => "0111001000001000",
31871 => "0111001000001100",
31872 => "0111001000010000",
31873 => "0111001000010100",
31874 => "0111001000011000",
31875 => "0111001000011100",
31876 => "0111001000011111",
31877 => "0111001000100011",
31878 => "0111001000100111",
31879 => "0111001000101011",
31880 => "0111001000101111",
31881 => "0111001000110011",
31882 => "0111001000110111",
31883 => "0111001000111011",
31884 => "0111001000111111",
31885 => "0111001001000011",
31886 => "0111001001000111",
31887 => "0111001001001011",
31888 => "0111001001001111",
31889 => "0111001001010011",
31890 => "0111001001010111",
31891 => "0111001001011011",
31892 => "0111001001011111",
31893 => "0111001001100011",
31894 => "0111001001100111",
31895 => "0111001001101011",
31896 => "0111001001101111",
31897 => "0111001001110010",
31898 => "0111001001110110",
31899 => "0111001001111010",
31900 => "0111001001111110",
31901 => "0111001010000010",
31902 => "0111001010000110",
31903 => "0111001010001010",
31904 => "0111001010001110",
31905 => "0111001010010010",
31906 => "0111001010010110",
31907 => "0111001010011010",
31908 => "0111001010011110",
31909 => "0111001010100010",
31910 => "0111001010100110",
31911 => "0111001010101010",
31912 => "0111001010101110",
31913 => "0111001010110010",
31914 => "0111001010110110",
31915 => "0111001010111010",
31916 => "0111001010111110",
31917 => "0111001011000010",
31918 => "0111001011000110",
31919 => "0111001011001010",
31920 => "0111001011001101",
31921 => "0111001011010001",
31922 => "0111001011010101",
31923 => "0111001011011001",
31924 => "0111001011011101",
31925 => "0111001011100001",
31926 => "0111001011100101",
31927 => "0111001011101001",
31928 => "0111001011101101",
31929 => "0111001011110001",
31930 => "0111001011110101",
31931 => "0111001011111001",
31932 => "0111001011111101",
31933 => "0111001100000001",
31934 => "0111001100000101",
31935 => "0111001100001001",
31936 => "0111001100001101",
31937 => "0111001100010001",
31938 => "0111001100010101",
31939 => "0111001100011001",
31940 => "0111001100011101",
31941 => "0111001100100001",
31942 => "0111001100100101",
31943 => "0111001100101001",
31944 => "0111001100101101",
31945 => "0111001100110000",
31946 => "0111001100110100",
31947 => "0111001100111000",
31948 => "0111001100111100",
31949 => "0111001101000000",
31950 => "0111001101000100",
31951 => "0111001101001000",
31952 => "0111001101001100",
31953 => "0111001101010000",
31954 => "0111001101010100",
31955 => "0111001101011000",
31956 => "0111001101011100",
31957 => "0111001101100000",
31958 => "0111001101100100",
31959 => "0111001101101000",
31960 => "0111001101101100",
31961 => "0111001101110000",
31962 => "0111001101110100",
31963 => "0111001101111000",
31964 => "0111001101111100",
31965 => "0111001110000000",
31966 => "0111001110000100",
31967 => "0111001110001000",
31968 => "0111001110001100",
31969 => "0111001110010000",
31970 => "0111001110010011",
31971 => "0111001110010111",
31972 => "0111001110011011",
31973 => "0111001110011111",
31974 => "0111001110100011",
31975 => "0111001110100111",
31976 => "0111001110101011",
31977 => "0111001110101111",
31978 => "0111001110110011",
31979 => "0111001110110111",
31980 => "0111001110111011",
31981 => "0111001110111111",
31982 => "0111001111000011",
31983 => "0111001111000111",
31984 => "0111001111001011",
31985 => "0111001111001111",
31986 => "0111001111010011",
31987 => "0111001111010111",
31988 => "0111001111011011",
31989 => "0111001111011111",
31990 => "0111001111100011",
31991 => "0111001111100111",
31992 => "0111001111101011",
31993 => "0111001111101111",
31994 => "0111001111110011",
31995 => "0111001111110111",
31996 => "0111001111111011",
31997 => "0111001111111111",
31998 => "0111010000000010",
31999 => "0111010000000110",
32000 => "0111010000001010",
32001 => "0111010000001110",
32002 => "0111010000010010",
32003 => "0111010000010110",
32004 => "0111010000011010",
32005 => "0111010000011110",
32006 => "0111010000100010",
32007 => "0111010000100110",
32008 => "0111010000101010",
32009 => "0111010000101110",
32010 => "0111010000110010",
32011 => "0111010000110110",
32012 => "0111010000111010",
32013 => "0111010000111110",
32014 => "0111010001000010",
32015 => "0111010001000110",
32016 => "0111010001001010",
32017 => "0111010001001110",
32018 => "0111010001010010",
32019 => "0111010001010110",
32020 => "0111010001011010",
32021 => "0111010001011110",
32022 => "0111010001100010",
32023 => "0111010001100110",
32024 => "0111010001101010",
32025 => "0111010001101110",
32026 => "0111010001110010",
32027 => "0111010001110101",
32028 => "0111010001111001",
32029 => "0111010001111101",
32030 => "0111010010000001",
32031 => "0111010010000101",
32032 => "0111010010001001",
32033 => "0111010010001101",
32034 => "0111010010010001",
32035 => "0111010010010101",
32036 => "0111010010011001",
32037 => "0111010010011101",
32038 => "0111010010100001",
32039 => "0111010010100101",
32040 => "0111010010101001",
32041 => "0111010010101101",
32042 => "0111010010110001",
32043 => "0111010010110101",
32044 => "0111010010111001",
32045 => "0111010010111101",
32046 => "0111010011000001",
32047 => "0111010011000101",
32048 => "0111010011001001",
32049 => "0111010011001101",
32050 => "0111010011010001",
32051 => "0111010011010101",
32052 => "0111010011011001",
32053 => "0111010011011101",
32054 => "0111010011100001",
32055 => "0111010011100101",
32056 => "0111010011101001",
32057 => "0111010011101101",
32058 => "0111010011110001",
32059 => "0111010011110101",
32060 => "0111010011111000",
32061 => "0111010011111100",
32062 => "0111010100000000",
32063 => "0111010100000100",
32064 => "0111010100001000",
32065 => "0111010100001100",
32066 => "0111010100010000",
32067 => "0111010100010100",
32068 => "0111010100011000",
32069 => "0111010100011100",
32070 => "0111010100100000",
32071 => "0111010100100100",
32072 => "0111010100101000",
32073 => "0111010100101100",
32074 => "0111010100110000",
32075 => "0111010100110100",
32076 => "0111010100111000",
32077 => "0111010100111100",
32078 => "0111010101000000",
32079 => "0111010101000100",
32080 => "0111010101001000",
32081 => "0111010101001100",
32082 => "0111010101010000",
32083 => "0111010101010100",
32084 => "0111010101011000",
32085 => "0111010101011100",
32086 => "0111010101100000",
32087 => "0111010101100100",
32088 => "0111010101101000",
32089 => "0111010101101100",
32090 => "0111010101110000",
32091 => "0111010101110100",
32092 => "0111010101111000",
32093 => "0111010101111100",
32094 => "0111010110000000",
32095 => "0111010110000011",
32096 => "0111010110000111",
32097 => "0111010110001011",
32098 => "0111010110001111",
32099 => "0111010110010011",
32100 => "0111010110010111",
32101 => "0111010110011011",
32102 => "0111010110011111",
32103 => "0111010110100011",
32104 => "0111010110100111",
32105 => "0111010110101011",
32106 => "0111010110101111",
32107 => "0111010110110011",
32108 => "0111010110110111",
32109 => "0111010110111011",
32110 => "0111010110111111",
32111 => "0111010111000011",
32112 => "0111010111000111",
32113 => "0111010111001011",
32114 => "0111010111001111",
32115 => "0111010111010011",
32116 => "0111010111010111",
32117 => "0111010111011011",
32118 => "0111010111011111",
32119 => "0111010111100011",
32120 => "0111010111100111",
32121 => "0111010111101011",
32122 => "0111010111101111",
32123 => "0111010111110011",
32124 => "0111010111110111",
32125 => "0111010111111011",
32126 => "0111010111111111",
32127 => "0111011000000011",
32128 => "0111011000000111",
32129 => "0111011000001011",
32130 => "0111011000001111",
32131 => "0111011000010011",
32132 => "0111011000010111",
32133 => "0111011000011011",
32134 => "0111011000011111",
32135 => "0111011000100010",
32136 => "0111011000100110",
32137 => "0111011000101010",
32138 => "0111011000101110",
32139 => "0111011000110010",
32140 => "0111011000110110",
32141 => "0111011000111010",
32142 => "0111011000111110",
32143 => "0111011001000010",
32144 => "0111011001000110",
32145 => "0111011001001010",
32146 => "0111011001001110",
32147 => "0111011001010010",
32148 => "0111011001010110",
32149 => "0111011001011010",
32150 => "0111011001011110",
32151 => "0111011001100010",
32152 => "0111011001100110",
32153 => "0111011001101010",
32154 => "0111011001101110",
32155 => "0111011001110010",
32156 => "0111011001110110",
32157 => "0111011001111010",
32158 => "0111011001111110",
32159 => "0111011010000010",
32160 => "0111011010000110",
32161 => "0111011010001010",
32162 => "0111011010001110",
32163 => "0111011010010010",
32164 => "0111011010010110",
32165 => "0111011010011010",
32166 => "0111011010011110",
32167 => "0111011010100010",
32168 => "0111011010100110",
32169 => "0111011010101010",
32170 => "0111011010101110",
32171 => "0111011010110010",
32172 => "0111011010110110",
32173 => "0111011010111010",
32174 => "0111011010111110",
32175 => "0111011011000010",
32176 => "0111011011000110",
32177 => "0111011011001010",
32178 => "0111011011001110",
32179 => "0111011011010010",
32180 => "0111011011010101",
32181 => "0111011011011001",
32182 => "0111011011011101",
32183 => "0111011011100001",
32184 => "0111011011100101",
32185 => "0111011011101001",
32186 => "0111011011101101",
32187 => "0111011011110001",
32188 => "0111011011110101",
32189 => "0111011011111001",
32190 => "0111011011111101",
32191 => "0111011100000001",
32192 => "0111011100000101",
32193 => "0111011100001001",
32194 => "0111011100001101",
32195 => "0111011100010001",
32196 => "0111011100010101",
32197 => "0111011100011001",
32198 => "0111011100011101",
32199 => "0111011100100001",
32200 => "0111011100100101",
32201 => "0111011100101001",
32202 => "0111011100101101",
32203 => "0111011100110001",
32204 => "0111011100110101",
32205 => "0111011100111001",
32206 => "0111011100111101",
32207 => "0111011101000001",
32208 => "0111011101000101",
32209 => "0111011101001001",
32210 => "0111011101001101",
32211 => "0111011101010001",
32212 => "0111011101010101",
32213 => "0111011101011001",
32214 => "0111011101011101",
32215 => "0111011101100001",
32216 => "0111011101100101",
32217 => "0111011101101001",
32218 => "0111011101101101",
32219 => "0111011101110001",
32220 => "0111011101110101",
32221 => "0111011101111001",
32222 => "0111011101111101",
32223 => "0111011110000001",
32224 => "0111011110000101",
32225 => "0111011110001001",
32226 => "0111011110001101",
32227 => "0111011110010001",
32228 => "0111011110010101",
32229 => "0111011110011001",
32230 => "0111011110011101",
32231 => "0111011110100001",
32232 => "0111011110100101",
32233 => "0111011110101000",
32234 => "0111011110101100",
32235 => "0111011110110000",
32236 => "0111011110110100",
32237 => "0111011110111000",
32238 => "0111011110111100",
32239 => "0111011111000000",
32240 => "0111011111000100",
32241 => "0111011111001000",
32242 => "0111011111001100",
32243 => "0111011111010000",
32244 => "0111011111010100",
32245 => "0111011111011000",
32246 => "0111011111011100",
32247 => "0111011111100000",
32248 => "0111011111100100",
32249 => "0111011111101000",
32250 => "0111011111101100",
32251 => "0111011111110000",
32252 => "0111011111110100",
32253 => "0111011111111000",
32254 => "0111011111111100",
32255 => "0111100000000000",
32256 => "0111100000000100",
32257 => "0111100000001000",
32258 => "0111100000001100",
32259 => "0111100000010000",
32260 => "0111100000010100",
32261 => "0111100000011000",
32262 => "0111100000011100",
32263 => "0111100000100000",
32264 => "0111100000100100",
32265 => "0111100000101000",
32266 => "0111100000101100",
32267 => "0111100000110000",
32268 => "0111100000110100",
32269 => "0111100000111000",
32270 => "0111100000111100",
32271 => "0111100001000000",
32272 => "0111100001000100",
32273 => "0111100001001000",
32274 => "0111100001001100",
32275 => "0111100001010000",
32276 => "0111100001010100",
32277 => "0111100001011000",
32278 => "0111100001011100",
32279 => "0111100001100000",
32280 => "0111100001100100",
32281 => "0111100001101000",
32282 => "0111100001101100",
32283 => "0111100001110000",
32284 => "0111100001110100",
32285 => "0111100001111000",
32286 => "0111100001111100",
32287 => "0111100010000000",
32288 => "0111100010000100",
32289 => "0111100010001000",
32290 => "0111100010001100",
32291 => "0111100010010000",
32292 => "0111100010010100",
32293 => "0111100010011000",
32294 => "0111100010011100",
32295 => "0111100010100000",
32296 => "0111100010100100",
32297 => "0111100010101000",
32298 => "0111100010101100",
32299 => "0111100010110000",
32300 => "0111100010110011",
32301 => "0111100010110111",
32302 => "0111100010111011",
32303 => "0111100010111111",
32304 => "0111100011000011",
32305 => "0111100011000111",
32306 => "0111100011001011",
32307 => "0111100011001111",
32308 => "0111100011010011",
32309 => "0111100011010111",
32310 => "0111100011011011",
32311 => "0111100011011111",
32312 => "0111100011100011",
32313 => "0111100011100111",
32314 => "0111100011101011",
32315 => "0111100011101111",
32316 => "0111100011110011",
32317 => "0111100011110111",
32318 => "0111100011111011",
32319 => "0111100011111111",
32320 => "0111100100000011",
32321 => "0111100100000111",
32322 => "0111100100001011",
32323 => "0111100100001111",
32324 => "0111100100010011",
32325 => "0111100100010111",
32326 => "0111100100011011",
32327 => "0111100100011111",
32328 => "0111100100100011",
32329 => "0111100100100111",
32330 => "0111100100101011",
32331 => "0111100100101111",
32332 => "0111100100110011",
32333 => "0111100100110111",
32334 => "0111100100111011",
32335 => "0111100100111111",
32336 => "0111100101000011",
32337 => "0111100101000111",
32338 => "0111100101001011",
32339 => "0111100101001111",
32340 => "0111100101010011",
32341 => "0111100101010111",
32342 => "0111100101011011",
32343 => "0111100101011111",
32344 => "0111100101100011",
32345 => "0111100101100111",
32346 => "0111100101101011",
32347 => "0111100101101111",
32348 => "0111100101110011",
32349 => "0111100101110111",
32350 => "0111100101111011",
32351 => "0111100101111111",
32352 => "0111100110000011",
32353 => "0111100110000111",
32354 => "0111100110001011",
32355 => "0111100110001111",
32356 => "0111100110010011",
32357 => "0111100110010111",
32358 => "0111100110011011",
32359 => "0111100110011111",
32360 => "0111100110100011",
32361 => "0111100110100111",
32362 => "0111100110101011",
32363 => "0111100110101111",
32364 => "0111100110110011",
32365 => "0111100110110111",
32366 => "0111100110111011",
32367 => "0111100110111111",
32368 => "0111100111000011",
32369 => "0111100111000111",
32370 => "0111100111001011",
32371 => "0111100111001111",
32372 => "0111100111010011",
32373 => "0111100111010111",
32374 => "0111100111011011",
32375 => "0111100111011111",
32376 => "0111100111100011",
32377 => "0111100111100111",
32378 => "0111100111101011",
32379 => "0111100111101111",
32380 => "0111100111110011",
32381 => "0111100111110111",
32382 => "0111100111111011",
32383 => "0111100111111111",
32384 => "0111101000000011",
32385 => "0111101000000111",
32386 => "0111101000001011",
32387 => "0111101000001111",
32388 => "0111101000010011",
32389 => "0111101000010111",
32390 => "0111101000011011",
32391 => "0111101000011111",
32392 => "0111101000100011",
32393 => "0111101000100111",
32394 => "0111101000101011",
32395 => "0111101000101111",
32396 => "0111101000110010",
32397 => "0111101000110110",
32398 => "0111101000111010",
32399 => "0111101000111110",
32400 => "0111101001000010",
32401 => "0111101001000110",
32402 => "0111101001001010",
32403 => "0111101001001110",
32404 => "0111101001010010",
32405 => "0111101001010110",
32406 => "0111101001011010",
32407 => "0111101001011110",
32408 => "0111101001100010",
32409 => "0111101001100110",
32410 => "0111101001101010",
32411 => "0111101001101110",
32412 => "0111101001110010",
32413 => "0111101001110110",
32414 => "0111101001111010",
32415 => "0111101001111110",
32416 => "0111101010000010",
32417 => "0111101010000110",
32418 => "0111101010001010",
32419 => "0111101010001110",
32420 => "0111101010010010",
32421 => "0111101010010110",
32422 => "0111101010011010",
32423 => "0111101010011110",
32424 => "0111101010100010",
32425 => "0111101010100110",
32426 => "0111101010101010",
32427 => "0111101010101110",
32428 => "0111101010110010",
32429 => "0111101010110110",
32430 => "0111101010111010",
32431 => "0111101010111110",
32432 => "0111101011000010",
32433 => "0111101011000110",
32434 => "0111101011001010",
32435 => "0111101011001110",
32436 => "0111101011010010",
32437 => "0111101011010110",
32438 => "0111101011011010",
32439 => "0111101011011110",
32440 => "0111101011100010",
32441 => "0111101011100110",
32442 => "0111101011101010",
32443 => "0111101011101110",
32444 => "0111101011110010",
32445 => "0111101011110110",
32446 => "0111101011111010",
32447 => "0111101011111110",
32448 => "0111101100000010",
32449 => "0111101100000110",
32450 => "0111101100001010",
32451 => "0111101100001110",
32452 => "0111101100010010",
32453 => "0111101100010110",
32454 => "0111101100011010",
32455 => "0111101100011110",
32456 => "0111101100100010",
32457 => "0111101100100110",
32458 => "0111101100101010",
32459 => "0111101100101110",
32460 => "0111101100110010",
32461 => "0111101100110110",
32462 => "0111101100111010",
32463 => "0111101100111110",
32464 => "0111101101000010",
32465 => "0111101101000110",
32466 => "0111101101001010",
32467 => "0111101101001110",
32468 => "0111101101010010",
32469 => "0111101101010110",
32470 => "0111101101011010",
32471 => "0111101101011110",
32472 => "0111101101100010",
32473 => "0111101101100110",
32474 => "0111101101101010",
32475 => "0111101101101110",
32476 => "0111101101110010",
32477 => "0111101101110110",
32478 => "0111101101111010",
32479 => "0111101101111110",
32480 => "0111101110000010",
32481 => "0111101110000110",
32482 => "0111101110001010",
32483 => "0111101110001110",
32484 => "0111101110010010",
32485 => "0111101110010110",
32486 => "0111101110011010",
32487 => "0111101110011110",
32488 => "0111101110100010",
32489 => "0111101110100110",
32490 => "0111101110101010",
32491 => "0111101110101110",
32492 => "0111101110110010",
32493 => "0111101110110110",
32494 => "0111101110111010",
32495 => "0111101110111110",
32496 => "0111101111000010",
32497 => "0111101111000110",
32498 => "0111101111001010",
32499 => "0111101111001110",
32500 => "0111101111010010",
32501 => "0111101111010110",
32502 => "0111101111011010",
32503 => "0111101111011110",
32504 => "0111101111100010",
32505 => "0111101111100110",
32506 => "0111101111101010",
32507 => "0111101111101110",
32508 => "0111101111110010",
32509 => "0111101111110110",
32510 => "0111101111111010",
32511 => "0111101111111110",
32512 => "0111110000000010",
32513 => "0111110000000110",
32514 => "0111110000001010",
32515 => "0111110000001110",
32516 => "0111110000010010",
32517 => "0111110000010110",
32518 => "0111110000011010",
32519 => "0111110000011110",
32520 => "0111110000100010",
32521 => "0111110000100110",
32522 => "0111110000101010",
32523 => "0111110000101110",
32524 => "0111110000110010",
32525 => "0111110000110110",
32526 => "0111110000111010",
32527 => "0111110000111110",
32528 => "0111110001000010",
32529 => "0111110001000110",
32530 => "0111110001001010",
32531 => "0111110001001110",
32532 => "0111110001010010",
32533 => "0111110001010110",
32534 => "0111110001011010",
32535 => "0111110001011110",
32536 => "0111110001100010",
32537 => "0111110001100110",
32538 => "0111110001101010",
32539 => "0111110001101110",
32540 => "0111110001110010",
32541 => "0111110001110110",
32542 => "0111110001111010",
32543 => "0111110001111110",
32544 => "0111110010000010",
32545 => "0111110010000110",
32546 => "0111110010001010",
32547 => "0111110010001110",
32548 => "0111110010010010",
32549 => "0111110010010110",
32550 => "0111110010011010",
32551 => "0111110010011110",
32552 => "0111110010100010",
32553 => "0111110010100110",
32554 => "0111110010101010",
32555 => "0111110010101110",
32556 => "0111110010110010",
32557 => "0111110010110110",
32558 => "0111110010111010",
32559 => "0111110010111110",
32560 => "0111110011000010",
32561 => "0111110011000110",
32562 => "0111110011001010",
32563 => "0111110011001110",
32564 => "0111110011010010",
32565 => "0111110011010110",
32566 => "0111110011011010",
32567 => "0111110011011110",
32568 => "0111110011100010",
32569 => "0111110011100110",
32570 => "0111110011101010",
32571 => "0111110011101110",
32572 => "0111110011110010",
32573 => "0111110011110110",
32574 => "0111110011111010",
32575 => "0111110011111110",
32576 => "0111110100000010",
32577 => "0111110100000110",
32578 => "0111110100001010",
32579 => "0111110100001110",
32580 => "0111110100010010",
32581 => "0111110100010110",
32582 => "0111110100011010",
32583 => "0111110100011110",
32584 => "0111110100100010",
32585 => "0111110100100110",
32586 => "0111110100101010",
32587 => "0111110100101110",
32588 => "0111110100110010",
32589 => "0111110100110110",
32590 => "0111110100111010",
32591 => "0111110100111110",
32592 => "0111110101000010",
32593 => "0111110101000110",
32594 => "0111110101001010",
32595 => "0111110101001110",
32596 => "0111110101010010",
32597 => "0111110101010110",
32598 => "0111110101011010",
32599 => "0111110101011110",
32600 => "0111110101100010",
32601 => "0111110101100110",
32602 => "0111110101101010",
32603 => "0111110101101110",
32604 => "0111110101110010",
32605 => "0111110101110110",
32606 => "0111110101111010",
32607 => "0111110101111110",
32608 => "0111110110000010",
32609 => "0111110110000110",
32610 => "0111110110001010",
32611 => "0111110110001110",
32612 => "0111110110010010",
32613 => "0111110110010110",
32614 => "0111110110011010",
32615 => "0111110110011110",
32616 => "0111110110100010",
32617 => "0111110110100110",
32618 => "0111110110101010",
32619 => "0111110110101110",
32620 => "0111110110110010",
32621 => "0111110110110110",
32622 => "0111110110111010",
32623 => "0111110110111110",
32624 => "0111110111000010",
32625 => "0111110111000110",
32626 => "0111110111001010",
32627 => "0111110111001110",
32628 => "0111110111010010",
32629 => "0111110111010110",
32630 => "0111110111011010",
32631 => "0111110111011110",
32632 => "0111110111100010",
32633 => "0111110111100110",
32634 => "0111110111101010",
32635 => "0111110111101110",
32636 => "0111110111110010",
32637 => "0111110111110110",
32638 => "0111110111111010",
32639 => "0111110111111110",
32640 => "0111111000000010",
32641 => "0111111000000110",
32642 => "0111111000001010",
32643 => "0111111000001110",
32644 => "0111111000010010",
32645 => "0111111000010110",
32646 => "0111111000011010",
32647 => "0111111000011110",
32648 => "0111111000100010",
32649 => "0111111000100110",
32650 => "0111111000101010",
32651 => "0111111000101110",
32652 => "0111111000110010",
32653 => "0111111000110110",
32654 => "0111111000111010",
32655 => "0111111000111110",
32656 => "0111111001000010",
32657 => "0111111001000110",
32658 => "0111111001001010",
32659 => "0111111001001110",
32660 => "0111111001010010",
32661 => "0111111001010110",
32662 => "0111111001011010",
32663 => "0111111001011110",
32664 => "0111111001100010",
32665 => "0111111001100110",
32666 => "0111111001101010",
32667 => "0111111001101110",
32668 => "0111111001110010",
32669 => "0111111001110110",
32670 => "0111111001111010",
32671 => "0111111001111110",
32672 => "0111111010000010",
32673 => "0111111010000110",
32674 => "0111111010001010",
32675 => "0111111010001110",
32676 => "0111111010010010",
32677 => "0111111010010110",
32678 => "0111111010011010",
32679 => "0111111010011110",
32680 => "0111111010100010",
32681 => "0111111010100110",
32682 => "0111111010101010",
32683 => "0111111010101110",
32684 => "0111111010110010",
32685 => "0111111010110110",
32686 => "0111111010111010",
32687 => "0111111010111110",
32688 => "0111111011000010",
32689 => "0111111011000110",
32690 => "0111111011001010",
32691 => "0111111011001110",
32692 => "0111111011010010",
32693 => "0111111011010110",
32694 => "0111111011011010",
32695 => "0111111011011110",
32696 => "0111111011100010",
32697 => "0111111011100110",
32698 => "0111111011101010",
32699 => "0111111011101110",
32700 => "0111111011110010",
32701 => "0111111011110110",
32702 => "0111111011111010",
32703 => "0111111011111110",
32704 => "0111111100000010",
32705 => "0111111100000110",
32706 => "0111111100001010",
32707 => "0111111100001110",
32708 => "0111111100010010",
32709 => "0111111100010110",
32710 => "0111111100011010",
32711 => "0111111100011110",
32712 => "0111111100100010",
32713 => "0111111100100101",
32714 => "0111111100101001",
32715 => "0111111100101101",
32716 => "0111111100110001",
32717 => "0111111100110101",
32718 => "0111111100111001",
32719 => "0111111100111101",
32720 => "0111111101000001",
32721 => "0111111101000101",
32722 => "0111111101001001",
32723 => "0111111101001101",
32724 => "0111111101010001",
32725 => "0111111101010101",
32726 => "0111111101011001",
32727 => "0111111101011101",
32728 => "0111111101100001",
32729 => "0111111101100101",
32730 => "0111111101101001",
32731 => "0111111101101101",
32732 => "0111111101110001",
32733 => "0111111101110101",
32734 => "0111111101111001",
32735 => "0111111101111101",
32736 => "0111111110000001",
32737 => "0111111110000101",
32738 => "0111111110001001",
32739 => "0111111110001101",
32740 => "0111111110010001",
32741 => "0111111110010101",
32742 => "0111111110011001",
32743 => "0111111110011101",
32744 => "0111111110100001",
32745 => "0111111110100101",
32746 => "0111111110101001",
32747 => "0111111110101101",
32748 => "0111111110110001",
32749 => "0111111110110101",
32750 => "0111111110111001",
32751 => "0111111110111101",
32752 => "0111111111000001",
32753 => "0111111111000101",
32754 => "0111111111001001",
32755 => "0111111111001101",
32756 => "0111111111010001",
32757 => "0111111111010101",
32758 => "0111111111011001",
32759 => "0111111111011101",
32760 => "0111111111100001",
32761 => "0111111111100101",
32762 => "0111111111101001",
32763 => "0111111111101101",
32764 => "0111111111110001",
32765 => "0111111111110101",
32766 => "0111111111111001",
32767 => "0111111111111101",
32768 => "1000000000000010",
32769 => "1000000000000110",
32770 => "1000000000001010",
32771 => "1000000000001110",
32772 => "1000000000010010",
32773 => "1000000000010110",
32774 => "1000000000011010",
32775 => "1000000000011110",
32776 => "1000000000100010",
32777 => "1000000000100110",
32778 => "1000000000101010",
32779 => "1000000000101110",
32780 => "1000000000110010",
32781 => "1000000000110110",
32782 => "1000000000111010",
32783 => "1000000000111110",
32784 => "1000000001000010",
32785 => "1000000001000110",
32786 => "1000000001001010",
32787 => "1000000001001110",
32788 => "1000000001010010",
32789 => "1000000001010110",
32790 => "1000000001011010",
32791 => "1000000001011110",
32792 => "1000000001100010",
32793 => "1000000001100110",
32794 => "1000000001101010",
32795 => "1000000001101110",
32796 => "1000000001110010",
32797 => "1000000001110110",
32798 => "1000000001111010",
32799 => "1000000001111110",
32800 => "1000000010000010",
32801 => "1000000010000110",
32802 => "1000000010001010",
32803 => "1000000010001110",
32804 => "1000000010010010",
32805 => "1000000010010110",
32806 => "1000000010011010",
32807 => "1000000010011110",
32808 => "1000000010100010",
32809 => "1000000010100110",
32810 => "1000000010101010",
32811 => "1000000010101110",
32812 => "1000000010110010",
32813 => "1000000010110110",
32814 => "1000000010111010",
32815 => "1000000010111110",
32816 => "1000000011000010",
32817 => "1000000011000110",
32818 => "1000000011001010",
32819 => "1000000011001110",
32820 => "1000000011010010",
32821 => "1000000011010110",
32822 => "1000000011011010",
32823 => "1000000011011101",
32824 => "1000000011100001",
32825 => "1000000011100101",
32826 => "1000000011101001",
32827 => "1000000011101101",
32828 => "1000000011110001",
32829 => "1000000011110101",
32830 => "1000000011111001",
32831 => "1000000011111101",
32832 => "1000000100000001",
32833 => "1000000100000101",
32834 => "1000000100001001",
32835 => "1000000100001101",
32836 => "1000000100010001",
32837 => "1000000100010101",
32838 => "1000000100011001",
32839 => "1000000100011101",
32840 => "1000000100100001",
32841 => "1000000100100101",
32842 => "1000000100101001",
32843 => "1000000100101101",
32844 => "1000000100110001",
32845 => "1000000100110101",
32846 => "1000000100111001",
32847 => "1000000100111101",
32848 => "1000000101000001",
32849 => "1000000101000101",
32850 => "1000000101001001",
32851 => "1000000101001101",
32852 => "1000000101010001",
32853 => "1000000101010101",
32854 => "1000000101011001",
32855 => "1000000101011101",
32856 => "1000000101100001",
32857 => "1000000101100101",
32858 => "1000000101101001",
32859 => "1000000101101101",
32860 => "1000000101110001",
32861 => "1000000101110101",
32862 => "1000000101111001",
32863 => "1000000101111101",
32864 => "1000000110000001",
32865 => "1000000110000101",
32866 => "1000000110001001",
32867 => "1000000110001101",
32868 => "1000000110010001",
32869 => "1000000110010101",
32870 => "1000000110011001",
32871 => "1000000110011101",
32872 => "1000000110100001",
32873 => "1000000110100101",
32874 => "1000000110101001",
32875 => "1000000110101101",
32876 => "1000000110110001",
32877 => "1000000110110101",
32878 => "1000000110111001",
32879 => "1000000110111101",
32880 => "1000000111000001",
32881 => "1000000111000101",
32882 => "1000000111001001",
32883 => "1000000111001101",
32884 => "1000000111010001",
32885 => "1000000111010101",
32886 => "1000000111011001",
32887 => "1000000111011101",
32888 => "1000000111100001",
32889 => "1000000111100101",
32890 => "1000000111101001",
32891 => "1000000111101101",
32892 => "1000000111110001",
32893 => "1000000111110101",
32894 => "1000000111111001",
32895 => "1000000111111101",
32896 => "1000001000000001",
32897 => "1000001000000101",
32898 => "1000001000001001",
32899 => "1000001000001101",
32900 => "1000001000010001",
32901 => "1000001000010101",
32902 => "1000001000011001",
32903 => "1000001000011101",
32904 => "1000001000100001",
32905 => "1000001000100101",
32906 => "1000001000101001",
32907 => "1000001000101101",
32908 => "1000001000110001",
32909 => "1000001000110101",
32910 => "1000001000111001",
32911 => "1000001000111101",
32912 => "1000001001000001",
32913 => "1000001001000101",
32914 => "1000001001001001",
32915 => "1000001001001101",
32916 => "1000001001010001",
32917 => "1000001001010101",
32918 => "1000001001011001",
32919 => "1000001001011101",
32920 => "1000001001100001",
32921 => "1000001001100101",
32922 => "1000001001101001",
32923 => "1000001001101101",
32924 => "1000001001110001",
32925 => "1000001001110101",
32926 => "1000001001111001",
32927 => "1000001001111101",
32928 => "1000001010000001",
32929 => "1000001010000101",
32930 => "1000001010001001",
32931 => "1000001010001101",
32932 => "1000001010010001",
32933 => "1000001010010101",
32934 => "1000001010011001",
32935 => "1000001010011101",
32936 => "1000001010100001",
32937 => "1000001010100101",
32938 => "1000001010101001",
32939 => "1000001010101101",
32940 => "1000001010110001",
32941 => "1000001010110101",
32942 => "1000001010111001",
32943 => "1000001010111101",
32944 => "1000001011000001",
32945 => "1000001011000101",
32946 => "1000001011001001",
32947 => "1000001011001101",
32948 => "1000001011010001",
32949 => "1000001011010101",
32950 => "1000001011011001",
32951 => "1000001011011101",
32952 => "1000001011100001",
32953 => "1000001011100101",
32954 => "1000001011101001",
32955 => "1000001011101101",
32956 => "1000001011110001",
32957 => "1000001011110101",
32958 => "1000001011111001",
32959 => "1000001011111101",
32960 => "1000001100000001",
32961 => "1000001100000101",
32962 => "1000001100001001",
32963 => "1000001100001101",
32964 => "1000001100010001",
32965 => "1000001100010101",
32966 => "1000001100011001",
32967 => "1000001100011101",
32968 => "1000001100100001",
32969 => "1000001100100101",
32970 => "1000001100101001",
32971 => "1000001100101101",
32972 => "1000001100110001",
32973 => "1000001100110101",
32974 => "1000001100111001",
32975 => "1000001100111101",
32976 => "1000001101000001",
32977 => "1000001101000101",
32978 => "1000001101001001",
32979 => "1000001101001101",
32980 => "1000001101010001",
32981 => "1000001101010101",
32982 => "1000001101011001",
32983 => "1000001101011101",
32984 => "1000001101100001",
32985 => "1000001101100101",
32986 => "1000001101101001",
32987 => "1000001101101101",
32988 => "1000001101110001",
32989 => "1000001101110101",
32990 => "1000001101111001",
32991 => "1000001101111101",
32992 => "1000001110000001",
32993 => "1000001110000101",
32994 => "1000001110001001",
32995 => "1000001110001101",
32996 => "1000001110010001",
32997 => "1000001110010101",
32998 => "1000001110011001",
32999 => "1000001110011101",
33000 => "1000001110100001",
33001 => "1000001110100101",
33002 => "1000001110101001",
33003 => "1000001110101101",
33004 => "1000001110110001",
33005 => "1000001110110101",
33006 => "1000001110111001",
33007 => "1000001110111101",
33008 => "1000001111000001",
33009 => "1000001111000101",
33010 => "1000001111001001",
33011 => "1000001111001101",
33012 => "1000001111010001",
33013 => "1000001111010101",
33014 => "1000001111011001",
33015 => "1000001111011101",
33016 => "1000001111100001",
33017 => "1000001111100101",
33018 => "1000001111101001",
33019 => "1000001111101101",
33020 => "1000001111110001",
33021 => "1000001111110101",
33022 => "1000001111111001",
33023 => "1000001111111101",
33024 => "1000010000000001",
33025 => "1000010000000101",
33026 => "1000010000001001",
33027 => "1000010000001101",
33028 => "1000010000010001",
33029 => "1000010000010101",
33030 => "1000010000011001",
33031 => "1000010000011101",
33032 => "1000010000100001",
33033 => "1000010000100101",
33034 => "1000010000101001",
33035 => "1000010000101101",
33036 => "1000010000110001",
33037 => "1000010000110101",
33038 => "1000010000111001",
33039 => "1000010000111101",
33040 => "1000010001000001",
33041 => "1000010001000101",
33042 => "1000010001001001",
33043 => "1000010001001101",
33044 => "1000010001010001",
33045 => "1000010001010101",
33046 => "1000010001011001",
33047 => "1000010001011101",
33048 => "1000010001100001",
33049 => "1000010001100101",
33050 => "1000010001101001",
33051 => "1000010001101101",
33052 => "1000010001110001",
33053 => "1000010001110101",
33054 => "1000010001111001",
33055 => "1000010001111101",
33056 => "1000010010000001",
33057 => "1000010010000101",
33058 => "1000010010001001",
33059 => "1000010010001101",
33060 => "1000010010010001",
33061 => "1000010010010101",
33062 => "1000010010011001",
33063 => "1000010010011101",
33064 => "1000010010100001",
33065 => "1000010010100101",
33066 => "1000010010101001",
33067 => "1000010010101101",
33068 => "1000010010110001",
33069 => "1000010010110101",
33070 => "1000010010111001",
33071 => "1000010010111101",
33072 => "1000010011000001",
33073 => "1000010011000101",
33074 => "1000010011001001",
33075 => "1000010011001101",
33076 => "1000010011010001",
33077 => "1000010011010101",
33078 => "1000010011011001",
33079 => "1000010011011101",
33080 => "1000010011100001",
33081 => "1000010011100101",
33082 => "1000010011101001",
33083 => "1000010011101101",
33084 => "1000010011110001",
33085 => "1000010011110101",
33086 => "1000010011111001",
33087 => "1000010011111101",
33088 => "1000010100000001",
33089 => "1000010100000101",
33090 => "1000010100001001",
33091 => "1000010100001101",
33092 => "1000010100010001",
33093 => "1000010100010101",
33094 => "1000010100011001",
33095 => "1000010100011101",
33096 => "1000010100100001",
33097 => "1000010100100101",
33098 => "1000010100101001",
33099 => "1000010100101101",
33100 => "1000010100110001",
33101 => "1000010100110101",
33102 => "1000010100111001",
33103 => "1000010100111101",
33104 => "1000010101000001",
33105 => "1000010101000101",
33106 => "1000010101001001",
33107 => "1000010101001101",
33108 => "1000010101010001",
33109 => "1000010101010101",
33110 => "1000010101011001",
33111 => "1000010101011101",
33112 => "1000010101100001",
33113 => "1000010101100101",
33114 => "1000010101101001",
33115 => "1000010101101101",
33116 => "1000010101110001",
33117 => "1000010101110101",
33118 => "1000010101111001",
33119 => "1000010101111101",
33120 => "1000010110000001",
33121 => "1000010110000101",
33122 => "1000010110001001",
33123 => "1000010110001101",
33124 => "1000010110010001",
33125 => "1000010110010101",
33126 => "1000010110011001",
33127 => "1000010110011101",
33128 => "1000010110100001",
33129 => "1000010110100101",
33130 => "1000010110101001",
33131 => "1000010110101101",
33132 => "1000010110110001",
33133 => "1000010110110101",
33134 => "1000010110111001",
33135 => "1000010110111101",
33136 => "1000010111000001",
33137 => "1000010111000101",
33138 => "1000010111001001",
33139 => "1000010111001101",
33140 => "1000010111010000",
33141 => "1000010111010100",
33142 => "1000010111011000",
33143 => "1000010111011100",
33144 => "1000010111100000",
33145 => "1000010111100100",
33146 => "1000010111101000",
33147 => "1000010111101100",
33148 => "1000010111110000",
33149 => "1000010111110100",
33150 => "1000010111111000",
33151 => "1000010111111100",
33152 => "1000011000000000",
33153 => "1000011000000100",
33154 => "1000011000001000",
33155 => "1000011000001100",
33156 => "1000011000010000",
33157 => "1000011000010100",
33158 => "1000011000011000",
33159 => "1000011000011100",
33160 => "1000011000100000",
33161 => "1000011000100100",
33162 => "1000011000101000",
33163 => "1000011000101100",
33164 => "1000011000110000",
33165 => "1000011000110100",
33166 => "1000011000111000",
33167 => "1000011000111100",
33168 => "1000011001000000",
33169 => "1000011001000100",
33170 => "1000011001001000",
33171 => "1000011001001100",
33172 => "1000011001010000",
33173 => "1000011001010100",
33174 => "1000011001011000",
33175 => "1000011001011100",
33176 => "1000011001100000",
33177 => "1000011001100100",
33178 => "1000011001101000",
33179 => "1000011001101100",
33180 => "1000011001110000",
33181 => "1000011001110100",
33182 => "1000011001111000",
33183 => "1000011001111100",
33184 => "1000011010000000",
33185 => "1000011010000100",
33186 => "1000011010001000",
33187 => "1000011010001100",
33188 => "1000011010010000",
33189 => "1000011010010100",
33190 => "1000011010011000",
33191 => "1000011010011100",
33192 => "1000011010100000",
33193 => "1000011010100100",
33194 => "1000011010101000",
33195 => "1000011010101100",
33196 => "1000011010110000",
33197 => "1000011010110100",
33198 => "1000011010111000",
33199 => "1000011010111100",
33200 => "1000011011000000",
33201 => "1000011011000100",
33202 => "1000011011001000",
33203 => "1000011011001100",
33204 => "1000011011010000",
33205 => "1000011011010100",
33206 => "1000011011011000",
33207 => "1000011011011100",
33208 => "1000011011100000",
33209 => "1000011011100100",
33210 => "1000011011101000",
33211 => "1000011011101100",
33212 => "1000011011110000",
33213 => "1000011011110100",
33214 => "1000011011111000",
33215 => "1000011011111100",
33216 => "1000011100000000",
33217 => "1000011100000100",
33218 => "1000011100001000",
33219 => "1000011100001100",
33220 => "1000011100010000",
33221 => "1000011100010100",
33222 => "1000011100011000",
33223 => "1000011100011100",
33224 => "1000011100100000",
33225 => "1000011100100100",
33226 => "1000011100101000",
33227 => "1000011100101100",
33228 => "1000011100110000",
33229 => "1000011100110100",
33230 => "1000011100111000",
33231 => "1000011100111100",
33232 => "1000011101000000",
33233 => "1000011101000100",
33234 => "1000011101001000",
33235 => "1000011101001100",
33236 => "1000011101001111",
33237 => "1000011101010011",
33238 => "1000011101010111",
33239 => "1000011101011011",
33240 => "1000011101011111",
33241 => "1000011101100011",
33242 => "1000011101100111",
33243 => "1000011101101011",
33244 => "1000011101101111",
33245 => "1000011101110011",
33246 => "1000011101110111",
33247 => "1000011101111011",
33248 => "1000011101111111",
33249 => "1000011110000011",
33250 => "1000011110000111",
33251 => "1000011110001011",
33252 => "1000011110001111",
33253 => "1000011110010011",
33254 => "1000011110010111",
33255 => "1000011110011011",
33256 => "1000011110011111",
33257 => "1000011110100011",
33258 => "1000011110100111",
33259 => "1000011110101011",
33260 => "1000011110101111",
33261 => "1000011110110011",
33262 => "1000011110110111",
33263 => "1000011110111011",
33264 => "1000011110111111",
33265 => "1000011111000011",
33266 => "1000011111000111",
33267 => "1000011111001011",
33268 => "1000011111001111",
33269 => "1000011111010011",
33270 => "1000011111010111",
33271 => "1000011111011011",
33272 => "1000011111011111",
33273 => "1000011111100011",
33274 => "1000011111100111",
33275 => "1000011111101011",
33276 => "1000011111101111",
33277 => "1000011111110011",
33278 => "1000011111110111",
33279 => "1000011111111011",
33280 => "1000011111111111",
33281 => "1000100000000011",
33282 => "1000100000000111",
33283 => "1000100000001011",
33284 => "1000100000001111",
33285 => "1000100000010011",
33286 => "1000100000010111",
33287 => "1000100000011011",
33288 => "1000100000011111",
33289 => "1000100000100011",
33290 => "1000100000100111",
33291 => "1000100000101011",
33292 => "1000100000101111",
33293 => "1000100000110011",
33294 => "1000100000110111",
33295 => "1000100000111011",
33296 => "1000100000111111",
33297 => "1000100001000011",
33298 => "1000100001000111",
33299 => "1000100001001011",
33300 => "1000100001001111",
33301 => "1000100001010011",
33302 => "1000100001010111",
33303 => "1000100001011010",
33304 => "1000100001011110",
33305 => "1000100001100010",
33306 => "1000100001100110",
33307 => "1000100001101010",
33308 => "1000100001101110",
33309 => "1000100001110010",
33310 => "1000100001110110",
33311 => "1000100001111010",
33312 => "1000100001111110",
33313 => "1000100010000010",
33314 => "1000100010000110",
33315 => "1000100010001010",
33316 => "1000100010001110",
33317 => "1000100010010010",
33318 => "1000100010010110",
33319 => "1000100010011010",
33320 => "1000100010011110",
33321 => "1000100010100010",
33322 => "1000100010100110",
33323 => "1000100010101010",
33324 => "1000100010101110",
33325 => "1000100010110010",
33326 => "1000100010110110",
33327 => "1000100010111010",
33328 => "1000100010111110",
33329 => "1000100011000010",
33330 => "1000100011000110",
33331 => "1000100011001010",
33332 => "1000100011001110",
33333 => "1000100011010010",
33334 => "1000100011010110",
33335 => "1000100011011010",
33336 => "1000100011011110",
33337 => "1000100011100010",
33338 => "1000100011100110",
33339 => "1000100011101010",
33340 => "1000100011101110",
33341 => "1000100011110010",
33342 => "1000100011110110",
33343 => "1000100011111010",
33344 => "1000100011111110",
33345 => "1000100100000010",
33346 => "1000100100000110",
33347 => "1000100100001010",
33348 => "1000100100001110",
33349 => "1000100100010010",
33350 => "1000100100010110",
33351 => "1000100100011010",
33352 => "1000100100011110",
33353 => "1000100100100010",
33354 => "1000100100100110",
33355 => "1000100100101010",
33356 => "1000100100101101",
33357 => "1000100100110001",
33358 => "1000100100110101",
33359 => "1000100100111001",
33360 => "1000100100111101",
33361 => "1000100101000001",
33362 => "1000100101000101",
33363 => "1000100101001001",
33364 => "1000100101001101",
33365 => "1000100101010001",
33366 => "1000100101010101",
33367 => "1000100101011001",
33368 => "1000100101011101",
33369 => "1000100101100001",
33370 => "1000100101100101",
33371 => "1000100101101001",
33372 => "1000100101101101",
33373 => "1000100101110001",
33374 => "1000100101110101",
33375 => "1000100101111001",
33376 => "1000100101111101",
33377 => "1000100110000001",
33378 => "1000100110000101",
33379 => "1000100110001001",
33380 => "1000100110001101",
33381 => "1000100110010001",
33382 => "1000100110010101",
33383 => "1000100110011001",
33384 => "1000100110011101",
33385 => "1000100110100001",
33386 => "1000100110100101",
33387 => "1000100110101001",
33388 => "1000100110101101",
33389 => "1000100110110001",
33390 => "1000100110110101",
33391 => "1000100110111001",
33392 => "1000100110111101",
33393 => "1000100111000001",
33394 => "1000100111000101",
33395 => "1000100111001001",
33396 => "1000100111001101",
33397 => "1000100111010001",
33398 => "1000100111010101",
33399 => "1000100111011001",
33400 => "1000100111011101",
33401 => "1000100111100000",
33402 => "1000100111100100",
33403 => "1000100111101000",
33404 => "1000100111101100",
33405 => "1000100111110000",
33406 => "1000100111110100",
33407 => "1000100111111000",
33408 => "1000100111111100",
33409 => "1000101000000000",
33410 => "1000101000000100",
33411 => "1000101000001000",
33412 => "1000101000001100",
33413 => "1000101000010000",
33414 => "1000101000010100",
33415 => "1000101000011000",
33416 => "1000101000011100",
33417 => "1000101000100000",
33418 => "1000101000100100",
33419 => "1000101000101000",
33420 => "1000101000101100",
33421 => "1000101000110000",
33422 => "1000101000110100",
33423 => "1000101000111000",
33424 => "1000101000111100",
33425 => "1000101001000000",
33426 => "1000101001000100",
33427 => "1000101001001000",
33428 => "1000101001001100",
33429 => "1000101001010000",
33430 => "1000101001010100",
33431 => "1000101001011000",
33432 => "1000101001011100",
33433 => "1000101001100000",
33434 => "1000101001100100",
33435 => "1000101001101000",
33436 => "1000101001101100",
33437 => "1000101001110000",
33438 => "1000101001110100",
33439 => "1000101001111000",
33440 => "1000101001111100",
33441 => "1000101001111111",
33442 => "1000101010000011",
33443 => "1000101010000111",
33444 => "1000101010001011",
33445 => "1000101010001111",
33446 => "1000101010010011",
33447 => "1000101010010111",
33448 => "1000101010011011",
33449 => "1000101010011111",
33450 => "1000101010100011",
33451 => "1000101010100111",
33452 => "1000101010101011",
33453 => "1000101010101111",
33454 => "1000101010110011",
33455 => "1000101010110111",
33456 => "1000101010111011",
33457 => "1000101010111111",
33458 => "1000101011000011",
33459 => "1000101011000111",
33460 => "1000101011001011",
33461 => "1000101011001111",
33462 => "1000101011010011",
33463 => "1000101011010111",
33464 => "1000101011011011",
33465 => "1000101011011111",
33466 => "1000101011100011",
33467 => "1000101011100111",
33468 => "1000101011101011",
33469 => "1000101011101111",
33470 => "1000101011110011",
33471 => "1000101011110111",
33472 => "1000101011111011",
33473 => "1000101011111111",
33474 => "1000101100000011",
33475 => "1000101100000111",
33476 => "1000101100001010",
33477 => "1000101100001110",
33478 => "1000101100010010",
33479 => "1000101100010110",
33480 => "1000101100011010",
33481 => "1000101100011110",
33482 => "1000101100100010",
33483 => "1000101100100110",
33484 => "1000101100101010",
33485 => "1000101100101110",
33486 => "1000101100110010",
33487 => "1000101100110110",
33488 => "1000101100111010",
33489 => "1000101100111110",
33490 => "1000101101000010",
33491 => "1000101101000110",
33492 => "1000101101001010",
33493 => "1000101101001110",
33494 => "1000101101010010",
33495 => "1000101101010110",
33496 => "1000101101011010",
33497 => "1000101101011110",
33498 => "1000101101100010",
33499 => "1000101101100110",
33500 => "1000101101101010",
33501 => "1000101101101110",
33502 => "1000101101110010",
33503 => "1000101101110110",
33504 => "1000101101111010",
33505 => "1000101101111110",
33506 => "1000101110000010",
33507 => "1000101110000110",
33508 => "1000101110001010",
33509 => "1000101110001101",
33510 => "1000101110010001",
33511 => "1000101110010101",
33512 => "1000101110011001",
33513 => "1000101110011101",
33514 => "1000101110100001",
33515 => "1000101110100101",
33516 => "1000101110101001",
33517 => "1000101110101101",
33518 => "1000101110110001",
33519 => "1000101110110101",
33520 => "1000101110111001",
33521 => "1000101110111101",
33522 => "1000101111000001",
33523 => "1000101111000101",
33524 => "1000101111001001",
33525 => "1000101111001101",
33526 => "1000101111010001",
33527 => "1000101111010101",
33528 => "1000101111011001",
33529 => "1000101111011101",
33530 => "1000101111100001",
33531 => "1000101111100101",
33532 => "1000101111101001",
33533 => "1000101111101101",
33534 => "1000101111110001",
33535 => "1000101111110101",
33536 => "1000101111111001",
33537 => "1000101111111101",
33538 => "1000110000000000",
33539 => "1000110000000100",
33540 => "1000110000001000",
33541 => "1000110000001100",
33542 => "1000110000010000",
33543 => "1000110000010100",
33544 => "1000110000011000",
33545 => "1000110000011100",
33546 => "1000110000100000",
33547 => "1000110000100100",
33548 => "1000110000101000",
33549 => "1000110000101100",
33550 => "1000110000110000",
33551 => "1000110000110100",
33552 => "1000110000111000",
33553 => "1000110000111100",
33554 => "1000110001000000",
33555 => "1000110001000100",
33556 => "1000110001001000",
33557 => "1000110001001100",
33558 => "1000110001010000",
33559 => "1000110001010100",
33560 => "1000110001011000",
33561 => "1000110001011100",
33562 => "1000110001100000",
33563 => "1000110001100100",
33564 => "1000110001101000",
33565 => "1000110001101100",
33566 => "1000110001101111",
33567 => "1000110001110011",
33568 => "1000110001110111",
33569 => "1000110001111011",
33570 => "1000110001111111",
33571 => "1000110010000011",
33572 => "1000110010000111",
33573 => "1000110010001011",
33574 => "1000110010001111",
33575 => "1000110010010011",
33576 => "1000110010010111",
33577 => "1000110010011011",
33578 => "1000110010011111",
33579 => "1000110010100011",
33580 => "1000110010100111",
33581 => "1000110010101011",
33582 => "1000110010101111",
33583 => "1000110010110011",
33584 => "1000110010110111",
33585 => "1000110010111011",
33586 => "1000110010111111",
33587 => "1000110011000011",
33588 => "1000110011000111",
33589 => "1000110011001011",
33590 => "1000110011001111",
33591 => "1000110011010010",
33592 => "1000110011010110",
33593 => "1000110011011010",
33594 => "1000110011011110",
33595 => "1000110011100010",
33596 => "1000110011100110",
33597 => "1000110011101010",
33598 => "1000110011101110",
33599 => "1000110011110010",
33600 => "1000110011110110",
33601 => "1000110011111010",
33602 => "1000110011111110",
33603 => "1000110100000010",
33604 => "1000110100000110",
33605 => "1000110100001010",
33606 => "1000110100001110",
33607 => "1000110100010010",
33608 => "1000110100010110",
33609 => "1000110100011010",
33610 => "1000110100011110",
33611 => "1000110100100010",
33612 => "1000110100100110",
33613 => "1000110100101010",
33614 => "1000110100101110",
33615 => "1000110100110010",
33616 => "1000110100110101",
33617 => "1000110100111001",
33618 => "1000110100111101",
33619 => "1000110101000001",
33620 => "1000110101000101",
33621 => "1000110101001001",
33622 => "1000110101001101",
33623 => "1000110101010001",
33624 => "1000110101010101",
33625 => "1000110101011001",
33626 => "1000110101011101",
33627 => "1000110101100001",
33628 => "1000110101100101",
33629 => "1000110101101001",
33630 => "1000110101101101",
33631 => "1000110101110001",
33632 => "1000110101110101",
33633 => "1000110101111001",
33634 => "1000110101111101",
33635 => "1000110110000001",
33636 => "1000110110000101",
33637 => "1000110110001001",
33638 => "1000110110001101",
33639 => "1000110110010000",
33640 => "1000110110010100",
33641 => "1000110110011000",
33642 => "1000110110011100",
33643 => "1000110110100000",
33644 => "1000110110100100",
33645 => "1000110110101000",
33646 => "1000110110101100",
33647 => "1000110110110000",
33648 => "1000110110110100",
33649 => "1000110110111000",
33650 => "1000110110111100",
33651 => "1000110111000000",
33652 => "1000110111000100",
33653 => "1000110111001000",
33654 => "1000110111001100",
33655 => "1000110111010000",
33656 => "1000110111010100",
33657 => "1000110111011000",
33658 => "1000110111011100",
33659 => "1000110111100000",
33660 => "1000110111100011",
33661 => "1000110111100111",
33662 => "1000110111101011",
33663 => "1000110111101111",
33664 => "1000110111110011",
33665 => "1000110111110111",
33666 => "1000110111111011",
33667 => "1000110111111111",
33668 => "1000111000000011",
33669 => "1000111000000111",
33670 => "1000111000001011",
33671 => "1000111000001111",
33672 => "1000111000010011",
33673 => "1000111000010111",
33674 => "1000111000011011",
33675 => "1000111000011111",
33676 => "1000111000100011",
33677 => "1000111000100111",
33678 => "1000111000101011",
33679 => "1000111000101111",
33680 => "1000111000110011",
33681 => "1000111000110110",
33682 => "1000111000111010",
33683 => "1000111000111110",
33684 => "1000111001000010",
33685 => "1000111001000110",
33686 => "1000111001001010",
33687 => "1000111001001110",
33688 => "1000111001010010",
33689 => "1000111001010110",
33690 => "1000111001011010",
33691 => "1000111001011110",
33692 => "1000111001100010",
33693 => "1000111001100110",
33694 => "1000111001101010",
33695 => "1000111001101110",
33696 => "1000111001110010",
33697 => "1000111001110110",
33698 => "1000111001111010",
33699 => "1000111001111110",
33700 => "1000111010000010",
33701 => "1000111010000101",
33702 => "1000111010001001",
33703 => "1000111010001101",
33704 => "1000111010010001",
33705 => "1000111010010101",
33706 => "1000111010011001",
33707 => "1000111010011101",
33708 => "1000111010100001",
33709 => "1000111010100101",
33710 => "1000111010101001",
33711 => "1000111010101101",
33712 => "1000111010110001",
33713 => "1000111010110101",
33714 => "1000111010111001",
33715 => "1000111010111101",
33716 => "1000111011000001",
33717 => "1000111011000101",
33718 => "1000111011001001",
33719 => "1000111011001101",
33720 => "1000111011010000",
33721 => "1000111011010100",
33722 => "1000111011011000",
33723 => "1000111011011100",
33724 => "1000111011100000",
33725 => "1000111011100100",
33726 => "1000111011101000",
33727 => "1000111011101100",
33728 => "1000111011110000",
33729 => "1000111011110100",
33730 => "1000111011111000",
33731 => "1000111011111100",
33732 => "1000111100000000",
33733 => "1000111100000100",
33734 => "1000111100001000",
33735 => "1000111100001100",
33736 => "1000111100010000",
33737 => "1000111100010100",
33738 => "1000111100010111",
33739 => "1000111100011011",
33740 => "1000111100011111",
33741 => "1000111100100011",
33742 => "1000111100100111",
33743 => "1000111100101011",
33744 => "1000111100101111",
33745 => "1000111100110011",
33746 => "1000111100110111",
33747 => "1000111100111011",
33748 => "1000111100111111",
33749 => "1000111101000011",
33750 => "1000111101000111",
33751 => "1000111101001011",
33752 => "1000111101001111",
33753 => "1000111101010011",
33754 => "1000111101010111",
33755 => "1000111101011011",
33756 => "1000111101011110",
33757 => "1000111101100010",
33758 => "1000111101100110",
33759 => "1000111101101010",
33760 => "1000111101101110",
33761 => "1000111101110010",
33762 => "1000111101110110",
33763 => "1000111101111010",
33764 => "1000111101111110",
33765 => "1000111110000010",
33766 => "1000111110000110",
33767 => "1000111110001010",
33768 => "1000111110001110",
33769 => "1000111110010010",
33770 => "1000111110010110",
33771 => "1000111110011010",
33772 => "1000111110011110",
33773 => "1000111110100001",
33774 => "1000111110100101",
33775 => "1000111110101001",
33776 => "1000111110101101",
33777 => "1000111110110001",
33778 => "1000111110110101",
33779 => "1000111110111001",
33780 => "1000111110111101",
33781 => "1000111111000001",
33782 => "1000111111000101",
33783 => "1000111111001001",
33784 => "1000111111001101",
33785 => "1000111111010001",
33786 => "1000111111010101",
33787 => "1000111111011001",
33788 => "1000111111011101",
33789 => "1000111111100001",
33790 => "1000111111100100",
33791 => "1000111111101000",
33792 => "1000111111101100",
33793 => "1000111111110000",
33794 => "1000111111110100",
33795 => "1000111111111000",
33796 => "1000111111111100",
33797 => "1001000000000000",
33798 => "1001000000000100",
33799 => "1001000000001000",
33800 => "1001000000001100",
33801 => "1001000000010000",
33802 => "1001000000010100",
33803 => "1001000000011000",
33804 => "1001000000011100",
33805 => "1001000000100000",
33806 => "1001000000100011",
33807 => "1001000000100111",
33808 => "1001000000101011",
33809 => "1001000000101111",
33810 => "1001000000110011",
33811 => "1001000000110111",
33812 => "1001000000111011",
33813 => "1001000000111111",
33814 => "1001000001000011",
33815 => "1001000001000111",
33816 => "1001000001001011",
33817 => "1001000001001111",
33818 => "1001000001010011",
33819 => "1001000001010111",
33820 => "1001000001011011",
33821 => "1001000001011110",
33822 => "1001000001100010",
33823 => "1001000001100110",
33824 => "1001000001101010",
33825 => "1001000001101110",
33826 => "1001000001110010",
33827 => "1001000001110110",
33828 => "1001000001111010",
33829 => "1001000001111110",
33830 => "1001000010000010",
33831 => "1001000010000110",
33832 => "1001000010001010",
33833 => "1001000010001110",
33834 => "1001000010010010",
33835 => "1001000010010110",
33836 => "1001000010011001",
33837 => "1001000010011101",
33838 => "1001000010100001",
33839 => "1001000010100101",
33840 => "1001000010101001",
33841 => "1001000010101101",
33842 => "1001000010110001",
33843 => "1001000010110101",
33844 => "1001000010111001",
33845 => "1001000010111101",
33846 => "1001000011000001",
33847 => "1001000011000101",
33848 => "1001000011001001",
33849 => "1001000011001101",
33850 => "1001000011010001",
33851 => "1001000011010100",
33852 => "1001000011011000",
33853 => "1001000011011100",
33854 => "1001000011100000",
33855 => "1001000011100100",
33856 => "1001000011101000",
33857 => "1001000011101100",
33858 => "1001000011110000",
33859 => "1001000011110100",
33860 => "1001000011111000",
33861 => "1001000011111100",
33862 => "1001000100000000",
33863 => "1001000100000100",
33864 => "1001000100001000",
33865 => "1001000100001011",
33866 => "1001000100001111",
33867 => "1001000100010011",
33868 => "1001000100010111",
33869 => "1001000100011011",
33870 => "1001000100011111",
33871 => "1001000100100011",
33872 => "1001000100100111",
33873 => "1001000100101011",
33874 => "1001000100101111",
33875 => "1001000100110011",
33876 => "1001000100110111",
33877 => "1001000100111011",
33878 => "1001000100111111",
33879 => "1001000101000010",
33880 => "1001000101000110",
33881 => "1001000101001010",
33882 => "1001000101001110",
33883 => "1001000101010010",
33884 => "1001000101010110",
33885 => "1001000101011010",
33886 => "1001000101011110",
33887 => "1001000101100010",
33888 => "1001000101100110",
33889 => "1001000101101010",
33890 => "1001000101101110",
33891 => "1001000101110010",
33892 => "1001000101110110",
33893 => "1001000101111001",
33894 => "1001000101111101",
33895 => "1001000110000001",
33896 => "1001000110000101",
33897 => "1001000110001001",
33898 => "1001000110001101",
33899 => "1001000110010001",
33900 => "1001000110010101",
33901 => "1001000110011001",
33902 => "1001000110011101",
33903 => "1001000110100001",
33904 => "1001000110100101",
33905 => "1001000110101001",
33906 => "1001000110101100",
33907 => "1001000110110000",
33908 => "1001000110110100",
33909 => "1001000110111000",
33910 => "1001000110111100",
33911 => "1001000111000000",
33912 => "1001000111000100",
33913 => "1001000111001000",
33914 => "1001000111001100",
33915 => "1001000111010000",
33916 => "1001000111010100",
33917 => "1001000111011000",
33918 => "1001000111011100",
33919 => "1001000111011111",
33920 => "1001000111100011",
33921 => "1001000111100111",
33922 => "1001000111101011",
33923 => "1001000111101111",
33924 => "1001000111110011",
33925 => "1001000111110111",
33926 => "1001000111111011",
33927 => "1001000111111111",
33928 => "1001001000000011",
33929 => "1001001000000111",
33930 => "1001001000001011",
33931 => "1001001000001111",
33932 => "1001001000010010",
33933 => "1001001000010110",
33934 => "1001001000011010",
33935 => "1001001000011110",
33936 => "1001001000100010",
33937 => "1001001000100110",
33938 => "1001001000101010",
33939 => "1001001000101110",
33940 => "1001001000110010",
33941 => "1001001000110110",
33942 => "1001001000111010",
33943 => "1001001000111110",
33944 => "1001001001000001",
33945 => "1001001001000101",
33946 => "1001001001001001",
33947 => "1001001001001101",
33948 => "1001001001010001",
33949 => "1001001001010101",
33950 => "1001001001011001",
33951 => "1001001001011101",
33952 => "1001001001100001",
33953 => "1001001001100101",
33954 => "1001001001101001",
33955 => "1001001001101101",
33956 => "1001001001110000",
33957 => "1001001001110100",
33958 => "1001001001111000",
33959 => "1001001001111100",
33960 => "1001001010000000",
33961 => "1001001010000100",
33962 => "1001001010001000",
33963 => "1001001010001100",
33964 => "1001001010010000",
33965 => "1001001010010100",
33966 => "1001001010011000",
33967 => "1001001010011100",
33968 => "1001001010011111",
33969 => "1001001010100011",
33970 => "1001001010100111",
33971 => "1001001010101011",
33972 => "1001001010101111",
33973 => "1001001010110011",
33974 => "1001001010110111",
33975 => "1001001010111011",
33976 => "1001001010111111",
33977 => "1001001011000011",
33978 => "1001001011000111",
33979 => "1001001011001011",
33980 => "1001001011001110",
33981 => "1001001011010010",
33982 => "1001001011010110",
33983 => "1001001011011010",
33984 => "1001001011011110",
33985 => "1001001011100010",
33986 => "1001001011100110",
33987 => "1001001011101010",
33988 => "1001001011101110",
33989 => "1001001011110010",
33990 => "1001001011110110",
33991 => "1001001011111010",
33992 => "1001001011111101",
33993 => "1001001100000001",
33994 => "1001001100000101",
33995 => "1001001100001001",
33996 => "1001001100001101",
33997 => "1001001100010001",
33998 => "1001001100010101",
33999 => "1001001100011001",
34000 => "1001001100011101",
34001 => "1001001100100001",
34002 => "1001001100100101",
34003 => "1001001100101000",
34004 => "1001001100101100",
34005 => "1001001100110000",
34006 => "1001001100110100",
34007 => "1001001100111000",
34008 => "1001001100111100",
34009 => "1001001101000000",
34010 => "1001001101000100",
34011 => "1001001101001000",
34012 => "1001001101001100",
34013 => "1001001101010000",
34014 => "1001001101010011",
34015 => "1001001101010111",
34016 => "1001001101011011",
34017 => "1001001101011111",
34018 => "1001001101100011",
34019 => "1001001101100111",
34020 => "1001001101101011",
34021 => "1001001101101111",
34022 => "1001001101110011",
34023 => "1001001101110111",
34024 => "1001001101111011",
34025 => "1001001101111110",
34026 => "1001001110000010",
34027 => "1001001110000110",
34028 => "1001001110001010",
34029 => "1001001110001110",
34030 => "1001001110010010",
34031 => "1001001110010110",
34032 => "1001001110011010",
34033 => "1001001110011110",
34034 => "1001001110100010",
34035 => "1001001110100110",
34036 => "1001001110101001",
34037 => "1001001110101101",
34038 => "1001001110110001",
34039 => "1001001110110101",
34040 => "1001001110111001",
34041 => "1001001110111101",
34042 => "1001001111000001",
34043 => "1001001111000101",
34044 => "1001001111001001",
34045 => "1001001111001101",
34046 => "1001001111010000",
34047 => "1001001111010100",
34048 => "1001001111011000",
34049 => "1001001111011100",
34050 => "1001001111100000",
34051 => "1001001111100100",
34052 => "1001001111101000",
34053 => "1001001111101100",
34054 => "1001001111110000",
34055 => "1001001111110100",
34056 => "1001001111110111",
34057 => "1001001111111011",
34058 => "1001001111111111",
34059 => "1001010000000011",
34060 => "1001010000000111",
34061 => "1001010000001011",
34062 => "1001010000001111",
34063 => "1001010000010011",
34064 => "1001010000010111",
34065 => "1001010000011011",
34066 => "1001010000011111",
34067 => "1001010000100010",
34068 => "1001010000100110",
34069 => "1001010000101010",
34070 => "1001010000101110",
34071 => "1001010000110010",
34072 => "1001010000110110",
34073 => "1001010000111010",
34074 => "1001010000111110",
34075 => "1001010001000010",
34076 => "1001010001000110",
34077 => "1001010001001001",
34078 => "1001010001001101",
34079 => "1001010001010001",
34080 => "1001010001010101",
34081 => "1001010001011001",
34082 => "1001010001011101",
34083 => "1001010001100001",
34084 => "1001010001100101",
34085 => "1001010001101001",
34086 => "1001010001101101",
34087 => "1001010001110000",
34088 => "1001010001110100",
34089 => "1001010001111000",
34090 => "1001010001111100",
34091 => "1001010010000000",
34092 => "1001010010000100",
34093 => "1001010010001000",
34094 => "1001010010001100",
34095 => "1001010010010000",
34096 => "1001010010010011",
34097 => "1001010010010111",
34098 => "1001010010011011",
34099 => "1001010010011111",
34100 => "1001010010100011",
34101 => "1001010010100111",
34102 => "1001010010101011",
34103 => "1001010010101111",
34104 => "1001010010110011",
34105 => "1001010010110111",
34106 => "1001010010111010",
34107 => "1001010010111110",
34108 => "1001010011000010",
34109 => "1001010011000110",
34110 => "1001010011001010",
34111 => "1001010011001110",
34112 => "1001010011010010",
34113 => "1001010011010110",
34114 => "1001010011011010",
34115 => "1001010011011101",
34116 => "1001010011100001",
34117 => "1001010011100101",
34118 => "1001010011101001",
34119 => "1001010011101101",
34120 => "1001010011110001",
34121 => "1001010011110101",
34122 => "1001010011111001",
34123 => "1001010011111101",
34124 => "1001010100000001",
34125 => "1001010100000100",
34126 => "1001010100001000",
34127 => "1001010100001100",
34128 => "1001010100010000",
34129 => "1001010100010100",
34130 => "1001010100011000",
34131 => "1001010100011100",
34132 => "1001010100100000",
34133 => "1001010100100100",
34134 => "1001010100100111",
34135 => "1001010100101011",
34136 => "1001010100101111",
34137 => "1001010100110011",
34138 => "1001010100110111",
34139 => "1001010100111011",
34140 => "1001010100111111",
34141 => "1001010101000011",
34142 => "1001010101000111",
34143 => "1001010101001010",
34144 => "1001010101001110",
34145 => "1001010101010010",
34146 => "1001010101010110",
34147 => "1001010101011010",
34148 => "1001010101011110",
34149 => "1001010101100010",
34150 => "1001010101100110",
34151 => "1001010101101010",
34152 => "1001010101101101",
34153 => "1001010101110001",
34154 => "1001010101110101",
34155 => "1001010101111001",
34156 => "1001010101111101",
34157 => "1001010110000001",
34158 => "1001010110000101",
34159 => "1001010110001001",
34160 => "1001010110001101",
34161 => "1001010110010000",
34162 => "1001010110010100",
34163 => "1001010110011000",
34164 => "1001010110011100",
34165 => "1001010110100000",
34166 => "1001010110100100",
34167 => "1001010110101000",
34168 => "1001010110101100",
34169 => "1001010110110000",
34170 => "1001010110110011",
34171 => "1001010110110111",
34172 => "1001010110111011",
34173 => "1001010110111111",
34174 => "1001010111000011",
34175 => "1001010111000111",
34176 => "1001010111001011",
34177 => "1001010111001111",
34178 => "1001010111010010",
34179 => "1001010111010110",
34180 => "1001010111011010",
34181 => "1001010111011110",
34182 => "1001010111100010",
34183 => "1001010111100110",
34184 => "1001010111101010",
34185 => "1001010111101110",
34186 => "1001010111110010",
34187 => "1001010111110101",
34188 => "1001010111111001",
34189 => "1001010111111101",
34190 => "1001011000000001",
34191 => "1001011000000101",
34192 => "1001011000001001",
34193 => "1001011000001101",
34194 => "1001011000010001",
34195 => "1001011000010100",
34196 => "1001011000011000",
34197 => "1001011000011100",
34198 => "1001011000100000",
34199 => "1001011000100100",
34200 => "1001011000101000",
34201 => "1001011000101100",
34202 => "1001011000110000",
34203 => "1001011000110100",
34204 => "1001011000110111",
34205 => "1001011000111011",
34206 => "1001011000111111",
34207 => "1001011001000011",
34208 => "1001011001000111",
34209 => "1001011001001011",
34210 => "1001011001001111",
34211 => "1001011001010011",
34212 => "1001011001010110",
34213 => "1001011001011010",
34214 => "1001011001011110",
34215 => "1001011001100010",
34216 => "1001011001100110",
34217 => "1001011001101010",
34218 => "1001011001101110",
34219 => "1001011001110010",
34220 => "1001011001110101",
34221 => "1001011001111001",
34222 => "1001011001111101",
34223 => "1001011010000001",
34224 => "1001011010000101",
34225 => "1001011010001001",
34226 => "1001011010001101",
34227 => "1001011010010001",
34228 => "1001011010010100",
34229 => "1001011010011000",
34230 => "1001011010011100",
34231 => "1001011010100000",
34232 => "1001011010100100",
34233 => "1001011010101000",
34234 => "1001011010101100",
34235 => "1001011010110000",
34236 => "1001011010110011",
34237 => "1001011010110111",
34238 => "1001011010111011",
34239 => "1001011010111111",
34240 => "1001011011000011",
34241 => "1001011011000111",
34242 => "1001011011001011",
34243 => "1001011011001111",
34244 => "1001011011010010",
34245 => "1001011011010110",
34246 => "1001011011011010",
34247 => "1001011011011110",
34248 => "1001011011100010",
34249 => "1001011011100110",
34250 => "1001011011101010",
34251 => "1001011011101110",
34252 => "1001011011110001",
34253 => "1001011011110101",
34254 => "1001011011111001",
34255 => "1001011011111101",
34256 => "1001011100000001",
34257 => "1001011100000101",
34258 => "1001011100001001",
34259 => "1001011100001101",
34260 => "1001011100010000",
34261 => "1001011100010100",
34262 => "1001011100011000",
34263 => "1001011100011100",
34264 => "1001011100100000",
34265 => "1001011100100100",
34266 => "1001011100101000",
34267 => "1001011100101011",
34268 => "1001011100101111",
34269 => "1001011100110011",
34270 => "1001011100110111",
34271 => "1001011100111011",
34272 => "1001011100111111",
34273 => "1001011101000011",
34274 => "1001011101000111",
34275 => "1001011101001010",
34276 => "1001011101001110",
34277 => "1001011101010010",
34278 => "1001011101010110",
34279 => "1001011101011010",
34280 => "1001011101011110",
34281 => "1001011101100010",
34282 => "1001011101100110",
34283 => "1001011101101001",
34284 => "1001011101101101",
34285 => "1001011101110001",
34286 => "1001011101110101",
34287 => "1001011101111001",
34288 => "1001011101111101",
34289 => "1001011110000001",
34290 => "1001011110000100",
34291 => "1001011110001000",
34292 => "1001011110001100",
34293 => "1001011110010000",
34294 => "1001011110010100",
34295 => "1001011110011000",
34296 => "1001011110011100",
34297 => "1001011110011111",
34298 => "1001011110100011",
34299 => "1001011110100111",
34300 => "1001011110101011",
34301 => "1001011110101111",
34302 => "1001011110110011",
34303 => "1001011110110111",
34304 => "1001011110111011",
34305 => "1001011110111110",
34306 => "1001011111000010",
34307 => "1001011111000110",
34308 => "1001011111001010",
34309 => "1001011111001110",
34310 => "1001011111010010",
34311 => "1001011111010110",
34312 => "1001011111011001",
34313 => "1001011111011101",
34314 => "1001011111100001",
34315 => "1001011111100101",
34316 => "1001011111101001",
34317 => "1001011111101101",
34318 => "1001011111110001",
34319 => "1001011111110100",
34320 => "1001011111111000",
34321 => "1001011111111100",
34322 => "1001100000000000",
34323 => "1001100000000100",
34324 => "1001100000001000",
34325 => "1001100000001100",
34326 => "1001100000001111",
34327 => "1001100000010011",
34328 => "1001100000010111",
34329 => "1001100000011011",
34330 => "1001100000011111",
34331 => "1001100000100011",
34332 => "1001100000100111",
34333 => "1001100000101010",
34334 => "1001100000101110",
34335 => "1001100000110010",
34336 => "1001100000110110",
34337 => "1001100000111010",
34338 => "1001100000111110",
34339 => "1001100001000010",
34340 => "1001100001000101",
34341 => "1001100001001001",
34342 => "1001100001001101",
34343 => "1001100001010001",
34344 => "1001100001010101",
34345 => "1001100001011001",
34346 => "1001100001011101",
34347 => "1001100001100000",
34348 => "1001100001100100",
34349 => "1001100001101000",
34350 => "1001100001101100",
34351 => "1001100001110000",
34352 => "1001100001110100",
34353 => "1001100001111000",
34354 => "1001100001111011",
34355 => "1001100001111111",
34356 => "1001100010000011",
34357 => "1001100010000111",
34358 => "1001100010001011",
34359 => "1001100010001111",
34360 => "1001100010010011",
34361 => "1001100010010110",
34362 => "1001100010011010",
34363 => "1001100010011110",
34364 => "1001100010100010",
34365 => "1001100010100110",
34366 => "1001100010101010",
34367 => "1001100010101110",
34368 => "1001100010110001",
34369 => "1001100010110101",
34370 => "1001100010111001",
34371 => "1001100010111101",
34372 => "1001100011000001",
34373 => "1001100011000101",
34374 => "1001100011001000",
34375 => "1001100011001100",
34376 => "1001100011010000",
34377 => "1001100011010100",
34378 => "1001100011011000",
34379 => "1001100011011100",
34380 => "1001100011100000",
34381 => "1001100011100011",
34382 => "1001100011100111",
34383 => "1001100011101011",
34384 => "1001100011101111",
34385 => "1001100011110011",
34386 => "1001100011110111",
34387 => "1001100011111011",
34388 => "1001100011111110",
34389 => "1001100100000010",
34390 => "1001100100000110",
34391 => "1001100100001010",
34392 => "1001100100001110",
34393 => "1001100100010010",
34394 => "1001100100010101",
34395 => "1001100100011001",
34396 => "1001100100011101",
34397 => "1001100100100001",
34398 => "1001100100100101",
34399 => "1001100100101001",
34400 => "1001100100101101",
34401 => "1001100100110000",
34402 => "1001100100110100",
34403 => "1001100100111000",
34404 => "1001100100111100",
34405 => "1001100101000000",
34406 => "1001100101000100",
34407 => "1001100101000111",
34408 => "1001100101001011",
34409 => "1001100101001111",
34410 => "1001100101010011",
34411 => "1001100101010111",
34412 => "1001100101011011",
34413 => "1001100101011110",
34414 => "1001100101100010",
34415 => "1001100101100110",
34416 => "1001100101101010",
34417 => "1001100101101110",
34418 => "1001100101110010",
34419 => "1001100101110110",
34420 => "1001100101111001",
34421 => "1001100101111101",
34422 => "1001100110000001",
34423 => "1001100110000101",
34424 => "1001100110001001",
34425 => "1001100110001101",
34426 => "1001100110010000",
34427 => "1001100110010100",
34428 => "1001100110011000",
34429 => "1001100110011100",
34430 => "1001100110100000",
34431 => "1001100110100100",
34432 => "1001100110100111",
34433 => "1001100110101011",
34434 => "1001100110101111",
34435 => "1001100110110011",
34436 => "1001100110110111",
34437 => "1001100110111011",
34438 => "1001100110111110",
34439 => "1001100111000010",
34440 => "1001100111000110",
34441 => "1001100111001010",
34442 => "1001100111001110",
34443 => "1001100111010010",
34444 => "1001100111010110",
34445 => "1001100111011001",
34446 => "1001100111011101",
34447 => "1001100111100001",
34448 => "1001100111100101",
34449 => "1001100111101001",
34450 => "1001100111101101",
34451 => "1001100111110000",
34452 => "1001100111110100",
34453 => "1001100111111000",
34454 => "1001100111111100",
34455 => "1001101000000000",
34456 => "1001101000000100",
34457 => "1001101000000111",
34458 => "1001101000001011",
34459 => "1001101000001111",
34460 => "1001101000010011",
34461 => "1001101000010111",
34462 => "1001101000011011",
34463 => "1001101000011110",
34464 => "1001101000100010",
34465 => "1001101000100110",
34466 => "1001101000101010",
34467 => "1001101000101110",
34468 => "1001101000110010",
34469 => "1001101000110101",
34470 => "1001101000111001",
34471 => "1001101000111101",
34472 => "1001101001000001",
34473 => "1001101001000101",
34474 => "1001101001001001",
34475 => "1001101001001100",
34476 => "1001101001010000",
34477 => "1001101001010100",
34478 => "1001101001011000",
34479 => "1001101001011100",
34480 => "1001101001100000",
34481 => "1001101001100011",
34482 => "1001101001100111",
34483 => "1001101001101011",
34484 => "1001101001101111",
34485 => "1001101001110011",
34486 => "1001101001110111",
34487 => "1001101001111010",
34488 => "1001101001111110",
34489 => "1001101010000010",
34490 => "1001101010000110",
34491 => "1001101010001010",
34492 => "1001101010001101",
34493 => "1001101010010001",
34494 => "1001101010010101",
34495 => "1001101010011001",
34496 => "1001101010011101",
34497 => "1001101010100001",
34498 => "1001101010100100",
34499 => "1001101010101000",
34500 => "1001101010101100",
34501 => "1001101010110000",
34502 => "1001101010110100",
34503 => "1001101010111000",
34504 => "1001101010111011",
34505 => "1001101010111111",
34506 => "1001101011000011",
34507 => "1001101011000111",
34508 => "1001101011001011",
34509 => "1001101011001111",
34510 => "1001101011010010",
34511 => "1001101011010110",
34512 => "1001101011011010",
34513 => "1001101011011110",
34514 => "1001101011100010",
34515 => "1001101011100101",
34516 => "1001101011101001",
34517 => "1001101011101101",
34518 => "1001101011110001",
34519 => "1001101011110101",
34520 => "1001101011111001",
34521 => "1001101011111100",
34522 => "1001101100000000",
34523 => "1001101100000100",
34524 => "1001101100001000",
34525 => "1001101100001100",
34526 => "1001101100010000",
34527 => "1001101100010011",
34528 => "1001101100010111",
34529 => "1001101100011011",
34530 => "1001101100011111",
34531 => "1001101100100011",
34532 => "1001101100100110",
34533 => "1001101100101010",
34534 => "1001101100101110",
34535 => "1001101100110010",
34536 => "1001101100110110",
34537 => "1001101100111010",
34538 => "1001101100111101",
34539 => "1001101101000001",
34540 => "1001101101000101",
34541 => "1001101101001001",
34542 => "1001101101001101",
34543 => "1001101101010000",
34544 => "1001101101010100",
34545 => "1001101101011000",
34546 => "1001101101011100",
34547 => "1001101101100000",
34548 => "1001101101100100",
34549 => "1001101101100111",
34550 => "1001101101101011",
34551 => "1001101101101111",
34552 => "1001101101110011",
34553 => "1001101101110111",
34554 => "1001101101111010",
34555 => "1001101101111110",
34556 => "1001101110000010",
34557 => "1001101110000110",
34558 => "1001101110001010",
34559 => "1001101110001110",
34560 => "1001101110010001",
34561 => "1001101110010101",
34562 => "1001101110011001",
34563 => "1001101110011101",
34564 => "1001101110100001",
34565 => "1001101110100100",
34566 => "1001101110101000",
34567 => "1001101110101100",
34568 => "1001101110110000",
34569 => "1001101110110100",
34570 => "1001101110110111",
34571 => "1001101110111011",
34572 => "1001101110111111",
34573 => "1001101111000011",
34574 => "1001101111000111",
34575 => "1001101111001011",
34576 => "1001101111001110",
34577 => "1001101111010010",
34578 => "1001101111010110",
34579 => "1001101111011010",
34580 => "1001101111011110",
34581 => "1001101111100001",
34582 => "1001101111100101",
34583 => "1001101111101001",
34584 => "1001101111101101",
34585 => "1001101111110001",
34586 => "1001101111110100",
34587 => "1001101111111000",
34588 => "1001101111111100",
34589 => "1001110000000000",
34590 => "1001110000000100",
34591 => "1001110000000111",
34592 => "1001110000001011",
34593 => "1001110000001111",
34594 => "1001110000010011",
34595 => "1001110000010111",
34596 => "1001110000011011",
34597 => "1001110000011110",
34598 => "1001110000100010",
34599 => "1001110000100110",
34600 => "1001110000101010",
34601 => "1001110000101110",
34602 => "1001110000110001",
34603 => "1001110000110101",
34604 => "1001110000111001",
34605 => "1001110000111101",
34606 => "1001110001000001",
34607 => "1001110001000100",
34608 => "1001110001001000",
34609 => "1001110001001100",
34610 => "1001110001010000",
34611 => "1001110001010100",
34612 => "1001110001010111",
34613 => "1001110001011011",
34614 => "1001110001011111",
34615 => "1001110001100011",
34616 => "1001110001100111",
34617 => "1001110001101010",
34618 => "1001110001101110",
34619 => "1001110001110010",
34620 => "1001110001110110",
34621 => "1001110001111010",
34622 => "1001110001111101",
34623 => "1001110010000001",
34624 => "1001110010000101",
34625 => "1001110010001001",
34626 => "1001110010001101",
34627 => "1001110010010000",
34628 => "1001110010010100",
34629 => "1001110010011000",
34630 => "1001110010011100",
34631 => "1001110010100000",
34632 => "1001110010100011",
34633 => "1001110010100111",
34634 => "1001110010101011",
34635 => "1001110010101111",
34636 => "1001110010110011",
34637 => "1001110010110110",
34638 => "1001110010111010",
34639 => "1001110010111110",
34640 => "1001110011000010",
34641 => "1001110011000110",
34642 => "1001110011001001",
34643 => "1001110011001101",
34644 => "1001110011010001",
34645 => "1001110011010101",
34646 => "1001110011011001",
34647 => "1001110011011100",
34648 => "1001110011100000",
34649 => "1001110011100100",
34650 => "1001110011101000",
34651 => "1001110011101100",
34652 => "1001110011101111",
34653 => "1001110011110011",
34654 => "1001110011110111",
34655 => "1001110011111011",
34656 => "1001110011111111",
34657 => "1001110100000010",
34658 => "1001110100000110",
34659 => "1001110100001010",
34660 => "1001110100001110",
34661 => "1001110100010010",
34662 => "1001110100010101",
34663 => "1001110100011001",
34664 => "1001110100011101",
34665 => "1001110100100001",
34666 => "1001110100100101",
34667 => "1001110100101000",
34668 => "1001110100101100",
34669 => "1001110100110000",
34670 => "1001110100110100",
34671 => "1001110100110111",
34672 => "1001110100111011",
34673 => "1001110100111111",
34674 => "1001110101000011",
34675 => "1001110101000111",
34676 => "1001110101001010",
34677 => "1001110101001110",
34678 => "1001110101010010",
34679 => "1001110101010110",
34680 => "1001110101011010",
34681 => "1001110101011101",
34682 => "1001110101100001",
34683 => "1001110101100101",
34684 => "1001110101101001",
34685 => "1001110101101101",
34686 => "1001110101110000",
34687 => "1001110101110100",
34688 => "1001110101111000",
34689 => "1001110101111100",
34690 => "1001110101111111",
34691 => "1001110110000011",
34692 => "1001110110000111",
34693 => "1001110110001011",
34694 => "1001110110001111",
34695 => "1001110110010010",
34696 => "1001110110010110",
34697 => "1001110110011010",
34698 => "1001110110011110",
34699 => "1001110110100010",
34700 => "1001110110100101",
34701 => "1001110110101001",
34702 => "1001110110101101",
34703 => "1001110110110001",
34704 => "1001110110110100",
34705 => "1001110110111000",
34706 => "1001110110111100",
34707 => "1001110111000000",
34708 => "1001110111000100",
34709 => "1001110111000111",
34710 => "1001110111001011",
34711 => "1001110111001111",
34712 => "1001110111010011",
34713 => "1001110111010111",
34714 => "1001110111011010",
34715 => "1001110111011110",
34716 => "1001110111100010",
34717 => "1001110111100110",
34718 => "1001110111101001",
34719 => "1001110111101101",
34720 => "1001110111110001",
34721 => "1001110111110101",
34722 => "1001110111111001",
34723 => "1001110111111100",
34724 => "1001111000000000",
34725 => "1001111000000100",
34726 => "1001111000001000",
34727 => "1001111000001011",
34728 => "1001111000001111",
34729 => "1001111000010011",
34730 => "1001111000010111",
34731 => "1001111000011011",
34732 => "1001111000011110",
34733 => "1001111000100010",
34734 => "1001111000100110",
34735 => "1001111000101010",
34736 => "1001111000101101",
34737 => "1001111000110001",
34738 => "1001111000110101",
34739 => "1001111000111001",
34740 => "1001111000111101",
34741 => "1001111001000000",
34742 => "1001111001000100",
34743 => "1001111001001000",
34744 => "1001111001001100",
34745 => "1001111001001111",
34746 => "1001111001010011",
34747 => "1001111001010111",
34748 => "1001111001011011",
34749 => "1001111001011111",
34750 => "1001111001100010",
34751 => "1001111001100110",
34752 => "1001111001101010",
34753 => "1001111001101110",
34754 => "1001111001110001",
34755 => "1001111001110101",
34756 => "1001111001111001",
34757 => "1001111001111101",
34758 => "1001111010000001",
34759 => "1001111010000100",
34760 => "1001111010001000",
34761 => "1001111010001100",
34762 => "1001111010010000",
34763 => "1001111010010011",
34764 => "1001111010010111",
34765 => "1001111010011011",
34766 => "1001111010011111",
34767 => "1001111010100010",
34768 => "1001111010100110",
34769 => "1001111010101010",
34770 => "1001111010101110",
34771 => "1001111010110010",
34772 => "1001111010110101",
34773 => "1001111010111001",
34774 => "1001111010111101",
34775 => "1001111011000001",
34776 => "1001111011000100",
34777 => "1001111011001000",
34778 => "1001111011001100",
34779 => "1001111011010000",
34780 => "1001111011010011",
34781 => "1001111011010111",
34782 => "1001111011011011",
34783 => "1001111011011111",
34784 => "1001111011100011",
34785 => "1001111011100110",
34786 => "1001111011101010",
34787 => "1001111011101110",
34788 => "1001111011110010",
34789 => "1001111011110101",
34790 => "1001111011111001",
34791 => "1001111011111101",
34792 => "1001111100000001",
34793 => "1001111100000100",
34794 => "1001111100001000",
34795 => "1001111100001100",
34796 => "1001111100010000",
34797 => "1001111100010100",
34798 => "1001111100010111",
34799 => "1001111100011011",
34800 => "1001111100011111",
34801 => "1001111100100011",
34802 => "1001111100100110",
34803 => "1001111100101010",
34804 => "1001111100101110",
34805 => "1001111100110010",
34806 => "1001111100110101",
34807 => "1001111100111001",
34808 => "1001111100111101",
34809 => "1001111101000001",
34810 => "1001111101000100",
34811 => "1001111101001000",
34812 => "1001111101001100",
34813 => "1001111101010000",
34814 => "1001111101010011",
34815 => "1001111101010111",
34816 => "1001111101011011",
34817 => "1001111101011111",
34818 => "1001111101100011",
34819 => "1001111101100110",
34820 => "1001111101101010",
34821 => "1001111101101110",
34822 => "1001111101110010",
34823 => "1001111101110101",
34824 => "1001111101111001",
34825 => "1001111101111101",
34826 => "1001111110000001",
34827 => "1001111110000100",
34828 => "1001111110001000",
34829 => "1001111110001100",
34830 => "1001111110010000",
34831 => "1001111110010011",
34832 => "1001111110010111",
34833 => "1001111110011011",
34834 => "1001111110011111",
34835 => "1001111110100010",
34836 => "1001111110100110",
34837 => "1001111110101010",
34838 => "1001111110101110",
34839 => "1001111110110001",
34840 => "1001111110110101",
34841 => "1001111110111001",
34842 => "1001111110111101",
34843 => "1001111111000000",
34844 => "1001111111000100",
34845 => "1001111111001000",
34846 => "1001111111001100",
34847 => "1001111111001111",
34848 => "1001111111010011",
34849 => "1001111111010111",
34850 => "1001111111011011",
34851 => "1001111111011110",
34852 => "1001111111100010",
34853 => "1001111111100110",
34854 => "1001111111101010",
34855 => "1001111111101101",
34856 => "1001111111110001",
34857 => "1001111111110101",
34858 => "1001111111111001",
34859 => "1001111111111100",
34860 => "1010000000000000",
34861 => "1010000000000100",
34862 => "1010000000001000",
34863 => "1010000000001011",
34864 => "1010000000001111",
34865 => "1010000000010011",
34866 => "1010000000010111",
34867 => "1010000000011010",
34868 => "1010000000011110",
34869 => "1010000000100010",
34870 => "1010000000100110",
34871 => "1010000000101001",
34872 => "1010000000101101",
34873 => "1010000000110001",
34874 => "1010000000110101",
34875 => "1010000000111000",
34876 => "1010000000111100",
34877 => "1010000001000000",
34878 => "1010000001000100",
34879 => "1010000001000111",
34880 => "1010000001001011",
34881 => "1010000001001111",
34882 => "1010000001010011",
34883 => "1010000001010110",
34884 => "1010000001011010",
34885 => "1010000001011110",
34886 => "1010000001100010",
34887 => "1010000001100101",
34888 => "1010000001101001",
34889 => "1010000001101101",
34890 => "1010000001110001",
34891 => "1010000001110100",
34892 => "1010000001111000",
34893 => "1010000001111100",
34894 => "1010000010000000",
34895 => "1010000010000011",
34896 => "1010000010000111",
34897 => "1010000010001011",
34898 => "1010000010001111",
34899 => "1010000010010010",
34900 => "1010000010010110",
34901 => "1010000010011010",
34902 => "1010000010011110",
34903 => "1010000010100001",
34904 => "1010000010100101",
34905 => "1010000010101001",
34906 => "1010000010101100",
34907 => "1010000010110000",
34908 => "1010000010110100",
34909 => "1010000010111000",
34910 => "1010000010111011",
34911 => "1010000010111111",
34912 => "1010000011000011",
34913 => "1010000011000111",
34914 => "1010000011001010",
34915 => "1010000011001110",
34916 => "1010000011010010",
34917 => "1010000011010110",
34918 => "1010000011011001",
34919 => "1010000011011101",
34920 => "1010000011100001",
34921 => "1010000011100101",
34922 => "1010000011101000",
34923 => "1010000011101100",
34924 => "1010000011110000",
34925 => "1010000011110011",
34926 => "1010000011110111",
34927 => "1010000011111011",
34928 => "1010000011111111",
34929 => "1010000100000010",
34930 => "1010000100000110",
34931 => "1010000100001010",
34932 => "1010000100001110",
34933 => "1010000100010001",
34934 => "1010000100010101",
34935 => "1010000100011001",
34936 => "1010000100011101",
34937 => "1010000100100000",
34938 => "1010000100100100",
34939 => "1010000100101000",
34940 => "1010000100101011",
34941 => "1010000100101111",
34942 => "1010000100110011",
34943 => "1010000100110111",
34944 => "1010000100111010",
34945 => "1010000100111110",
34946 => "1010000101000010",
34947 => "1010000101000110",
34948 => "1010000101001001",
34949 => "1010000101001101",
34950 => "1010000101010001",
34951 => "1010000101010101",
34952 => "1010000101011000",
34953 => "1010000101011100",
34954 => "1010000101100000",
34955 => "1010000101100011",
34956 => "1010000101100111",
34957 => "1010000101101011",
34958 => "1010000101101111",
34959 => "1010000101110010",
34960 => "1010000101110110",
34961 => "1010000101111010",
34962 => "1010000101111110",
34963 => "1010000110000001",
34964 => "1010000110000101",
34965 => "1010000110001001",
34966 => "1010000110001100",
34967 => "1010000110010000",
34968 => "1010000110010100",
34969 => "1010000110011000",
34970 => "1010000110011011",
34971 => "1010000110011111",
34972 => "1010000110100011",
34973 => "1010000110100110",
34974 => "1010000110101010",
34975 => "1010000110101110",
34976 => "1010000110110010",
34977 => "1010000110110101",
34978 => "1010000110111001",
34979 => "1010000110111101",
34980 => "1010000111000001",
34981 => "1010000111000100",
34982 => "1010000111001000",
34983 => "1010000111001100",
34984 => "1010000111001111",
34985 => "1010000111010011",
34986 => "1010000111010111",
34987 => "1010000111011011",
34988 => "1010000111011110",
34989 => "1010000111100010",
34990 => "1010000111100110",
34991 => "1010000111101001",
34992 => "1010000111101101",
34993 => "1010000111110001",
34994 => "1010000111110101",
34995 => "1010000111111000",
34996 => "1010000111111100",
34997 => "1010001000000000",
34998 => "1010001000000011",
34999 => "1010001000000111",
35000 => "1010001000001011",
35001 => "1010001000001111",
35002 => "1010001000010010",
35003 => "1010001000010110",
35004 => "1010001000011010",
35005 => "1010001000011110",
35006 => "1010001000100001",
35007 => "1010001000100101",
35008 => "1010001000101001",
35009 => "1010001000101100",
35010 => "1010001000110000",
35011 => "1010001000110100",
35012 => "1010001000111000",
35013 => "1010001000111011",
35014 => "1010001000111111",
35015 => "1010001001000011",
35016 => "1010001001000110",
35017 => "1010001001001010",
35018 => "1010001001001110",
35019 => "1010001001010010",
35020 => "1010001001010101",
35021 => "1010001001011001",
35022 => "1010001001011101",
35023 => "1010001001100000",
35024 => "1010001001100100",
35025 => "1010001001101000",
35026 => "1010001001101011",
35027 => "1010001001101111",
35028 => "1010001001110011",
35029 => "1010001001110111",
35030 => "1010001001111010",
35031 => "1010001001111110",
35032 => "1010001010000010",
35033 => "1010001010000101",
35034 => "1010001010001001",
35035 => "1010001010001101",
35036 => "1010001010010001",
35037 => "1010001010010100",
35038 => "1010001010011000",
35039 => "1010001010011100",
35040 => "1010001010011111",
35041 => "1010001010100011",
35042 => "1010001010100111",
35043 => "1010001010101011",
35044 => "1010001010101110",
35045 => "1010001010110010",
35046 => "1010001010110110",
35047 => "1010001010111001",
35048 => "1010001010111101",
35049 => "1010001011000001",
35050 => "1010001011000100",
35051 => "1010001011001000",
35052 => "1010001011001100",
35053 => "1010001011010000",
35054 => "1010001011010011",
35055 => "1010001011010111",
35056 => "1010001011011011",
35057 => "1010001011011110",
35058 => "1010001011100010",
35059 => "1010001011100110",
35060 => "1010001011101010",
35061 => "1010001011101101",
35062 => "1010001011110001",
35063 => "1010001011110101",
35064 => "1010001011111000",
35065 => "1010001011111100",
35066 => "1010001100000000",
35067 => "1010001100000011",
35068 => "1010001100000111",
35069 => "1010001100001011",
35070 => "1010001100001111",
35071 => "1010001100010010",
35072 => "1010001100010110",
35073 => "1010001100011010",
35074 => "1010001100011101",
35075 => "1010001100100001",
35076 => "1010001100100101",
35077 => "1010001100101000",
35078 => "1010001100101100",
35079 => "1010001100110000",
35080 => "1010001100110100",
35081 => "1010001100110111",
35082 => "1010001100111011",
35083 => "1010001100111111",
35084 => "1010001101000010",
35085 => "1010001101000110",
35086 => "1010001101001010",
35087 => "1010001101001101",
35088 => "1010001101010001",
35089 => "1010001101010101",
35090 => "1010001101011000",
35091 => "1010001101011100",
35092 => "1010001101100000",
35093 => "1010001101100100",
35094 => "1010001101100111",
35095 => "1010001101101011",
35096 => "1010001101101111",
35097 => "1010001101110010",
35098 => "1010001101110110",
35099 => "1010001101111010",
35100 => "1010001101111101",
35101 => "1010001110000001",
35102 => "1010001110000101",
35103 => "1010001110001000",
35104 => "1010001110001100",
35105 => "1010001110010000",
35106 => "1010001110010100",
35107 => "1010001110010111",
35108 => "1010001110011011",
35109 => "1010001110011111",
35110 => "1010001110100010",
35111 => "1010001110100110",
35112 => "1010001110101010",
35113 => "1010001110101101",
35114 => "1010001110110001",
35115 => "1010001110110101",
35116 => "1010001110111000",
35117 => "1010001110111100",
35118 => "1010001111000000",
35119 => "1010001111000100",
35120 => "1010001111000111",
35121 => "1010001111001011",
35122 => "1010001111001111",
35123 => "1010001111010010",
35124 => "1010001111010110",
35125 => "1010001111011010",
35126 => "1010001111011101",
35127 => "1010001111100001",
35128 => "1010001111100101",
35129 => "1010001111101000",
35130 => "1010001111101100",
35131 => "1010001111110000",
35132 => "1010001111110011",
35133 => "1010001111110111",
35134 => "1010001111111011",
35135 => "1010001111111111",
35136 => "1010010000000010",
35137 => "1010010000000110",
35138 => "1010010000001010",
35139 => "1010010000001101",
35140 => "1010010000010001",
35141 => "1010010000010101",
35142 => "1010010000011000",
35143 => "1010010000011100",
35144 => "1010010000100000",
35145 => "1010010000100011",
35146 => "1010010000100111",
35147 => "1010010000101011",
35148 => "1010010000101110",
35149 => "1010010000110010",
35150 => "1010010000110110",
35151 => "1010010000111001",
35152 => "1010010000111101",
35153 => "1010010001000001",
35154 => "1010010001000100",
35155 => "1010010001001000",
35156 => "1010010001001100",
35157 => "1010010001001111",
35158 => "1010010001010011",
35159 => "1010010001010111",
35160 => "1010010001011011",
35161 => "1010010001011110",
35162 => "1010010001100010",
35163 => "1010010001100110",
35164 => "1010010001101001",
35165 => "1010010001101101",
35166 => "1010010001110001",
35167 => "1010010001110100",
35168 => "1010010001111000",
35169 => "1010010001111100",
35170 => "1010010001111111",
35171 => "1010010010000011",
35172 => "1010010010000111",
35173 => "1010010010001010",
35174 => "1010010010001110",
35175 => "1010010010010010",
35176 => "1010010010010101",
35177 => "1010010010011001",
35178 => "1010010010011101",
35179 => "1010010010100000",
35180 => "1010010010100100",
35181 => "1010010010101000",
35182 => "1010010010101011",
35183 => "1010010010101111",
35184 => "1010010010110011",
35185 => "1010010010110110",
35186 => "1010010010111010",
35187 => "1010010010111110",
35188 => "1010010011000001",
35189 => "1010010011000101",
35190 => "1010010011001001",
35191 => "1010010011001100",
35192 => "1010010011010000",
35193 => "1010010011010100",
35194 => "1010010011010111",
35195 => "1010010011011011",
35196 => "1010010011011111",
35197 => "1010010011100010",
35198 => "1010010011100110",
35199 => "1010010011101010",
35200 => "1010010011101101",
35201 => "1010010011110001",
35202 => "1010010011110101",
35203 => "1010010011111000",
35204 => "1010010011111100",
35205 => "1010010100000000",
35206 => "1010010100000011",
35207 => "1010010100000111",
35208 => "1010010100001011",
35209 => "1010010100001110",
35210 => "1010010100010010",
35211 => "1010010100010110",
35212 => "1010010100011001",
35213 => "1010010100011101",
35214 => "1010010100100001",
35215 => "1010010100100100",
35216 => "1010010100101000",
35217 => "1010010100101100",
35218 => "1010010100101111",
35219 => "1010010100110011",
35220 => "1010010100110111",
35221 => "1010010100111010",
35222 => "1010010100111110",
35223 => "1010010101000010",
35224 => "1010010101000101",
35225 => "1010010101001001",
35226 => "1010010101001101",
35227 => "1010010101010000",
35228 => "1010010101010100",
35229 => "1010010101011000",
35230 => "1010010101011011",
35231 => "1010010101011111",
35232 => "1010010101100011",
35233 => "1010010101100110",
35234 => "1010010101101010",
35235 => "1010010101101110",
35236 => "1010010101110001",
35237 => "1010010101110101",
35238 => "1010010101111001",
35239 => "1010010101111100",
35240 => "1010010110000000",
35241 => "1010010110000100",
35242 => "1010010110000111",
35243 => "1010010110001011",
35244 => "1010010110001111",
35245 => "1010010110010010",
35246 => "1010010110010110",
35247 => "1010010110011001",
35248 => "1010010110011101",
35249 => "1010010110100001",
35250 => "1010010110100100",
35251 => "1010010110101000",
35252 => "1010010110101100",
35253 => "1010010110101111",
35254 => "1010010110110011",
35255 => "1010010110110111",
35256 => "1010010110111010",
35257 => "1010010110111110",
35258 => "1010010111000010",
35259 => "1010010111000101",
35260 => "1010010111001001",
35261 => "1010010111001101",
35262 => "1010010111010000",
35263 => "1010010111010100",
35264 => "1010010111011000",
35265 => "1010010111011011",
35266 => "1010010111011111",
35267 => "1010010111100011",
35268 => "1010010111100110",
35269 => "1010010111101010",
35270 => "1010010111101101",
35271 => "1010010111110001",
35272 => "1010010111110101",
35273 => "1010010111111000",
35274 => "1010010111111100",
35275 => "1010011000000000",
35276 => "1010011000000011",
35277 => "1010011000000111",
35278 => "1010011000001011",
35279 => "1010011000001110",
35280 => "1010011000010010",
35281 => "1010011000010110",
35282 => "1010011000011001",
35283 => "1010011000011101",
35284 => "1010011000100001",
35285 => "1010011000100100",
35286 => "1010011000101000",
35287 => "1010011000101011",
35288 => "1010011000101111",
35289 => "1010011000110011",
35290 => "1010011000110110",
35291 => "1010011000111010",
35292 => "1010011000111110",
35293 => "1010011001000001",
35294 => "1010011001000101",
35295 => "1010011001001001",
35296 => "1010011001001100",
35297 => "1010011001010000",
35298 => "1010011001010100",
35299 => "1010011001010111",
35300 => "1010011001011011",
35301 => "1010011001011110",
35302 => "1010011001100010",
35303 => "1010011001100110",
35304 => "1010011001101001",
35305 => "1010011001101101",
35306 => "1010011001110001",
35307 => "1010011001110100",
35308 => "1010011001111000",
35309 => "1010011001111100",
35310 => "1010011001111111",
35311 => "1010011010000011",
35312 => "1010011010000110",
35313 => "1010011010001010",
35314 => "1010011010001110",
35315 => "1010011010010001",
35316 => "1010011010010101",
35317 => "1010011010011001",
35318 => "1010011010011100",
35319 => "1010011010100000",
35320 => "1010011010100100",
35321 => "1010011010100111",
35322 => "1010011010101011",
35323 => "1010011010101110",
35324 => "1010011010110010",
35325 => "1010011010110110",
35326 => "1010011010111001",
35327 => "1010011010111101",
35328 => "1010011011000001",
35329 => "1010011011000100",
35330 => "1010011011001000",
35331 => "1010011011001100",
35332 => "1010011011001111",
35333 => "1010011011010011",
35334 => "1010011011010110",
35335 => "1010011011011010",
35336 => "1010011011011110",
35337 => "1010011011100001",
35338 => "1010011011100101",
35339 => "1010011011101001",
35340 => "1010011011101100",
35341 => "1010011011110000",
35342 => "1010011011110011",
35343 => "1010011011110111",
35344 => "1010011011111011",
35345 => "1010011011111110",
35346 => "1010011100000010",
35347 => "1010011100000110",
35348 => "1010011100001001",
35349 => "1010011100001101",
35350 => "1010011100010001",
35351 => "1010011100010100",
35352 => "1010011100011000",
35353 => "1010011100011011",
35354 => "1010011100011111",
35355 => "1010011100100011",
35356 => "1010011100100110",
35357 => "1010011100101010",
35358 => "1010011100101110",
35359 => "1010011100110001",
35360 => "1010011100110101",
35361 => "1010011100111000",
35362 => "1010011100111100",
35363 => "1010011101000000",
35364 => "1010011101000011",
35365 => "1010011101000111",
35366 => "1010011101001011",
35367 => "1010011101001110",
35368 => "1010011101010010",
35369 => "1010011101010101",
35370 => "1010011101011001",
35371 => "1010011101011101",
35372 => "1010011101100000",
35373 => "1010011101100100",
35374 => "1010011101101000",
35375 => "1010011101101011",
35376 => "1010011101101111",
35377 => "1010011101110010",
35378 => "1010011101110110",
35379 => "1010011101111010",
35380 => "1010011101111101",
35381 => "1010011110000001",
35382 => "1010011110000100",
35383 => "1010011110001000",
35384 => "1010011110001100",
35385 => "1010011110001111",
35386 => "1010011110010011",
35387 => "1010011110010111",
35388 => "1010011110011010",
35389 => "1010011110011110",
35390 => "1010011110100001",
35391 => "1010011110100101",
35392 => "1010011110101001",
35393 => "1010011110101100",
35394 => "1010011110110000",
35395 => "1010011110110011",
35396 => "1010011110110111",
35397 => "1010011110111011",
35398 => "1010011110111110",
35399 => "1010011111000010",
35400 => "1010011111000110",
35401 => "1010011111001001",
35402 => "1010011111001101",
35403 => "1010011111010000",
35404 => "1010011111010100",
35405 => "1010011111011000",
35406 => "1010011111011011",
35407 => "1010011111011111",
35408 => "1010011111100010",
35409 => "1010011111100110",
35410 => "1010011111101010",
35411 => "1010011111101101",
35412 => "1010011111110001",
35413 => "1010011111110101",
35414 => "1010011111111000",
35415 => "1010011111111100",
35416 => "1010011111111111",
35417 => "1010100000000011",
35418 => "1010100000000111",
35419 => "1010100000001010",
35420 => "1010100000001110",
35421 => "1010100000010001",
35422 => "1010100000010101",
35423 => "1010100000011001",
35424 => "1010100000011100",
35425 => "1010100000100000",
35426 => "1010100000100011",
35427 => "1010100000100111",
35428 => "1010100000101011",
35429 => "1010100000101110",
35430 => "1010100000110010",
35431 => "1010100000110101",
35432 => "1010100000111001",
35433 => "1010100000111101",
35434 => "1010100001000000",
35435 => "1010100001000100",
35436 => "1010100001000111",
35437 => "1010100001001011",
35438 => "1010100001001111",
35439 => "1010100001010010",
35440 => "1010100001010110",
35441 => "1010100001011001",
35442 => "1010100001011101",
35443 => "1010100001100001",
35444 => "1010100001100100",
35445 => "1010100001101000",
35446 => "1010100001101011",
35447 => "1010100001101111",
35448 => "1010100001110011",
35449 => "1010100001110110",
35450 => "1010100001111010",
35451 => "1010100001111110",
35452 => "1010100010000001",
35453 => "1010100010000101",
35454 => "1010100010001000",
35455 => "1010100010001100",
35456 => "1010100010001111",
35457 => "1010100010010011",
35458 => "1010100010010111",
35459 => "1010100010011010",
35460 => "1010100010011110",
35461 => "1010100010100001",
35462 => "1010100010100101",
35463 => "1010100010101001",
35464 => "1010100010101100",
35465 => "1010100010110000",
35466 => "1010100010110011",
35467 => "1010100010110111",
35468 => "1010100010111011",
35469 => "1010100010111110",
35470 => "1010100011000010",
35471 => "1010100011000101",
35472 => "1010100011001001",
35473 => "1010100011001101",
35474 => "1010100011010000",
35475 => "1010100011010100",
35476 => "1010100011010111",
35477 => "1010100011011011",
35478 => "1010100011011111",
35479 => "1010100011100010",
35480 => "1010100011100110",
35481 => "1010100011101001",
35482 => "1010100011101101",
35483 => "1010100011110001",
35484 => "1010100011110100",
35485 => "1010100011111000",
35486 => "1010100011111011",
35487 => "1010100011111111",
35488 => "1010100100000011",
35489 => "1010100100000110",
35490 => "1010100100001010",
35491 => "1010100100001101",
35492 => "1010100100010001",
35493 => "1010100100010100",
35494 => "1010100100011000",
35495 => "1010100100011100",
35496 => "1010100100011111",
35497 => "1010100100100011",
35498 => "1010100100100110",
35499 => "1010100100101010",
35500 => "1010100100101110",
35501 => "1010100100110001",
35502 => "1010100100110101",
35503 => "1010100100111000",
35504 => "1010100100111100",
35505 => "1010100100111111",
35506 => "1010100101000011",
35507 => "1010100101000111",
35508 => "1010100101001010",
35509 => "1010100101001110",
35510 => "1010100101010001",
35511 => "1010100101010101",
35512 => "1010100101011001",
35513 => "1010100101011100",
35514 => "1010100101100000",
35515 => "1010100101100011",
35516 => "1010100101100111",
35517 => "1010100101101010",
35518 => "1010100101101110",
35519 => "1010100101110010",
35520 => "1010100101110101",
35521 => "1010100101111001",
35522 => "1010100101111100",
35523 => "1010100110000000",
35524 => "1010100110000100",
35525 => "1010100110000111",
35526 => "1010100110001011",
35527 => "1010100110001110",
35528 => "1010100110010010",
35529 => "1010100110010101",
35530 => "1010100110011001",
35531 => "1010100110011101",
35532 => "1010100110100000",
35533 => "1010100110100100",
35534 => "1010100110100111",
35535 => "1010100110101011",
35536 => "1010100110101110",
35537 => "1010100110110010",
35538 => "1010100110110110",
35539 => "1010100110111001",
35540 => "1010100110111101",
35541 => "1010100111000000",
35542 => "1010100111000100",
35543 => "1010100111000111",
35544 => "1010100111001011",
35545 => "1010100111001111",
35546 => "1010100111010010",
35547 => "1010100111010110",
35548 => "1010100111011001",
35549 => "1010100111011101",
35550 => "1010100111100001",
35551 => "1010100111100100",
35552 => "1010100111101000",
35553 => "1010100111101011",
35554 => "1010100111101111",
35555 => "1010100111110010",
35556 => "1010100111110110",
35557 => "1010100111111001",
35558 => "1010100111111101",
35559 => "1010101000000001",
35560 => "1010101000000100",
35561 => "1010101000001000",
35562 => "1010101000001011",
35563 => "1010101000001111",
35564 => "1010101000010010",
35565 => "1010101000010110",
35566 => "1010101000011010",
35567 => "1010101000011101",
35568 => "1010101000100001",
35569 => "1010101000100100",
35570 => "1010101000101000",
35571 => "1010101000101011",
35572 => "1010101000101111",
35573 => "1010101000110011",
35574 => "1010101000110110",
35575 => "1010101000111010",
35576 => "1010101000111101",
35577 => "1010101001000001",
35578 => "1010101001000100",
35579 => "1010101001001000",
35580 => "1010101001001100",
35581 => "1010101001001111",
35582 => "1010101001010011",
35583 => "1010101001010110",
35584 => "1010101001011010",
35585 => "1010101001011101",
35586 => "1010101001100001",
35587 => "1010101001100100",
35588 => "1010101001101000",
35589 => "1010101001101100",
35590 => "1010101001101111",
35591 => "1010101001110011",
35592 => "1010101001110110",
35593 => "1010101001111010",
35594 => "1010101001111101",
35595 => "1010101010000001",
35596 => "1010101010000101",
35597 => "1010101010001000",
35598 => "1010101010001100",
35599 => "1010101010001111",
35600 => "1010101010010011",
35601 => "1010101010010110",
35602 => "1010101010011010",
35603 => "1010101010011101",
35604 => "1010101010100001",
35605 => "1010101010100101",
35606 => "1010101010101000",
35607 => "1010101010101100",
35608 => "1010101010101111",
35609 => "1010101010110011",
35610 => "1010101010110110",
35611 => "1010101010111010",
35612 => "1010101010111101",
35613 => "1010101011000001",
35614 => "1010101011000101",
35615 => "1010101011001000",
35616 => "1010101011001100",
35617 => "1010101011001111",
35618 => "1010101011010011",
35619 => "1010101011010110",
35620 => "1010101011011010",
35621 => "1010101011011101",
35622 => "1010101011100001",
35623 => "1010101011100100",
35624 => "1010101011101000",
35625 => "1010101011101100",
35626 => "1010101011101111",
35627 => "1010101011110011",
35628 => "1010101011110110",
35629 => "1010101011111010",
35630 => "1010101011111101",
35631 => "1010101100000001",
35632 => "1010101100000100",
35633 => "1010101100001000",
35634 => "1010101100001100",
35635 => "1010101100001111",
35636 => "1010101100010011",
35637 => "1010101100010110",
35638 => "1010101100011010",
35639 => "1010101100011101",
35640 => "1010101100100001",
35641 => "1010101100100100",
35642 => "1010101100101000",
35643 => "1010101100101011",
35644 => "1010101100101111",
35645 => "1010101100110011",
35646 => "1010101100110110",
35647 => "1010101100111010",
35648 => "1010101100111101",
35649 => "1010101101000001",
35650 => "1010101101000100",
35651 => "1010101101001000",
35652 => "1010101101001011",
35653 => "1010101101001111",
35654 => "1010101101010010",
35655 => "1010101101010110",
35656 => "1010101101011010",
35657 => "1010101101011101",
35658 => "1010101101100001",
35659 => "1010101101100100",
35660 => "1010101101101000",
35661 => "1010101101101011",
35662 => "1010101101101111",
35663 => "1010101101110010",
35664 => "1010101101110110",
35665 => "1010101101111001",
35666 => "1010101101111101",
35667 => "1010101110000000",
35668 => "1010101110000100",
35669 => "1010101110001000",
35670 => "1010101110001011",
35671 => "1010101110001111",
35672 => "1010101110010010",
35673 => "1010101110010110",
35674 => "1010101110011001",
35675 => "1010101110011101",
35676 => "1010101110100000",
35677 => "1010101110100100",
35678 => "1010101110100111",
35679 => "1010101110101011",
35680 => "1010101110101110",
35681 => "1010101110110010",
35682 => "1010101110110101",
35683 => "1010101110111001",
35684 => "1010101110111101",
35685 => "1010101111000000",
35686 => "1010101111000100",
35687 => "1010101111000111",
35688 => "1010101111001011",
35689 => "1010101111001110",
35690 => "1010101111010010",
35691 => "1010101111010101",
35692 => "1010101111011001",
35693 => "1010101111011100",
35694 => "1010101111100000",
35695 => "1010101111100011",
35696 => "1010101111100111",
35697 => "1010101111101010",
35698 => "1010101111101110",
35699 => "1010101111110010",
35700 => "1010101111110101",
35701 => "1010101111111001",
35702 => "1010101111111100",
35703 => "1010110000000000",
35704 => "1010110000000011",
35705 => "1010110000000111",
35706 => "1010110000001010",
35707 => "1010110000001110",
35708 => "1010110000010001",
35709 => "1010110000010101",
35710 => "1010110000011000",
35711 => "1010110000011100",
35712 => "1010110000011111",
35713 => "1010110000100011",
35714 => "1010110000100110",
35715 => "1010110000101010",
35716 => "1010110000101101",
35717 => "1010110000110001",
35718 => "1010110000110100",
35719 => "1010110000111000",
35720 => "1010110000111100",
35721 => "1010110000111111",
35722 => "1010110001000011",
35723 => "1010110001000110",
35724 => "1010110001001010",
35725 => "1010110001001101",
35726 => "1010110001010001",
35727 => "1010110001010100",
35728 => "1010110001011000",
35729 => "1010110001011011",
35730 => "1010110001011111",
35731 => "1010110001100010",
35732 => "1010110001100110",
35733 => "1010110001101001",
35734 => "1010110001101101",
35735 => "1010110001110000",
35736 => "1010110001110100",
35737 => "1010110001110111",
35738 => "1010110001111011",
35739 => "1010110001111110",
35740 => "1010110010000010",
35741 => "1010110010000101",
35742 => "1010110010001001",
35743 => "1010110010001100",
35744 => "1010110010010000",
35745 => "1010110010010100",
35746 => "1010110010010111",
35747 => "1010110010011011",
35748 => "1010110010011110",
35749 => "1010110010100010",
35750 => "1010110010100101",
35751 => "1010110010101001",
35752 => "1010110010101100",
35753 => "1010110010110000",
35754 => "1010110010110011",
35755 => "1010110010110111",
35756 => "1010110010111010",
35757 => "1010110010111110",
35758 => "1010110011000001",
35759 => "1010110011000101",
35760 => "1010110011001000",
35761 => "1010110011001100",
35762 => "1010110011001111",
35763 => "1010110011010011",
35764 => "1010110011010110",
35765 => "1010110011011010",
35766 => "1010110011011101",
35767 => "1010110011100001",
35768 => "1010110011100100",
35769 => "1010110011101000",
35770 => "1010110011101011",
35771 => "1010110011101111",
35772 => "1010110011110010",
35773 => "1010110011110110",
35774 => "1010110011111001",
35775 => "1010110011111101",
35776 => "1010110100000000",
35777 => "1010110100000100",
35778 => "1010110100000111",
35779 => "1010110100001011",
35780 => "1010110100001110",
35781 => "1010110100010010",
35782 => "1010110100010101",
35783 => "1010110100011001",
35784 => "1010110100011100",
35785 => "1010110100100000",
35786 => "1010110100100011",
35787 => "1010110100100111",
35788 => "1010110100101010",
35789 => "1010110100101110",
35790 => "1010110100110001",
35791 => "1010110100110101",
35792 => "1010110100111000",
35793 => "1010110100111100",
35794 => "1010110100111111",
35795 => "1010110101000011",
35796 => "1010110101000110",
35797 => "1010110101001010",
35798 => "1010110101001101",
35799 => "1010110101010001",
35800 => "1010110101010100",
35801 => "1010110101011000",
35802 => "1010110101011011",
35803 => "1010110101011111",
35804 => "1010110101100010",
35805 => "1010110101100110",
35806 => "1010110101101001",
35807 => "1010110101101101",
35808 => "1010110101110000",
35809 => "1010110101110100",
35810 => "1010110101110111",
35811 => "1010110101111011",
35812 => "1010110101111110",
35813 => "1010110110000010",
35814 => "1010110110000101",
35815 => "1010110110001001",
35816 => "1010110110001100",
35817 => "1010110110010000",
35818 => "1010110110010011",
35819 => "1010110110010111",
35820 => "1010110110011010",
35821 => "1010110110011110",
35822 => "1010110110100001",
35823 => "1010110110100101",
35824 => "1010110110101000",
35825 => "1010110110101100",
35826 => "1010110110101111",
35827 => "1010110110110011",
35828 => "1010110110110110",
35829 => "1010110110111010",
35830 => "1010110110111101",
35831 => "1010110111000001",
35832 => "1010110111000100",
35833 => "1010110111001000",
35834 => "1010110111001011",
35835 => "1010110111001111",
35836 => "1010110111010010",
35837 => "1010110111010110",
35838 => "1010110111011001",
35839 => "1010110111011101",
35840 => "1010110111100000",
35841 => "1010110111100100",
35842 => "1010110111100111",
35843 => "1010110111101011",
35844 => "1010110111101110",
35845 => "1010110111110001",
35846 => "1010110111110101",
35847 => "1010110111111000",
35848 => "1010110111111100",
35849 => "1010110111111111",
35850 => "1010111000000011",
35851 => "1010111000000110",
35852 => "1010111000001010",
35853 => "1010111000001101",
35854 => "1010111000010001",
35855 => "1010111000010100",
35856 => "1010111000011000",
35857 => "1010111000011011",
35858 => "1010111000011111",
35859 => "1010111000100010",
35860 => "1010111000100110",
35861 => "1010111000101001",
35862 => "1010111000101101",
35863 => "1010111000110000",
35864 => "1010111000110100",
35865 => "1010111000110111",
35866 => "1010111000111011",
35867 => "1010111000111110",
35868 => "1010111001000010",
35869 => "1010111001000101",
35870 => "1010111001001001",
35871 => "1010111001001100",
35872 => "1010111001001111",
35873 => "1010111001010011",
35874 => "1010111001010110",
35875 => "1010111001011010",
35876 => "1010111001011101",
35877 => "1010111001100001",
35878 => "1010111001100100",
35879 => "1010111001101000",
35880 => "1010111001101011",
35881 => "1010111001101111",
35882 => "1010111001110010",
35883 => "1010111001110110",
35884 => "1010111001111001",
35885 => "1010111001111101",
35886 => "1010111010000000",
35887 => "1010111010000100",
35888 => "1010111010000111",
35889 => "1010111010001011",
35890 => "1010111010001110",
35891 => "1010111010010001",
35892 => "1010111010010101",
35893 => "1010111010011000",
35894 => "1010111010011100",
35895 => "1010111010011111",
35896 => "1010111010100011",
35897 => "1010111010100110",
35898 => "1010111010101010",
35899 => "1010111010101101",
35900 => "1010111010110001",
35901 => "1010111010110100",
35902 => "1010111010111000",
35903 => "1010111010111011",
35904 => "1010111010111111",
35905 => "1010111011000010",
35906 => "1010111011000101",
35907 => "1010111011001001",
35908 => "1010111011001100",
35909 => "1010111011010000",
35910 => "1010111011010011",
35911 => "1010111011010111",
35912 => "1010111011011010",
35913 => "1010111011011110",
35914 => "1010111011100001",
35915 => "1010111011100101",
35916 => "1010111011101000",
35917 => "1010111011101100",
35918 => "1010111011101111",
35919 => "1010111011110011",
35920 => "1010111011110110",
35921 => "1010111011111001",
35922 => "1010111011111101",
35923 => "1010111100000000",
35924 => "1010111100000100",
35925 => "1010111100000111",
35926 => "1010111100001011",
35927 => "1010111100001110",
35928 => "1010111100010010",
35929 => "1010111100010101",
35930 => "1010111100011001",
35931 => "1010111100011100",
35932 => "1010111100011111",
35933 => "1010111100100011",
35934 => "1010111100100110",
35935 => "1010111100101010",
35936 => "1010111100101101",
35937 => "1010111100110001",
35938 => "1010111100110100",
35939 => "1010111100111000",
35940 => "1010111100111011",
35941 => "1010111100111111",
35942 => "1010111101000010",
35943 => "1010111101000110",
35944 => "1010111101001001",
35945 => "1010111101001100",
35946 => "1010111101010000",
35947 => "1010111101010011",
35948 => "1010111101010111",
35949 => "1010111101011010",
35950 => "1010111101011110",
35951 => "1010111101100001",
35952 => "1010111101100101",
35953 => "1010111101101000",
35954 => "1010111101101011",
35955 => "1010111101101111",
35956 => "1010111101110010",
35957 => "1010111101110110",
35958 => "1010111101111001",
35959 => "1010111101111101",
35960 => "1010111110000000",
35961 => "1010111110000100",
35962 => "1010111110000111",
35963 => "1010111110001011",
35964 => "1010111110001110",
35965 => "1010111110010001",
35966 => "1010111110010101",
35967 => "1010111110011000",
35968 => "1010111110011100",
35969 => "1010111110011111",
35970 => "1010111110100011",
35971 => "1010111110100110",
35972 => "1010111110101010",
35973 => "1010111110101101",
35974 => "1010111110110000",
35975 => "1010111110110100",
35976 => "1010111110110111",
35977 => "1010111110111011",
35978 => "1010111110111110",
35979 => "1010111111000010",
35980 => "1010111111000101",
35981 => "1010111111001001",
35982 => "1010111111001100",
35983 => "1010111111001111",
35984 => "1010111111010011",
35985 => "1010111111010110",
35986 => "1010111111011010",
35987 => "1010111111011101",
35988 => "1010111111100001",
35989 => "1010111111100100",
35990 => "1010111111101000",
35991 => "1010111111101011",
35992 => "1010111111101110",
35993 => "1010111111110010",
35994 => "1010111111110101",
35995 => "1010111111111001",
35996 => "1010111111111100",
35997 => "1011000000000000",
35998 => "1011000000000011",
35999 => "1011000000000110",
36000 => "1011000000001010",
36001 => "1011000000001101",
36002 => "1011000000010001",
36003 => "1011000000010100",
36004 => "1011000000011000",
36005 => "1011000000011011",
36006 => "1011000000011111",
36007 => "1011000000100010",
36008 => "1011000000100101",
36009 => "1011000000101001",
36010 => "1011000000101100",
36011 => "1011000000110000",
36012 => "1011000000110011",
36013 => "1011000000110111",
36014 => "1011000000111010",
36015 => "1011000000111101",
36016 => "1011000001000001",
36017 => "1011000001000100",
36018 => "1011000001001000",
36019 => "1011000001001011",
36020 => "1011000001001111",
36021 => "1011000001010010",
36022 => "1011000001010101",
36023 => "1011000001011001",
36024 => "1011000001011100",
36025 => "1011000001100000",
36026 => "1011000001100011",
36027 => "1011000001100111",
36028 => "1011000001101010",
36029 => "1011000001101101",
36030 => "1011000001110001",
36031 => "1011000001110100",
36032 => "1011000001111000",
36033 => "1011000001111011",
36034 => "1011000001111111",
36035 => "1011000010000010",
36036 => "1011000010000101",
36037 => "1011000010001001",
36038 => "1011000010001100",
36039 => "1011000010010000",
36040 => "1011000010010011",
36041 => "1011000010010111",
36042 => "1011000010011010",
36043 => "1011000010011101",
36044 => "1011000010100001",
36045 => "1011000010100100",
36046 => "1011000010101000",
36047 => "1011000010101011",
36048 => "1011000010101111",
36049 => "1011000010110010",
36050 => "1011000010110101",
36051 => "1011000010111001",
36052 => "1011000010111100",
36053 => "1011000011000000",
36054 => "1011000011000011",
36055 => "1011000011000110",
36056 => "1011000011001010",
36057 => "1011000011001101",
36058 => "1011000011010001",
36059 => "1011000011010100",
36060 => "1011000011011000",
36061 => "1011000011011011",
36062 => "1011000011011110",
36063 => "1011000011100010",
36064 => "1011000011100101",
36065 => "1011000011101001",
36066 => "1011000011101100",
36067 => "1011000011101111",
36068 => "1011000011110011",
36069 => "1011000011110110",
36070 => "1011000011111010",
36071 => "1011000011111101",
36072 => "1011000100000001",
36073 => "1011000100000100",
36074 => "1011000100000111",
36075 => "1011000100001011",
36076 => "1011000100001110",
36077 => "1011000100010010",
36078 => "1011000100010101",
36079 => "1011000100011000",
36080 => "1011000100011100",
36081 => "1011000100011111",
36082 => "1011000100100011",
36083 => "1011000100100110",
36084 => "1011000100101001",
36085 => "1011000100101101",
36086 => "1011000100110000",
36087 => "1011000100110100",
36088 => "1011000100110111",
36089 => "1011000100111011",
36090 => "1011000100111110",
36091 => "1011000101000001",
36092 => "1011000101000101",
36093 => "1011000101001000",
36094 => "1011000101001100",
36095 => "1011000101001111",
36096 => "1011000101010010",
36097 => "1011000101010110",
36098 => "1011000101011001",
36099 => "1011000101011101",
36100 => "1011000101100000",
36101 => "1011000101100011",
36102 => "1011000101100111",
36103 => "1011000101101010",
36104 => "1011000101101110",
36105 => "1011000101110001",
36106 => "1011000101110100",
36107 => "1011000101111000",
36108 => "1011000101111011",
36109 => "1011000101111111",
36110 => "1011000110000010",
36111 => "1011000110000101",
36112 => "1011000110001001",
36113 => "1011000110001100",
36114 => "1011000110010000",
36115 => "1011000110010011",
36116 => "1011000110010110",
36117 => "1011000110011010",
36118 => "1011000110011101",
36119 => "1011000110100001",
36120 => "1011000110100100",
36121 => "1011000110100111",
36122 => "1011000110101011",
36123 => "1011000110101110",
36124 => "1011000110110010",
36125 => "1011000110110101",
36126 => "1011000110111000",
36127 => "1011000110111100",
36128 => "1011000110111111",
36129 => "1011000111000011",
36130 => "1011000111000110",
36131 => "1011000111001001",
36132 => "1011000111001101",
36133 => "1011000111010000",
36134 => "1011000111010100",
36135 => "1011000111010111",
36136 => "1011000111011010",
36137 => "1011000111011110",
36138 => "1011000111100001",
36139 => "1011000111100101",
36140 => "1011000111101000",
36141 => "1011000111101011",
36142 => "1011000111101111",
36143 => "1011000111110010",
36144 => "1011000111110101",
36145 => "1011000111111001",
36146 => "1011000111111100",
36147 => "1011001000000000",
36148 => "1011001000000011",
36149 => "1011001000000110",
36150 => "1011001000001010",
36151 => "1011001000001101",
36152 => "1011001000010001",
36153 => "1011001000010100",
36154 => "1011001000010111",
36155 => "1011001000011011",
36156 => "1011001000011110",
36157 => "1011001000100010",
36158 => "1011001000100101",
36159 => "1011001000101000",
36160 => "1011001000101100",
36161 => "1011001000101111",
36162 => "1011001000110010",
36163 => "1011001000110110",
36164 => "1011001000111001",
36165 => "1011001000111101",
36166 => "1011001001000000",
36167 => "1011001001000011",
36168 => "1011001001000111",
36169 => "1011001001001010",
36170 => "1011001001001110",
36171 => "1011001001010001",
36172 => "1011001001010100",
36173 => "1011001001011000",
36174 => "1011001001011011",
36175 => "1011001001011110",
36176 => "1011001001100010",
36177 => "1011001001100101",
36178 => "1011001001101001",
36179 => "1011001001101100",
36180 => "1011001001101111",
36181 => "1011001001110011",
36182 => "1011001001110110",
36183 => "1011001001111001",
36184 => "1011001001111101",
36185 => "1011001010000000",
36186 => "1011001010000100",
36187 => "1011001010000111",
36188 => "1011001010001010",
36189 => "1011001010001110",
36190 => "1011001010010001",
36191 => "1011001010010100",
36192 => "1011001010011000",
36193 => "1011001010011011",
36194 => "1011001010011111",
36195 => "1011001010100010",
36196 => "1011001010100101",
36197 => "1011001010101001",
36198 => "1011001010101100",
36199 => "1011001010101111",
36200 => "1011001010110011",
36201 => "1011001010110110",
36202 => "1011001010111010",
36203 => "1011001010111101",
36204 => "1011001011000000",
36205 => "1011001011000100",
36206 => "1011001011000111",
36207 => "1011001011001010",
36208 => "1011001011001110",
36209 => "1011001011010001",
36210 => "1011001011010101",
36211 => "1011001011011000",
36212 => "1011001011011011",
36213 => "1011001011011111",
36214 => "1011001011100010",
36215 => "1011001011100101",
36216 => "1011001011101001",
36217 => "1011001011101100",
36218 => "1011001011110000",
36219 => "1011001011110011",
36220 => "1011001011110110",
36221 => "1011001011111010",
36222 => "1011001011111101",
36223 => "1011001100000000",
36224 => "1011001100000100",
36225 => "1011001100000111",
36226 => "1011001100001010",
36227 => "1011001100001110",
36228 => "1011001100010001",
36229 => "1011001100010101",
36230 => "1011001100011000",
36231 => "1011001100011011",
36232 => "1011001100011111",
36233 => "1011001100100010",
36234 => "1011001100100101",
36235 => "1011001100101001",
36236 => "1011001100101100",
36237 => "1011001100101111",
36238 => "1011001100110011",
36239 => "1011001100110110",
36240 => "1011001100111001",
36241 => "1011001100111101",
36242 => "1011001101000000",
36243 => "1011001101000100",
36244 => "1011001101000111",
36245 => "1011001101001010",
36246 => "1011001101001110",
36247 => "1011001101010001",
36248 => "1011001101010100",
36249 => "1011001101011000",
36250 => "1011001101011011",
36251 => "1011001101011110",
36252 => "1011001101100010",
36253 => "1011001101100101",
36254 => "1011001101101000",
36255 => "1011001101101100",
36256 => "1011001101101111",
36257 => "1011001101110011",
36258 => "1011001101110110",
36259 => "1011001101111001",
36260 => "1011001101111101",
36261 => "1011001110000000",
36262 => "1011001110000011",
36263 => "1011001110000111",
36264 => "1011001110001010",
36265 => "1011001110001101",
36266 => "1011001110010001",
36267 => "1011001110010100",
36268 => "1011001110010111",
36269 => "1011001110011011",
36270 => "1011001110011110",
36271 => "1011001110100001",
36272 => "1011001110100101",
36273 => "1011001110101000",
36274 => "1011001110101100",
36275 => "1011001110101111",
36276 => "1011001110110010",
36277 => "1011001110110110",
36278 => "1011001110111001",
36279 => "1011001110111100",
36280 => "1011001111000000",
36281 => "1011001111000011",
36282 => "1011001111000110",
36283 => "1011001111001010",
36284 => "1011001111001101",
36285 => "1011001111010000",
36286 => "1011001111010100",
36287 => "1011001111010111",
36288 => "1011001111011010",
36289 => "1011001111011110",
36290 => "1011001111100001",
36291 => "1011001111100100",
36292 => "1011001111101000",
36293 => "1011001111101011",
36294 => "1011001111101110",
36295 => "1011001111110010",
36296 => "1011001111110101",
36297 => "1011001111111000",
36298 => "1011001111111100",
36299 => "1011001111111111",
36300 => "1011010000000010",
36301 => "1011010000000110",
36302 => "1011010000001001",
36303 => "1011010000001100",
36304 => "1011010000010000",
36305 => "1011010000010011",
36306 => "1011010000010110",
36307 => "1011010000011010",
36308 => "1011010000011101",
36309 => "1011010000100001",
36310 => "1011010000100100",
36311 => "1011010000100111",
36312 => "1011010000101011",
36313 => "1011010000101110",
36314 => "1011010000110001",
36315 => "1011010000110101",
36316 => "1011010000111000",
36317 => "1011010000111011",
36318 => "1011010000111111",
36319 => "1011010001000010",
36320 => "1011010001000101",
36321 => "1011010001001001",
36322 => "1011010001001100",
36323 => "1011010001001111",
36324 => "1011010001010011",
36325 => "1011010001010110",
36326 => "1011010001011001",
36327 => "1011010001011101",
36328 => "1011010001100000",
36329 => "1011010001100011",
36330 => "1011010001100110",
36331 => "1011010001101010",
36332 => "1011010001101101",
36333 => "1011010001110000",
36334 => "1011010001110100",
36335 => "1011010001110111",
36336 => "1011010001111010",
36337 => "1011010001111110",
36338 => "1011010010000001",
36339 => "1011010010000100",
36340 => "1011010010001000",
36341 => "1011010010001011",
36342 => "1011010010001110",
36343 => "1011010010010010",
36344 => "1011010010010101",
36345 => "1011010010011000",
36346 => "1011010010011100",
36347 => "1011010010011111",
36348 => "1011010010100010",
36349 => "1011010010100110",
36350 => "1011010010101001",
36351 => "1011010010101100",
36352 => "1011010010110000",
36353 => "1011010010110011",
36354 => "1011010010110110",
36355 => "1011010010111010",
36356 => "1011010010111101",
36357 => "1011010011000000",
36358 => "1011010011000100",
36359 => "1011010011000111",
36360 => "1011010011001010",
36361 => "1011010011001110",
36362 => "1011010011010001",
36363 => "1011010011010100",
36364 => "1011010011011000",
36365 => "1011010011011011",
36366 => "1011010011011110",
36367 => "1011010011100001",
36368 => "1011010011100101",
36369 => "1011010011101000",
36370 => "1011010011101011",
36371 => "1011010011101111",
36372 => "1011010011110010",
36373 => "1011010011110101",
36374 => "1011010011111001",
36375 => "1011010011111100",
36376 => "1011010011111111",
36377 => "1011010100000011",
36378 => "1011010100000110",
36379 => "1011010100001001",
36380 => "1011010100001101",
36381 => "1011010100010000",
36382 => "1011010100010011",
36383 => "1011010100010111",
36384 => "1011010100011010",
36385 => "1011010100011101",
36386 => "1011010100100000",
36387 => "1011010100100100",
36388 => "1011010100100111",
36389 => "1011010100101010",
36390 => "1011010100101110",
36391 => "1011010100110001",
36392 => "1011010100110100",
36393 => "1011010100111000",
36394 => "1011010100111011",
36395 => "1011010100111110",
36396 => "1011010101000010",
36397 => "1011010101000101",
36398 => "1011010101001000",
36399 => "1011010101001011",
36400 => "1011010101001111",
36401 => "1011010101010010",
36402 => "1011010101010101",
36403 => "1011010101011001",
36404 => "1011010101011100",
36405 => "1011010101011111",
36406 => "1011010101100011",
36407 => "1011010101100110",
36408 => "1011010101101001",
36409 => "1011010101101100",
36410 => "1011010101110000",
36411 => "1011010101110011",
36412 => "1011010101110110",
36413 => "1011010101111010",
36414 => "1011010101111101",
36415 => "1011010110000000",
36416 => "1011010110000100",
36417 => "1011010110000111",
36418 => "1011010110001010",
36419 => "1011010110001110",
36420 => "1011010110010001",
36421 => "1011010110010100",
36422 => "1011010110010111",
36423 => "1011010110011011",
36424 => "1011010110011110",
36425 => "1011010110100001",
36426 => "1011010110100101",
36427 => "1011010110101000",
36428 => "1011010110101011",
36429 => "1011010110101110",
36430 => "1011010110110010",
36431 => "1011010110110101",
36432 => "1011010110111000",
36433 => "1011010110111100",
36434 => "1011010110111111",
36435 => "1011010111000010",
36436 => "1011010111000110",
36437 => "1011010111001001",
36438 => "1011010111001100",
36439 => "1011010111001111",
36440 => "1011010111010011",
36441 => "1011010111010110",
36442 => "1011010111011001",
36443 => "1011010111011101",
36444 => "1011010111100000",
36445 => "1011010111100011",
36446 => "1011010111100110",
36447 => "1011010111101010",
36448 => "1011010111101101",
36449 => "1011010111110000",
36450 => "1011010111110100",
36451 => "1011010111110111",
36452 => "1011010111111010",
36453 => "1011010111111110",
36454 => "1011011000000001",
36455 => "1011011000000100",
36456 => "1011011000000111",
36457 => "1011011000001011",
36458 => "1011011000001110",
36459 => "1011011000010001",
36460 => "1011011000010101",
36461 => "1011011000011000",
36462 => "1011011000011011",
36463 => "1011011000011110",
36464 => "1011011000100010",
36465 => "1011011000100101",
36466 => "1011011000101000",
36467 => "1011011000101100",
36468 => "1011011000101111",
36469 => "1011011000110010",
36470 => "1011011000110101",
36471 => "1011011000111001",
36472 => "1011011000111100",
36473 => "1011011000111111",
36474 => "1011011001000010",
36475 => "1011011001000110",
36476 => "1011011001001001",
36477 => "1011011001001100",
36478 => "1011011001010000",
36479 => "1011011001010011",
36480 => "1011011001010110",
36481 => "1011011001011001",
36482 => "1011011001011101",
36483 => "1011011001100000",
36484 => "1011011001100011",
36485 => "1011011001100111",
36486 => "1011011001101010",
36487 => "1011011001101101",
36488 => "1011011001110000",
36489 => "1011011001110100",
36490 => "1011011001110111",
36491 => "1011011001111010",
36492 => "1011011001111101",
36493 => "1011011010000001",
36494 => "1011011010000100",
36495 => "1011011010000111",
36496 => "1011011010001011",
36497 => "1011011010001110",
36498 => "1011011010010001",
36499 => "1011011010010100",
36500 => "1011011010011000",
36501 => "1011011010011011",
36502 => "1011011010011110",
36503 => "1011011010100010",
36504 => "1011011010100101",
36505 => "1011011010101000",
36506 => "1011011010101011",
36507 => "1011011010101111",
36508 => "1011011010110010",
36509 => "1011011010110101",
36510 => "1011011010111000",
36511 => "1011011010111100",
36512 => "1011011010111111",
36513 => "1011011011000010",
36514 => "1011011011000101",
36515 => "1011011011001001",
36516 => "1011011011001100",
36517 => "1011011011001111",
36518 => "1011011011010011",
36519 => "1011011011010110",
36520 => "1011011011011001",
36521 => "1011011011011100",
36522 => "1011011011100000",
36523 => "1011011011100011",
36524 => "1011011011100110",
36525 => "1011011011101001",
36526 => "1011011011101101",
36527 => "1011011011110000",
36528 => "1011011011110011",
36529 => "1011011011110110",
36530 => "1011011011111010",
36531 => "1011011011111101",
36532 => "1011011100000000",
36533 => "1011011100000011",
36534 => "1011011100000111",
36535 => "1011011100001010",
36536 => "1011011100001101",
36537 => "1011011100010001",
36538 => "1011011100010100",
36539 => "1011011100010111",
36540 => "1011011100011010",
36541 => "1011011100011110",
36542 => "1011011100100001",
36543 => "1011011100100100",
36544 => "1011011100100111",
36545 => "1011011100101011",
36546 => "1011011100101110",
36547 => "1011011100110001",
36548 => "1011011100110100",
36549 => "1011011100111000",
36550 => "1011011100111011",
36551 => "1011011100111110",
36552 => "1011011101000001",
36553 => "1011011101000101",
36554 => "1011011101001000",
36555 => "1011011101001011",
36556 => "1011011101001110",
36557 => "1011011101010010",
36558 => "1011011101010101",
36559 => "1011011101011000",
36560 => "1011011101011011",
36561 => "1011011101011111",
36562 => "1011011101100010",
36563 => "1011011101100101",
36564 => "1011011101101000",
36565 => "1011011101101100",
36566 => "1011011101101111",
36567 => "1011011101110010",
36568 => "1011011101110101",
36569 => "1011011101111001",
36570 => "1011011101111100",
36571 => "1011011101111111",
36572 => "1011011110000010",
36573 => "1011011110000110",
36574 => "1011011110001001",
36575 => "1011011110001100",
36576 => "1011011110001111",
36577 => "1011011110010011",
36578 => "1011011110010110",
36579 => "1011011110011001",
36580 => "1011011110011100",
36581 => "1011011110100000",
36582 => "1011011110100011",
36583 => "1011011110100110",
36584 => "1011011110101001",
36585 => "1011011110101101",
36586 => "1011011110110000",
36587 => "1011011110110011",
36588 => "1011011110110110",
36589 => "1011011110111010",
36590 => "1011011110111101",
36591 => "1011011111000000",
36592 => "1011011111000011",
36593 => "1011011111000111",
36594 => "1011011111001010",
36595 => "1011011111001101",
36596 => "1011011111010000",
36597 => "1011011111010011",
36598 => "1011011111010111",
36599 => "1011011111011010",
36600 => "1011011111011101",
36601 => "1011011111100000",
36602 => "1011011111100100",
36603 => "1011011111100111",
36604 => "1011011111101010",
36605 => "1011011111101101",
36606 => "1011011111110001",
36607 => "1011011111110100",
36608 => "1011011111110111",
36609 => "1011011111111010",
36610 => "1011011111111110",
36611 => "1011100000000001",
36612 => "1011100000000100",
36613 => "1011100000000111",
36614 => "1011100000001011",
36615 => "1011100000001110",
36616 => "1011100000010001",
36617 => "1011100000010100",
36618 => "1011100000010111",
36619 => "1011100000011011",
36620 => "1011100000011110",
36621 => "1011100000100001",
36622 => "1011100000100100",
36623 => "1011100000101000",
36624 => "1011100000101011",
36625 => "1011100000101110",
36626 => "1011100000110001",
36627 => "1011100000110101",
36628 => "1011100000111000",
36629 => "1011100000111011",
36630 => "1011100000111110",
36631 => "1011100001000001",
36632 => "1011100001000101",
36633 => "1011100001001000",
36634 => "1011100001001011",
36635 => "1011100001001110",
36636 => "1011100001010010",
36637 => "1011100001010101",
36638 => "1011100001011000",
36639 => "1011100001011011",
36640 => "1011100001011110",
36641 => "1011100001100010",
36642 => "1011100001100101",
36643 => "1011100001101000",
36644 => "1011100001101011",
36645 => "1011100001101111",
36646 => "1011100001110010",
36647 => "1011100001110101",
36648 => "1011100001111000",
36649 => "1011100001111011",
36650 => "1011100001111111",
36651 => "1011100010000010",
36652 => "1011100010000101",
36653 => "1011100010001000",
36654 => "1011100010001100",
36655 => "1011100010001111",
36656 => "1011100010010010",
36657 => "1011100010010101",
36658 => "1011100010011000",
36659 => "1011100010011100",
36660 => "1011100010011111",
36661 => "1011100010100010",
36662 => "1011100010100101",
36663 => "1011100010101001",
36664 => "1011100010101100",
36665 => "1011100010101111",
36666 => "1011100010110010",
36667 => "1011100010110101",
36668 => "1011100010111001",
36669 => "1011100010111100",
36670 => "1011100010111111",
36671 => "1011100011000010",
36672 => "1011100011000101",
36673 => "1011100011001001",
36674 => "1011100011001100",
36675 => "1011100011001111",
36676 => "1011100011010010",
36677 => "1011100011010110",
36678 => "1011100011011001",
36679 => "1011100011011100",
36680 => "1011100011011111",
36681 => "1011100011100010",
36682 => "1011100011100110",
36683 => "1011100011101001",
36684 => "1011100011101100",
36685 => "1011100011101111",
36686 => "1011100011110010",
36687 => "1011100011110110",
36688 => "1011100011111001",
36689 => "1011100011111100",
36690 => "1011100011111111",
36691 => "1011100100000010",
36692 => "1011100100000110",
36693 => "1011100100001001",
36694 => "1011100100001100",
36695 => "1011100100001111",
36696 => "1011100100010010",
36697 => "1011100100010110",
36698 => "1011100100011001",
36699 => "1011100100011100",
36700 => "1011100100011111",
36701 => "1011100100100010",
36702 => "1011100100100110",
36703 => "1011100100101001",
36704 => "1011100100101100",
36705 => "1011100100101111",
36706 => "1011100100110011",
36707 => "1011100100110110",
36708 => "1011100100111001",
36709 => "1011100100111100",
36710 => "1011100100111111",
36711 => "1011100101000011",
36712 => "1011100101000110",
36713 => "1011100101001001",
36714 => "1011100101001100",
36715 => "1011100101001111",
36716 => "1011100101010011",
36717 => "1011100101010110",
36718 => "1011100101011001",
36719 => "1011100101011100",
36720 => "1011100101011111",
36721 => "1011100101100010",
36722 => "1011100101100110",
36723 => "1011100101101001",
36724 => "1011100101101100",
36725 => "1011100101101111",
36726 => "1011100101110010",
36727 => "1011100101110110",
36728 => "1011100101111001",
36729 => "1011100101111100",
36730 => "1011100101111111",
36731 => "1011100110000010",
36732 => "1011100110000110",
36733 => "1011100110001001",
36734 => "1011100110001100",
36735 => "1011100110001111",
36736 => "1011100110010010",
36737 => "1011100110010110",
36738 => "1011100110011001",
36739 => "1011100110011100",
36740 => "1011100110011111",
36741 => "1011100110100010",
36742 => "1011100110100110",
36743 => "1011100110101001",
36744 => "1011100110101100",
36745 => "1011100110101111",
36746 => "1011100110110010",
36747 => "1011100110110101",
36748 => "1011100110111001",
36749 => "1011100110111100",
36750 => "1011100110111111",
36751 => "1011100111000010",
36752 => "1011100111000101",
36753 => "1011100111001001",
36754 => "1011100111001100",
36755 => "1011100111001111",
36756 => "1011100111010010",
36757 => "1011100111010101",
36758 => "1011100111011000",
36759 => "1011100111011100",
36760 => "1011100111011111",
36761 => "1011100111100010",
36762 => "1011100111100101",
36763 => "1011100111101000",
36764 => "1011100111101100",
36765 => "1011100111101111",
36766 => "1011100111110010",
36767 => "1011100111110101",
36768 => "1011100111111000",
36769 => "1011100111111011",
36770 => "1011100111111111",
36771 => "1011101000000010",
36772 => "1011101000000101",
36773 => "1011101000001000",
36774 => "1011101000001011",
36775 => "1011101000001111",
36776 => "1011101000010010",
36777 => "1011101000010101",
36778 => "1011101000011000",
36779 => "1011101000011011",
36780 => "1011101000011110",
36781 => "1011101000100010",
36782 => "1011101000100101",
36783 => "1011101000101000",
36784 => "1011101000101011",
36785 => "1011101000101110",
36786 => "1011101000110001",
36787 => "1011101000110101",
36788 => "1011101000111000",
36789 => "1011101000111011",
36790 => "1011101000111110",
36791 => "1011101001000001",
36792 => "1011101001000101",
36793 => "1011101001001000",
36794 => "1011101001001011",
36795 => "1011101001001110",
36796 => "1011101001010001",
36797 => "1011101001010100",
36798 => "1011101001011000",
36799 => "1011101001011011",
36800 => "1011101001011110",
36801 => "1011101001100001",
36802 => "1011101001100100",
36803 => "1011101001100111",
36804 => "1011101001101011",
36805 => "1011101001101110",
36806 => "1011101001110001",
36807 => "1011101001110100",
36808 => "1011101001110111",
36809 => "1011101001111010",
36810 => "1011101001111110",
36811 => "1011101010000001",
36812 => "1011101010000100",
36813 => "1011101010000111",
36814 => "1011101010001010",
36815 => "1011101010001101",
36816 => "1011101010010001",
36817 => "1011101010010100",
36818 => "1011101010010111",
36819 => "1011101010011010",
36820 => "1011101010011101",
36821 => "1011101010100000",
36822 => "1011101010100011",
36823 => "1011101010100111",
36824 => "1011101010101010",
36825 => "1011101010101101",
36826 => "1011101010110000",
36827 => "1011101010110011",
36828 => "1011101010110110",
36829 => "1011101010111010",
36830 => "1011101010111101",
36831 => "1011101011000000",
36832 => "1011101011000011",
36833 => "1011101011000110",
36834 => "1011101011001001",
36835 => "1011101011001101",
36836 => "1011101011010000",
36837 => "1011101011010011",
36838 => "1011101011010110",
36839 => "1011101011011001",
36840 => "1011101011011100",
36841 => "1011101011011111",
36842 => "1011101011100011",
36843 => "1011101011100110",
36844 => "1011101011101001",
36845 => "1011101011101100",
36846 => "1011101011101111",
36847 => "1011101011110010",
36848 => "1011101011110110",
36849 => "1011101011111001",
36850 => "1011101011111100",
36851 => "1011101011111111",
36852 => "1011101100000010",
36853 => "1011101100000101",
36854 => "1011101100001000",
36855 => "1011101100001100",
36856 => "1011101100001111",
36857 => "1011101100010010",
36858 => "1011101100010101",
36859 => "1011101100011000",
36860 => "1011101100011011",
36861 => "1011101100011110",
36862 => "1011101100100010",
36863 => "1011101100100101",
36864 => "1011101100101000",
36865 => "1011101100101011",
36866 => "1011101100101110",
36867 => "1011101100110001",
36868 => "1011101100110101",
36869 => "1011101100111000",
36870 => "1011101100111011",
36871 => "1011101100111110",
36872 => "1011101101000001",
36873 => "1011101101000100",
36874 => "1011101101000111",
36875 => "1011101101001011",
36876 => "1011101101001110",
36877 => "1011101101010001",
36878 => "1011101101010100",
36879 => "1011101101010111",
36880 => "1011101101011010",
36881 => "1011101101011101",
36882 => "1011101101100000",
36883 => "1011101101100100",
36884 => "1011101101100111",
36885 => "1011101101101010",
36886 => "1011101101101101",
36887 => "1011101101110000",
36888 => "1011101101110011",
36889 => "1011101101110110",
36890 => "1011101101111010",
36891 => "1011101101111101",
36892 => "1011101110000000",
36893 => "1011101110000011",
36894 => "1011101110000110",
36895 => "1011101110001001",
36896 => "1011101110001100",
36897 => "1011101110010000",
36898 => "1011101110010011",
36899 => "1011101110010110",
36900 => "1011101110011001",
36901 => "1011101110011100",
36902 => "1011101110011111",
36903 => "1011101110100010",
36904 => "1011101110100101",
36905 => "1011101110101001",
36906 => "1011101110101100",
36907 => "1011101110101111",
36908 => "1011101110110010",
36909 => "1011101110110101",
36910 => "1011101110111000",
36911 => "1011101110111011",
36912 => "1011101110111111",
36913 => "1011101111000010",
36914 => "1011101111000101",
36915 => "1011101111001000",
36916 => "1011101111001011",
36917 => "1011101111001110",
36918 => "1011101111010001",
36919 => "1011101111010100",
36920 => "1011101111011000",
36921 => "1011101111011011",
36922 => "1011101111011110",
36923 => "1011101111100001",
36924 => "1011101111100100",
36925 => "1011101111100111",
36926 => "1011101111101010",
36927 => "1011101111101101",
36928 => "1011101111110001",
36929 => "1011101111110100",
36930 => "1011101111110111",
36931 => "1011101111111010",
36932 => "1011101111111101",
36933 => "1011110000000000",
36934 => "1011110000000011",
36935 => "1011110000000110",
36936 => "1011110000001001",
36937 => "1011110000001101",
36938 => "1011110000010000",
36939 => "1011110000010011",
36940 => "1011110000010110",
36941 => "1011110000011001",
36942 => "1011110000011100",
36943 => "1011110000011111",
36944 => "1011110000100010",
36945 => "1011110000100110",
36946 => "1011110000101001",
36947 => "1011110000101100",
36948 => "1011110000101111",
36949 => "1011110000110010",
36950 => "1011110000110101",
36951 => "1011110000111000",
36952 => "1011110000111011",
36953 => "1011110000111110",
36954 => "1011110001000010",
36955 => "1011110001000101",
36956 => "1011110001001000",
36957 => "1011110001001011",
36958 => "1011110001001110",
36959 => "1011110001010001",
36960 => "1011110001010100",
36961 => "1011110001010111",
36962 => "1011110001011010",
36963 => "1011110001011110",
36964 => "1011110001100001",
36965 => "1011110001100100",
36966 => "1011110001100111",
36967 => "1011110001101010",
36968 => "1011110001101101",
36969 => "1011110001110000",
36970 => "1011110001110011",
36971 => "1011110001110110",
36972 => "1011110001111010",
36973 => "1011110001111101",
36974 => "1011110010000000",
36975 => "1011110010000011",
36976 => "1011110010000110",
36977 => "1011110010001001",
36978 => "1011110010001100",
36979 => "1011110010001111",
36980 => "1011110010010010",
36981 => "1011110010010110",
36982 => "1011110010011001",
36983 => "1011110010011100",
36984 => "1011110010011111",
36985 => "1011110010100010",
36986 => "1011110010100101",
36987 => "1011110010101000",
36988 => "1011110010101011",
36989 => "1011110010101110",
36990 => "1011110010110001",
36991 => "1011110010110101",
36992 => "1011110010111000",
36993 => "1011110010111011",
36994 => "1011110010111110",
36995 => "1011110011000001",
36996 => "1011110011000100",
36997 => "1011110011000111",
36998 => "1011110011001010",
36999 => "1011110011001101",
37000 => "1011110011010000",
37001 => "1011110011010100",
37002 => "1011110011010111",
37003 => "1011110011011010",
37004 => "1011110011011101",
37005 => "1011110011100000",
37006 => "1011110011100011",
37007 => "1011110011100110",
37008 => "1011110011101001",
37009 => "1011110011101100",
37010 => "1011110011101111",
37011 => "1011110011110010",
37012 => "1011110011110110",
37013 => "1011110011111001",
37014 => "1011110011111100",
37015 => "1011110011111111",
37016 => "1011110100000010",
37017 => "1011110100000101",
37018 => "1011110100001000",
37019 => "1011110100001011",
37020 => "1011110100001110",
37021 => "1011110100010001",
37022 => "1011110100010100",
37023 => "1011110100011000",
37024 => "1011110100011011",
37025 => "1011110100011110",
37026 => "1011110100100001",
37027 => "1011110100100100",
37028 => "1011110100100111",
37029 => "1011110100101010",
37030 => "1011110100101101",
37031 => "1011110100110000",
37032 => "1011110100110011",
37033 => "1011110100110110",
37034 => "1011110100111010",
37035 => "1011110100111101",
37036 => "1011110101000000",
37037 => "1011110101000011",
37038 => "1011110101000110",
37039 => "1011110101001001",
37040 => "1011110101001100",
37041 => "1011110101001111",
37042 => "1011110101010010",
37043 => "1011110101010101",
37044 => "1011110101011000",
37045 => "1011110101011011",
37046 => "1011110101011111",
37047 => "1011110101100010",
37048 => "1011110101100101",
37049 => "1011110101101000",
37050 => "1011110101101011",
37051 => "1011110101101110",
37052 => "1011110101110001",
37053 => "1011110101110100",
37054 => "1011110101110111",
37055 => "1011110101111010",
37056 => "1011110101111101",
37057 => "1011110110000000",
37058 => "1011110110000011",
37059 => "1011110110000111",
37060 => "1011110110001010",
37061 => "1011110110001101",
37062 => "1011110110010000",
37063 => "1011110110010011",
37064 => "1011110110010110",
37065 => "1011110110011001",
37066 => "1011110110011100",
37067 => "1011110110011111",
37068 => "1011110110100010",
37069 => "1011110110100101",
37070 => "1011110110101000",
37071 => "1011110110101011",
37072 => "1011110110101110",
37073 => "1011110110110010",
37074 => "1011110110110101",
37075 => "1011110110111000",
37076 => "1011110110111011",
37077 => "1011110110111110",
37078 => "1011110111000001",
37079 => "1011110111000100",
37080 => "1011110111000111",
37081 => "1011110111001010",
37082 => "1011110111001101",
37083 => "1011110111010000",
37084 => "1011110111010011",
37085 => "1011110111010110",
37086 => "1011110111011001",
37087 => "1011110111011101",
37088 => "1011110111100000",
37089 => "1011110111100011",
37090 => "1011110111100110",
37091 => "1011110111101001",
37092 => "1011110111101100",
37093 => "1011110111101111",
37094 => "1011110111110010",
37095 => "1011110111110101",
37096 => "1011110111111000",
37097 => "1011110111111011",
37098 => "1011110111111110",
37099 => "1011111000000001",
37100 => "1011111000000100",
37101 => "1011111000000111",
37102 => "1011111000001010",
37103 => "1011111000001110",
37104 => "1011111000010001",
37105 => "1011111000010100",
37106 => "1011111000010111",
37107 => "1011111000011010",
37108 => "1011111000011101",
37109 => "1011111000100000",
37110 => "1011111000100011",
37111 => "1011111000100110",
37112 => "1011111000101001",
37113 => "1011111000101100",
37114 => "1011111000101111",
37115 => "1011111000110010",
37116 => "1011111000110101",
37117 => "1011111000111000",
37118 => "1011111000111011",
37119 => "1011111000111110",
37120 => "1011111001000001",
37121 => "1011111001000101",
37122 => "1011111001001000",
37123 => "1011111001001011",
37124 => "1011111001001110",
37125 => "1011111001010001",
37126 => "1011111001010100",
37127 => "1011111001010111",
37128 => "1011111001011010",
37129 => "1011111001011101",
37130 => "1011111001100000",
37131 => "1011111001100011",
37132 => "1011111001100110",
37133 => "1011111001101001",
37134 => "1011111001101100",
37135 => "1011111001101111",
37136 => "1011111001110010",
37137 => "1011111001110101",
37138 => "1011111001111000",
37139 => "1011111001111011",
37140 => "1011111001111110",
37141 => "1011111010000010",
37142 => "1011111010000101",
37143 => "1011111010001000",
37144 => "1011111010001011",
37145 => "1011111010001110",
37146 => "1011111010010001",
37147 => "1011111010010100",
37148 => "1011111010010111",
37149 => "1011111010011010",
37150 => "1011111010011101",
37151 => "1011111010100000",
37152 => "1011111010100011",
37153 => "1011111010100110",
37154 => "1011111010101001",
37155 => "1011111010101100",
37156 => "1011111010101111",
37157 => "1011111010110010",
37158 => "1011111010110101",
37159 => "1011111010111000",
37160 => "1011111010111011",
37161 => "1011111010111110",
37162 => "1011111011000001",
37163 => "1011111011000100",
37164 => "1011111011001000",
37165 => "1011111011001011",
37166 => "1011111011001110",
37167 => "1011111011010001",
37168 => "1011111011010100",
37169 => "1011111011010111",
37170 => "1011111011011010",
37171 => "1011111011011101",
37172 => "1011111011100000",
37173 => "1011111011100011",
37174 => "1011111011100110",
37175 => "1011111011101001",
37176 => "1011111011101100",
37177 => "1011111011101111",
37178 => "1011111011110010",
37179 => "1011111011110101",
37180 => "1011111011111000",
37181 => "1011111011111011",
37182 => "1011111011111110",
37183 => "1011111100000001",
37184 => "1011111100000100",
37185 => "1011111100000111",
37186 => "1011111100001010",
37187 => "1011111100001101",
37188 => "1011111100010000",
37189 => "1011111100010011",
37190 => "1011111100010110",
37191 => "1011111100011001",
37192 => "1011111100011100",
37193 => "1011111100011111",
37194 => "1011111100100010",
37195 => "1011111100100101",
37196 => "1011111100101001",
37197 => "1011111100101100",
37198 => "1011111100101111",
37199 => "1011111100110010",
37200 => "1011111100110101",
37201 => "1011111100111000",
37202 => "1011111100111011",
37203 => "1011111100111110",
37204 => "1011111101000001",
37205 => "1011111101000100",
37206 => "1011111101000111",
37207 => "1011111101001010",
37208 => "1011111101001101",
37209 => "1011111101010000",
37210 => "1011111101010011",
37211 => "1011111101010110",
37212 => "1011111101011001",
37213 => "1011111101011100",
37214 => "1011111101011111",
37215 => "1011111101100010",
37216 => "1011111101100101",
37217 => "1011111101101000",
37218 => "1011111101101011",
37219 => "1011111101101110",
37220 => "1011111101110001",
37221 => "1011111101110100",
37222 => "1011111101110111",
37223 => "1011111101111010",
37224 => "1011111101111101",
37225 => "1011111110000000",
37226 => "1011111110000011",
37227 => "1011111110000110",
37228 => "1011111110001001",
37229 => "1011111110001100",
37230 => "1011111110001111",
37231 => "1011111110010010",
37232 => "1011111110010101",
37233 => "1011111110011000",
37234 => "1011111110011011",
37235 => "1011111110011110",
37236 => "1011111110100001",
37237 => "1011111110100100",
37238 => "1011111110100111",
37239 => "1011111110101010",
37240 => "1011111110101101",
37241 => "1011111110110000",
37242 => "1011111110110011",
37243 => "1011111110110110",
37244 => "1011111110111001",
37245 => "1011111110111100",
37246 => "1011111110111111",
37247 => "1011111111000010",
37248 => "1011111111000101",
37249 => "1011111111001000",
37250 => "1011111111001011",
37251 => "1011111111001110",
37252 => "1011111111010001",
37253 => "1011111111010100",
37254 => "1011111111010111",
37255 => "1011111111011010",
37256 => "1011111111011101",
37257 => "1011111111100000",
37258 => "1011111111100011",
37259 => "1011111111100110",
37260 => "1011111111101001",
37261 => "1011111111101100",
37262 => "1011111111101111",
37263 => "1011111111110010",
37264 => "1011111111110101",
37265 => "1011111111111000",
37266 => "1011111111111011",
37267 => "1011111111111110",
37268 => "1100000000000001",
37269 => "1100000000000100",
37270 => "1100000000000111",
37271 => "1100000000001010",
37272 => "1100000000001101",
37273 => "1100000000010000",
37274 => "1100000000010011",
37275 => "1100000000010110",
37276 => "1100000000011001",
37277 => "1100000000011100",
37278 => "1100000000011111",
37279 => "1100000000100010",
37280 => "1100000000100101",
37281 => "1100000000101000",
37282 => "1100000000101011",
37283 => "1100000000101110",
37284 => "1100000000110001",
37285 => "1100000000110100",
37286 => "1100000000110111",
37287 => "1100000000111010",
37288 => "1100000000111101",
37289 => "1100000001000000",
37290 => "1100000001000011",
37291 => "1100000001000110",
37292 => "1100000001001001",
37293 => "1100000001001100",
37294 => "1100000001001111",
37295 => "1100000001010010",
37296 => "1100000001010101",
37297 => "1100000001011000",
37298 => "1100000001011011",
37299 => "1100000001011110",
37300 => "1100000001100001",
37301 => "1100000001100100",
37302 => "1100000001100111",
37303 => "1100000001101010",
37304 => "1100000001101101",
37305 => "1100000001110000",
37306 => "1100000001110011",
37307 => "1100000001110110",
37308 => "1100000001111001",
37309 => "1100000001111100",
37310 => "1100000001111111",
37311 => "1100000010000010",
37312 => "1100000010000101",
37313 => "1100000010001000",
37314 => "1100000010001011",
37315 => "1100000010001110",
37316 => "1100000010010001",
37317 => "1100000010010100",
37318 => "1100000010010111",
37319 => "1100000010011010",
37320 => "1100000010011101",
37321 => "1100000010100000",
37322 => "1100000010100011",
37323 => "1100000010100110",
37324 => "1100000010101001",
37325 => "1100000010101100",
37326 => "1100000010101111",
37327 => "1100000010110010",
37328 => "1100000010110101",
37329 => "1100000010111000",
37330 => "1100000010111011",
37331 => "1100000010111110",
37332 => "1100000011000001",
37333 => "1100000011000100",
37334 => "1100000011000111",
37335 => "1100000011001010",
37336 => "1100000011001101",
37337 => "1100000011010000",
37338 => "1100000011010011",
37339 => "1100000011010110",
37340 => "1100000011011000",
37341 => "1100000011011011",
37342 => "1100000011011110",
37343 => "1100000011100001",
37344 => "1100000011100100",
37345 => "1100000011100111",
37346 => "1100000011101010",
37347 => "1100000011101101",
37348 => "1100000011110000",
37349 => "1100000011110011",
37350 => "1100000011110110",
37351 => "1100000011111001",
37352 => "1100000011111100",
37353 => "1100000011111111",
37354 => "1100000100000010",
37355 => "1100000100000101",
37356 => "1100000100001000",
37357 => "1100000100001011",
37358 => "1100000100001110",
37359 => "1100000100010001",
37360 => "1100000100010100",
37361 => "1100000100010111",
37362 => "1100000100011010",
37363 => "1100000100011101",
37364 => "1100000100100000",
37365 => "1100000100100011",
37366 => "1100000100100110",
37367 => "1100000100101001",
37368 => "1100000100101100",
37369 => "1100000100101111",
37370 => "1100000100110010",
37371 => "1100000100110100",
37372 => "1100000100110111",
37373 => "1100000100111010",
37374 => "1100000100111101",
37375 => "1100000101000000",
37376 => "1100000101000011",
37377 => "1100000101000110",
37378 => "1100000101001001",
37379 => "1100000101001100",
37380 => "1100000101001111",
37381 => "1100000101010010",
37382 => "1100000101010101",
37383 => "1100000101011000",
37384 => "1100000101011011",
37385 => "1100000101011110",
37386 => "1100000101100001",
37387 => "1100000101100100",
37388 => "1100000101100111",
37389 => "1100000101101010",
37390 => "1100000101101101",
37391 => "1100000101110000",
37392 => "1100000101110011",
37393 => "1100000101110110",
37394 => "1100000101111001",
37395 => "1100000101111011",
37396 => "1100000101111110",
37397 => "1100000110000001",
37398 => "1100000110000100",
37399 => "1100000110000111",
37400 => "1100000110001010",
37401 => "1100000110001101",
37402 => "1100000110010000",
37403 => "1100000110010011",
37404 => "1100000110010110",
37405 => "1100000110011001",
37406 => "1100000110011100",
37407 => "1100000110011111",
37408 => "1100000110100010",
37409 => "1100000110100101",
37410 => "1100000110101000",
37411 => "1100000110101011",
37412 => "1100000110101110",
37413 => "1100000110110001",
37414 => "1100000110110100",
37415 => "1100000110110110",
37416 => "1100000110111001",
37417 => "1100000110111100",
37418 => "1100000110111111",
37419 => "1100000111000010",
37420 => "1100000111000101",
37421 => "1100000111001000",
37422 => "1100000111001011",
37423 => "1100000111001110",
37424 => "1100000111010001",
37425 => "1100000111010100",
37426 => "1100000111010111",
37427 => "1100000111011010",
37428 => "1100000111011101",
37429 => "1100000111100000",
37430 => "1100000111100011",
37431 => "1100000111100110",
37432 => "1100000111101000",
37433 => "1100000111101011",
37434 => "1100000111101110",
37435 => "1100000111110001",
37436 => "1100000111110100",
37437 => "1100000111110111",
37438 => "1100000111111010",
37439 => "1100000111111101",
37440 => "1100001000000000",
37441 => "1100001000000011",
37442 => "1100001000000110",
37443 => "1100001000001001",
37444 => "1100001000001100",
37445 => "1100001000001111",
37446 => "1100001000010010",
37447 => "1100001000010101",
37448 => "1100001000010111",
37449 => "1100001000011010",
37450 => "1100001000011101",
37451 => "1100001000100000",
37452 => "1100001000100011",
37453 => "1100001000100110",
37454 => "1100001000101001",
37455 => "1100001000101100",
37456 => "1100001000101111",
37457 => "1100001000110010",
37458 => "1100001000110101",
37459 => "1100001000111000",
37460 => "1100001000111011",
37461 => "1100001000111110",
37462 => "1100001001000001",
37463 => "1100001001000011",
37464 => "1100001001000110",
37465 => "1100001001001001",
37466 => "1100001001001100",
37467 => "1100001001001111",
37468 => "1100001001010010",
37469 => "1100001001010101",
37470 => "1100001001011000",
37471 => "1100001001011011",
37472 => "1100001001011110",
37473 => "1100001001100001",
37474 => "1100001001100100",
37475 => "1100001001100111",
37476 => "1100001001101001",
37477 => "1100001001101100",
37478 => "1100001001101111",
37479 => "1100001001110010",
37480 => "1100001001110101",
37481 => "1100001001111000",
37482 => "1100001001111011",
37483 => "1100001001111110",
37484 => "1100001010000001",
37485 => "1100001010000100",
37486 => "1100001010000111",
37487 => "1100001010001010",
37488 => "1100001010001101",
37489 => "1100001010001111",
37490 => "1100001010010010",
37491 => "1100001010010101",
37492 => "1100001010011000",
37493 => "1100001010011011",
37494 => "1100001010011110",
37495 => "1100001010100001",
37496 => "1100001010100100",
37497 => "1100001010100111",
37498 => "1100001010101010",
37499 => "1100001010101101",
37500 => "1100001010110000",
37501 => "1100001010110010",
37502 => "1100001010110101",
37503 => "1100001010111000",
37504 => "1100001010111011",
37505 => "1100001010111110",
37506 => "1100001011000001",
37507 => "1100001011000100",
37508 => "1100001011000111",
37509 => "1100001011001010",
37510 => "1100001011001101",
37511 => "1100001011010000",
37512 => "1100001011010010",
37513 => "1100001011010101",
37514 => "1100001011011000",
37515 => "1100001011011011",
37516 => "1100001011011110",
37517 => "1100001011100001",
37518 => "1100001011100100",
37519 => "1100001011100111",
37520 => "1100001011101010",
37521 => "1100001011101101",
37522 => "1100001011110000",
37523 => "1100001011110010",
37524 => "1100001011110101",
37525 => "1100001011111000",
37526 => "1100001011111011",
37527 => "1100001011111110",
37528 => "1100001100000001",
37529 => "1100001100000100",
37530 => "1100001100000111",
37531 => "1100001100001010",
37532 => "1100001100001101",
37533 => "1100001100001111",
37534 => "1100001100010010",
37535 => "1100001100010101",
37536 => "1100001100011000",
37537 => "1100001100011011",
37538 => "1100001100011110",
37539 => "1100001100100001",
37540 => "1100001100100100",
37541 => "1100001100100111",
37542 => "1100001100101010",
37543 => "1100001100101100",
37544 => "1100001100101111",
37545 => "1100001100110010",
37546 => "1100001100110101",
37547 => "1100001100111000",
37548 => "1100001100111011",
37549 => "1100001100111110",
37550 => "1100001101000001",
37551 => "1100001101000100",
37552 => "1100001101000111",
37553 => "1100001101001001",
37554 => "1100001101001100",
37555 => "1100001101001111",
37556 => "1100001101010010",
37557 => "1100001101010101",
37558 => "1100001101011000",
37559 => "1100001101011011",
37560 => "1100001101011110",
37561 => "1100001101100001",
37562 => "1100001101100011",
37563 => "1100001101100110",
37564 => "1100001101101001",
37565 => "1100001101101100",
37566 => "1100001101101111",
37567 => "1100001101110010",
37568 => "1100001101110101",
37569 => "1100001101111000",
37570 => "1100001101111011",
37571 => "1100001101111101",
37572 => "1100001110000000",
37573 => "1100001110000011",
37574 => "1100001110000110",
37575 => "1100001110001001",
37576 => "1100001110001100",
37577 => "1100001110001111",
37578 => "1100001110010010",
37579 => "1100001110010101",
37580 => "1100001110010111",
37581 => "1100001110011010",
37582 => "1100001110011101",
37583 => "1100001110100000",
37584 => "1100001110100011",
37585 => "1100001110100110",
37586 => "1100001110101001",
37587 => "1100001110101100",
37588 => "1100001110101111",
37589 => "1100001110110001",
37590 => "1100001110110100",
37591 => "1100001110110111",
37592 => "1100001110111010",
37593 => "1100001110111101",
37594 => "1100001111000000",
37595 => "1100001111000011",
37596 => "1100001111000110",
37597 => "1100001111001000",
37598 => "1100001111001011",
37599 => "1100001111001110",
37600 => "1100001111010001",
37601 => "1100001111010100",
37602 => "1100001111010111",
37603 => "1100001111011010",
37604 => "1100001111011101",
37605 => "1100001111011111",
37606 => "1100001111100010",
37607 => "1100001111100101",
37608 => "1100001111101000",
37609 => "1100001111101011",
37610 => "1100001111101110",
37611 => "1100001111110001",
37612 => "1100001111110100",
37613 => "1100001111110110",
37614 => "1100001111111001",
37615 => "1100001111111100",
37616 => "1100001111111111",
37617 => "1100010000000010",
37618 => "1100010000000101",
37619 => "1100010000001000",
37620 => "1100010000001011",
37621 => "1100010000001101",
37622 => "1100010000010000",
37623 => "1100010000010011",
37624 => "1100010000010110",
37625 => "1100010000011001",
37626 => "1100010000011100",
37627 => "1100010000011111",
37628 => "1100010000100010",
37629 => "1100010000100100",
37630 => "1100010000100111",
37631 => "1100010000101010",
37632 => "1100010000101101",
37633 => "1100010000110000",
37634 => "1100010000110011",
37635 => "1100010000110110",
37636 => "1100010000111000",
37637 => "1100010000111011",
37638 => "1100010000111110",
37639 => "1100010001000001",
37640 => "1100010001000100",
37641 => "1100010001000111",
37642 => "1100010001001010",
37643 => "1100010001001100",
37644 => "1100010001001111",
37645 => "1100010001010010",
37646 => "1100010001010101",
37647 => "1100010001011000",
37648 => "1100010001011011",
37649 => "1100010001011110",
37650 => "1100010001100000",
37651 => "1100010001100011",
37652 => "1100010001100110",
37653 => "1100010001101001",
37654 => "1100010001101100",
37655 => "1100010001101111",
37656 => "1100010001110010",
37657 => "1100010001110100",
37658 => "1100010001110111",
37659 => "1100010001111010",
37660 => "1100010001111101",
37661 => "1100010010000000",
37662 => "1100010010000011",
37663 => "1100010010000110",
37664 => "1100010010001000",
37665 => "1100010010001011",
37666 => "1100010010001110",
37667 => "1100010010010001",
37668 => "1100010010010100",
37669 => "1100010010010111",
37670 => "1100010010011010",
37671 => "1100010010011100",
37672 => "1100010010011111",
37673 => "1100010010100010",
37674 => "1100010010100101",
37675 => "1100010010101000",
37676 => "1100010010101011",
37677 => "1100010010101110",
37678 => "1100010010110000",
37679 => "1100010010110011",
37680 => "1100010010110110",
37681 => "1100010010111001",
37682 => "1100010010111100",
37683 => "1100010010111111",
37684 => "1100010011000001",
37685 => "1100010011000100",
37686 => "1100010011000111",
37687 => "1100010011001010",
37688 => "1100010011001101",
37689 => "1100010011010000",
37690 => "1100010011010011",
37691 => "1100010011010101",
37692 => "1100010011011000",
37693 => "1100010011011011",
37694 => "1100010011011110",
37695 => "1100010011100001",
37696 => "1100010011100100",
37697 => "1100010011100110",
37698 => "1100010011101001",
37699 => "1100010011101100",
37700 => "1100010011101111",
37701 => "1100010011110010",
37702 => "1100010011110101",
37703 => "1100010011110111",
37704 => "1100010011111010",
37705 => "1100010011111101",
37706 => "1100010100000000",
37707 => "1100010100000011",
37708 => "1100010100000110",
37709 => "1100010100001000",
37710 => "1100010100001011",
37711 => "1100010100001110",
37712 => "1100010100010001",
37713 => "1100010100010100",
37714 => "1100010100010111",
37715 => "1100010100011001",
37716 => "1100010100011100",
37717 => "1100010100011111",
37718 => "1100010100100010",
37719 => "1100010100100101",
37720 => "1100010100101000",
37721 => "1100010100101010",
37722 => "1100010100101101",
37723 => "1100010100110000",
37724 => "1100010100110011",
37725 => "1100010100110110",
37726 => "1100010100111001",
37727 => "1100010100111011",
37728 => "1100010100111110",
37729 => "1100010101000001",
37730 => "1100010101000100",
37731 => "1100010101000111",
37732 => "1100010101001010",
37733 => "1100010101001100",
37734 => "1100010101001111",
37735 => "1100010101010010",
37736 => "1100010101010101",
37737 => "1100010101011000",
37738 => "1100010101011011",
37739 => "1100010101011101",
37740 => "1100010101100000",
37741 => "1100010101100011",
37742 => "1100010101100110",
37743 => "1100010101101001",
37744 => "1100010101101100",
37745 => "1100010101101110",
37746 => "1100010101110001",
37747 => "1100010101110100",
37748 => "1100010101110111",
37749 => "1100010101111010",
37750 => "1100010101111100",
37751 => "1100010101111111",
37752 => "1100010110000010",
37753 => "1100010110000101",
37754 => "1100010110001000",
37755 => "1100010110001011",
37756 => "1100010110001101",
37757 => "1100010110010000",
37758 => "1100010110010011",
37759 => "1100010110010110",
37760 => "1100010110011001",
37761 => "1100010110011011",
37762 => "1100010110011110",
37763 => "1100010110100001",
37764 => "1100010110100100",
37765 => "1100010110100111",
37766 => "1100010110101010",
37767 => "1100010110101100",
37768 => "1100010110101111",
37769 => "1100010110110010",
37770 => "1100010110110101",
37771 => "1100010110111000",
37772 => "1100010110111010",
37773 => "1100010110111101",
37774 => "1100010111000000",
37775 => "1100010111000011",
37776 => "1100010111000110",
37777 => "1100010111001001",
37778 => "1100010111001011",
37779 => "1100010111001110",
37780 => "1100010111010001",
37781 => "1100010111010100",
37782 => "1100010111010111",
37783 => "1100010111011001",
37784 => "1100010111011100",
37785 => "1100010111011111",
37786 => "1100010111100010",
37787 => "1100010111100101",
37788 => "1100010111100111",
37789 => "1100010111101010",
37790 => "1100010111101101",
37791 => "1100010111110000",
37792 => "1100010111110011",
37793 => "1100010111110101",
37794 => "1100010111111000",
37795 => "1100010111111011",
37796 => "1100010111111110",
37797 => "1100011000000001",
37798 => "1100011000000011",
37799 => "1100011000000110",
37800 => "1100011000001001",
37801 => "1100011000001100",
37802 => "1100011000001111",
37803 => "1100011000010001",
37804 => "1100011000010100",
37805 => "1100011000010111",
37806 => "1100011000011010",
37807 => "1100011000011101",
37808 => "1100011000011111",
37809 => "1100011000100010",
37810 => "1100011000100101",
37811 => "1100011000101000",
37812 => "1100011000101011",
37813 => "1100011000101101",
37814 => "1100011000110000",
37815 => "1100011000110011",
37816 => "1100011000110110",
37817 => "1100011000111001",
37818 => "1100011000111011",
37819 => "1100011000111110",
37820 => "1100011001000001",
37821 => "1100011001000100",
37822 => "1100011001000111",
37823 => "1100011001001001",
37824 => "1100011001001100",
37825 => "1100011001001111",
37826 => "1100011001010010",
37827 => "1100011001010101",
37828 => "1100011001010111",
37829 => "1100011001011010",
37830 => "1100011001011101",
37831 => "1100011001100000",
37832 => "1100011001100011",
37833 => "1100011001100101",
37834 => "1100011001101000",
37835 => "1100011001101011",
37836 => "1100011001101110",
37837 => "1100011001110000",
37838 => "1100011001110011",
37839 => "1100011001110110",
37840 => "1100011001111001",
37841 => "1100011001111100",
37842 => "1100011001111110",
37843 => "1100011010000001",
37844 => "1100011010000100",
37845 => "1100011010000111",
37846 => "1100011010001010",
37847 => "1100011010001100",
37848 => "1100011010001111",
37849 => "1100011010010010",
37850 => "1100011010010101",
37851 => "1100011010010111",
37852 => "1100011010011010",
37853 => "1100011010011101",
37854 => "1100011010100000",
37855 => "1100011010100011",
37856 => "1100011010100101",
37857 => "1100011010101000",
37858 => "1100011010101011",
37859 => "1100011010101110",
37860 => "1100011010110001",
37861 => "1100011010110011",
37862 => "1100011010110110",
37863 => "1100011010111001",
37864 => "1100011010111100",
37865 => "1100011010111110",
37866 => "1100011011000001",
37867 => "1100011011000100",
37868 => "1100011011000111",
37869 => "1100011011001010",
37870 => "1100011011001100",
37871 => "1100011011001111",
37872 => "1100011011010010",
37873 => "1100011011010101",
37874 => "1100011011010111",
37875 => "1100011011011010",
37876 => "1100011011011101",
37877 => "1100011011100000",
37878 => "1100011011100011",
37879 => "1100011011100101",
37880 => "1100011011101000",
37881 => "1100011011101011",
37882 => "1100011011101110",
37883 => "1100011011110000",
37884 => "1100011011110011",
37885 => "1100011011110110",
37886 => "1100011011111001",
37887 => "1100011011111011",
37888 => "1100011011111110",
37889 => "1100011100000001",
37890 => "1100011100000100",
37891 => "1100011100000111",
37892 => "1100011100001001",
37893 => "1100011100001100",
37894 => "1100011100001111",
37895 => "1100011100010010",
37896 => "1100011100010100",
37897 => "1100011100010111",
37898 => "1100011100011010",
37899 => "1100011100011101",
37900 => "1100011100011111",
37901 => "1100011100100010",
37902 => "1100011100100101",
37903 => "1100011100101000",
37904 => "1100011100101010",
37905 => "1100011100101101",
37906 => "1100011100110000",
37907 => "1100011100110011",
37908 => "1100011100110110",
37909 => "1100011100111000",
37910 => "1100011100111011",
37911 => "1100011100111110",
37912 => "1100011101000001",
37913 => "1100011101000011",
37914 => "1100011101000110",
37915 => "1100011101001001",
37916 => "1100011101001100",
37917 => "1100011101001110",
37918 => "1100011101010001",
37919 => "1100011101010100",
37920 => "1100011101010111",
37921 => "1100011101011001",
37922 => "1100011101011100",
37923 => "1100011101011111",
37924 => "1100011101100010",
37925 => "1100011101100100",
37926 => "1100011101100111",
37927 => "1100011101101010",
37928 => "1100011101101101",
37929 => "1100011101101111",
37930 => "1100011101110010",
37931 => "1100011101110101",
37932 => "1100011101111000",
37933 => "1100011101111010",
37934 => "1100011101111101",
37935 => "1100011110000000",
37936 => "1100011110000011",
37937 => "1100011110000101",
37938 => "1100011110001000",
37939 => "1100011110001011",
37940 => "1100011110001110",
37941 => "1100011110010000",
37942 => "1100011110010011",
37943 => "1100011110010110",
37944 => "1100011110011001",
37945 => "1100011110011011",
37946 => "1100011110011110",
37947 => "1100011110100001",
37948 => "1100011110100100",
37949 => "1100011110100110",
37950 => "1100011110101001",
37951 => "1100011110101100",
37952 => "1100011110101111",
37953 => "1100011110110001",
37954 => "1100011110110100",
37955 => "1100011110110111",
37956 => "1100011110111010",
37957 => "1100011110111100",
37958 => "1100011110111111",
37959 => "1100011111000010",
37960 => "1100011111000101",
37961 => "1100011111000111",
37962 => "1100011111001010",
37963 => "1100011111001101",
37964 => "1100011111010000",
37965 => "1100011111010010",
37966 => "1100011111010101",
37967 => "1100011111011000",
37968 => "1100011111011011",
37969 => "1100011111011101",
37970 => "1100011111100000",
37971 => "1100011111100011",
37972 => "1100011111100110",
37973 => "1100011111101000",
37974 => "1100011111101011",
37975 => "1100011111101110",
37976 => "1100011111110000",
37977 => "1100011111110011",
37978 => "1100011111110110",
37979 => "1100011111111001",
37980 => "1100011111111011",
37981 => "1100011111111110",
37982 => "1100100000000001",
37983 => "1100100000000100",
37984 => "1100100000000110",
37985 => "1100100000001001",
37986 => "1100100000001100",
37987 => "1100100000001111",
37988 => "1100100000010001",
37989 => "1100100000010100",
37990 => "1100100000010111",
37991 => "1100100000011001",
37992 => "1100100000011100",
37993 => "1100100000011111",
37994 => "1100100000100010",
37995 => "1100100000100100",
37996 => "1100100000100111",
37997 => "1100100000101010",
37998 => "1100100000101101",
37999 => "1100100000101111",
38000 => "1100100000110010",
38001 => "1100100000110101",
38002 => "1100100000111000",
38003 => "1100100000111010",
38004 => "1100100000111101",
38005 => "1100100001000000",
38006 => "1100100001000010",
38007 => "1100100001000101",
38008 => "1100100001001000",
38009 => "1100100001001011",
38010 => "1100100001001101",
38011 => "1100100001010000",
38012 => "1100100001010011",
38013 => "1100100001010101",
38014 => "1100100001011000",
38015 => "1100100001011011",
38016 => "1100100001011110",
38017 => "1100100001100000",
38018 => "1100100001100011",
38019 => "1100100001100110",
38020 => "1100100001101001",
38021 => "1100100001101011",
38022 => "1100100001101110",
38023 => "1100100001110001",
38024 => "1100100001110011",
38025 => "1100100001110110",
38026 => "1100100001111001",
38027 => "1100100001111100",
38028 => "1100100001111110",
38029 => "1100100010000001",
38030 => "1100100010000100",
38031 => "1100100010000110",
38032 => "1100100010001001",
38033 => "1100100010001100",
38034 => "1100100010001111",
38035 => "1100100010010001",
38036 => "1100100010010100",
38037 => "1100100010010111",
38038 => "1100100010011001",
38039 => "1100100010011100",
38040 => "1100100010011111",
38041 => "1100100010100010",
38042 => "1100100010100100",
38043 => "1100100010100111",
38044 => "1100100010101010",
38045 => "1100100010101100",
38046 => "1100100010101111",
38047 => "1100100010110010",
38048 => "1100100010110101",
38049 => "1100100010110111",
38050 => "1100100010111010",
38051 => "1100100010111101",
38052 => "1100100010111111",
38053 => "1100100011000010",
38054 => "1100100011000101",
38055 => "1100100011000111",
38056 => "1100100011001010",
38057 => "1100100011001101",
38058 => "1100100011010000",
38059 => "1100100011010010",
38060 => "1100100011010101",
38061 => "1100100011011000",
38062 => "1100100011011010",
38063 => "1100100011011101",
38064 => "1100100011100000",
38065 => "1100100011100011",
38066 => "1100100011100101",
38067 => "1100100011101000",
38068 => "1100100011101011",
38069 => "1100100011101101",
38070 => "1100100011110000",
38071 => "1100100011110011",
38072 => "1100100011110101",
38073 => "1100100011111000",
38074 => "1100100011111011",
38075 => "1100100011111110",
38076 => "1100100100000000",
38077 => "1100100100000011",
38078 => "1100100100000110",
38079 => "1100100100001000",
38080 => "1100100100001011",
38081 => "1100100100001110",
38082 => "1100100100010000",
38083 => "1100100100010011",
38084 => "1100100100010110",
38085 => "1100100100011001",
38086 => "1100100100011011",
38087 => "1100100100011110",
38088 => "1100100100100001",
38089 => "1100100100100011",
38090 => "1100100100100110",
38091 => "1100100100101001",
38092 => "1100100100101011",
38093 => "1100100100101110",
38094 => "1100100100110001",
38095 => "1100100100110011",
38096 => "1100100100110110",
38097 => "1100100100111001",
38098 => "1100100100111100",
38099 => "1100100100111110",
38100 => "1100100101000001",
38101 => "1100100101000100",
38102 => "1100100101000110",
38103 => "1100100101001001",
38104 => "1100100101001100",
38105 => "1100100101001110",
38106 => "1100100101010001",
38107 => "1100100101010100",
38108 => "1100100101010110",
38109 => "1100100101011001",
38110 => "1100100101011100",
38111 => "1100100101011110",
38112 => "1100100101100001",
38113 => "1100100101100100",
38114 => "1100100101100111",
38115 => "1100100101101001",
38116 => "1100100101101100",
38117 => "1100100101101111",
38118 => "1100100101110001",
38119 => "1100100101110100",
38120 => "1100100101110111",
38121 => "1100100101111001",
38122 => "1100100101111100",
38123 => "1100100101111111",
38124 => "1100100110000001",
38125 => "1100100110000100",
38126 => "1100100110000111",
38127 => "1100100110001001",
38128 => "1100100110001100",
38129 => "1100100110001111",
38130 => "1100100110010001",
38131 => "1100100110010100",
38132 => "1100100110010111",
38133 => "1100100110011001",
38134 => "1100100110011100",
38135 => "1100100110011111",
38136 => "1100100110100010",
38137 => "1100100110100100",
38138 => "1100100110100111",
38139 => "1100100110101010",
38140 => "1100100110101100",
38141 => "1100100110101111",
38142 => "1100100110110010",
38143 => "1100100110110100",
38144 => "1100100110110111",
38145 => "1100100110111010",
38146 => "1100100110111100",
38147 => "1100100110111111",
38148 => "1100100111000010",
38149 => "1100100111000100",
38150 => "1100100111000111",
38151 => "1100100111001010",
38152 => "1100100111001100",
38153 => "1100100111001111",
38154 => "1100100111010010",
38155 => "1100100111010100",
38156 => "1100100111010111",
38157 => "1100100111011010",
38158 => "1100100111011100",
38159 => "1100100111011111",
38160 => "1100100111100010",
38161 => "1100100111100100",
38162 => "1100100111100111",
38163 => "1100100111101010",
38164 => "1100100111101100",
38165 => "1100100111101111",
38166 => "1100100111110010",
38167 => "1100100111110100",
38168 => "1100100111110111",
38169 => "1100100111111010",
38170 => "1100100111111100",
38171 => "1100100111111111",
38172 => "1100101000000010",
38173 => "1100101000000100",
38174 => "1100101000000111",
38175 => "1100101000001010",
38176 => "1100101000001100",
38177 => "1100101000001111",
38178 => "1100101000010010",
38179 => "1100101000010100",
38180 => "1100101000010111",
38181 => "1100101000011010",
38182 => "1100101000011100",
38183 => "1100101000011111",
38184 => "1100101000100010",
38185 => "1100101000100100",
38186 => "1100101000100111",
38187 => "1100101000101010",
38188 => "1100101000101100",
38189 => "1100101000101111",
38190 => "1100101000110001",
38191 => "1100101000110100",
38192 => "1100101000110111",
38193 => "1100101000111001",
38194 => "1100101000111100",
38195 => "1100101000111111",
38196 => "1100101001000001",
38197 => "1100101001000100",
38198 => "1100101001000111",
38199 => "1100101001001001",
38200 => "1100101001001100",
38201 => "1100101001001111",
38202 => "1100101001010001",
38203 => "1100101001010100",
38204 => "1100101001010111",
38205 => "1100101001011001",
38206 => "1100101001011100",
38207 => "1100101001011111",
38208 => "1100101001100001",
38209 => "1100101001100100",
38210 => "1100101001100111",
38211 => "1100101001101001",
38212 => "1100101001101100",
38213 => "1100101001101110",
38214 => "1100101001110001",
38215 => "1100101001110100",
38216 => "1100101001110110",
38217 => "1100101001111001",
38218 => "1100101001111100",
38219 => "1100101001111110",
38220 => "1100101010000001",
38221 => "1100101010000100",
38222 => "1100101010000110",
38223 => "1100101010001001",
38224 => "1100101010001100",
38225 => "1100101010001110",
38226 => "1100101010010001",
38227 => "1100101010010100",
38228 => "1100101010010110",
38229 => "1100101010011001",
38230 => "1100101010011011",
38231 => "1100101010011110",
38232 => "1100101010100001",
38233 => "1100101010100011",
38234 => "1100101010100110",
38235 => "1100101010101001",
38236 => "1100101010101011",
38237 => "1100101010101110",
38238 => "1100101010110001",
38239 => "1100101010110011",
38240 => "1100101010110110",
38241 => "1100101010111000",
38242 => "1100101010111011",
38243 => "1100101010111110",
38244 => "1100101011000000",
38245 => "1100101011000011",
38246 => "1100101011000110",
38247 => "1100101011001000",
38248 => "1100101011001011",
38249 => "1100101011001110",
38250 => "1100101011010000",
38251 => "1100101011010011",
38252 => "1100101011010101",
38253 => "1100101011011000",
38254 => "1100101011011011",
38255 => "1100101011011101",
38256 => "1100101011100000",
38257 => "1100101011100011",
38258 => "1100101011100101",
38259 => "1100101011101000",
38260 => "1100101011101010",
38261 => "1100101011101101",
38262 => "1100101011110000",
38263 => "1100101011110010",
38264 => "1100101011110101",
38265 => "1100101011111000",
38266 => "1100101011111010",
38267 => "1100101011111101",
38268 => "1100101100000000",
38269 => "1100101100000010",
38270 => "1100101100000101",
38271 => "1100101100000111",
38272 => "1100101100001010",
38273 => "1100101100001101",
38274 => "1100101100001111",
38275 => "1100101100010010",
38276 => "1100101100010101",
38277 => "1100101100010111",
38278 => "1100101100011010",
38279 => "1100101100011100",
38280 => "1100101100011111",
38281 => "1100101100100010",
38282 => "1100101100100100",
38283 => "1100101100100111",
38284 => "1100101100101010",
38285 => "1100101100101100",
38286 => "1100101100101111",
38287 => "1100101100110001",
38288 => "1100101100110100",
38289 => "1100101100110111",
38290 => "1100101100111001",
38291 => "1100101100111100",
38292 => "1100101100111110",
38293 => "1100101101000001",
38294 => "1100101101000100",
38295 => "1100101101000110",
38296 => "1100101101001001",
38297 => "1100101101001100",
38298 => "1100101101001110",
38299 => "1100101101010001",
38300 => "1100101101010011",
38301 => "1100101101010110",
38302 => "1100101101011001",
38303 => "1100101101011011",
38304 => "1100101101011110",
38305 => "1100101101100000",
38306 => "1100101101100011",
38307 => "1100101101100110",
38308 => "1100101101101000",
38309 => "1100101101101011",
38310 => "1100101101101110",
38311 => "1100101101110000",
38312 => "1100101101110011",
38313 => "1100101101110101",
38314 => "1100101101111000",
38315 => "1100101101111011",
38316 => "1100101101111101",
38317 => "1100101110000000",
38318 => "1100101110000010",
38319 => "1100101110000101",
38320 => "1100101110001000",
38321 => "1100101110001010",
38322 => "1100101110001101",
38323 => "1100101110001111",
38324 => "1100101110010010",
38325 => "1100101110010101",
38326 => "1100101110010111",
38327 => "1100101110011010",
38328 => "1100101110011100",
38329 => "1100101110011111",
38330 => "1100101110100010",
38331 => "1100101110100100",
38332 => "1100101110100111",
38333 => "1100101110101001",
38334 => "1100101110101100",
38335 => "1100101110101111",
38336 => "1100101110110001",
38337 => "1100101110110100",
38338 => "1100101110110110",
38339 => "1100101110111001",
38340 => "1100101110111100",
38341 => "1100101110111110",
38342 => "1100101111000001",
38343 => "1100101111000011",
38344 => "1100101111000110",
38345 => "1100101111001001",
38346 => "1100101111001011",
38347 => "1100101111001110",
38348 => "1100101111010000",
38349 => "1100101111010011",
38350 => "1100101111010110",
38351 => "1100101111011000",
38352 => "1100101111011011",
38353 => "1100101111011101",
38354 => "1100101111100000",
38355 => "1100101111100011",
38356 => "1100101111100101",
38357 => "1100101111101000",
38358 => "1100101111101010",
38359 => "1100101111101101",
38360 => "1100101111110000",
38361 => "1100101111110010",
38362 => "1100101111110101",
38363 => "1100101111110111",
38364 => "1100101111111010",
38365 => "1100101111111101",
38366 => "1100101111111111",
38367 => "1100110000000010",
38368 => "1100110000000100",
38369 => "1100110000000111",
38370 => "1100110000001001",
38371 => "1100110000001100",
38372 => "1100110000001111",
38373 => "1100110000010001",
38374 => "1100110000010100",
38375 => "1100110000010110",
38376 => "1100110000011001",
38377 => "1100110000011100",
38378 => "1100110000011110",
38379 => "1100110000100001",
38380 => "1100110000100011",
38381 => "1100110000100110",
38382 => "1100110000101001",
38383 => "1100110000101011",
38384 => "1100110000101110",
38385 => "1100110000110000",
38386 => "1100110000110011",
38387 => "1100110000110101",
38388 => "1100110000111000",
38389 => "1100110000111011",
38390 => "1100110000111101",
38391 => "1100110001000000",
38392 => "1100110001000010",
38393 => "1100110001000101",
38394 => "1100110001001000",
38395 => "1100110001001010",
38396 => "1100110001001101",
38397 => "1100110001001111",
38398 => "1100110001010010",
38399 => "1100110001010100",
38400 => "1100110001010111",
38401 => "1100110001011010",
38402 => "1100110001011100",
38403 => "1100110001011111",
38404 => "1100110001100001",
38405 => "1100110001100100",
38406 => "1100110001100110",
38407 => "1100110001101001",
38408 => "1100110001101100",
38409 => "1100110001101110",
38410 => "1100110001110001",
38411 => "1100110001110011",
38412 => "1100110001110110",
38413 => "1100110001111000",
38414 => "1100110001111011",
38415 => "1100110001111110",
38416 => "1100110010000000",
38417 => "1100110010000011",
38418 => "1100110010000101",
38419 => "1100110010001000",
38420 => "1100110010001010",
38421 => "1100110010001101",
38422 => "1100110010010000",
38423 => "1100110010010010",
38424 => "1100110010010101",
38425 => "1100110010010111",
38426 => "1100110010011010",
38427 => "1100110010011100",
38428 => "1100110010011111",
38429 => "1100110010100010",
38430 => "1100110010100100",
38431 => "1100110010100111",
38432 => "1100110010101001",
38433 => "1100110010101100",
38434 => "1100110010101110",
38435 => "1100110010110001",
38436 => "1100110010110100",
38437 => "1100110010110110",
38438 => "1100110010111001",
38439 => "1100110010111011",
38440 => "1100110010111110",
38441 => "1100110011000000",
38442 => "1100110011000011",
38443 => "1100110011000101",
38444 => "1100110011001000",
38445 => "1100110011001011",
38446 => "1100110011001101",
38447 => "1100110011010000",
38448 => "1100110011010010",
38449 => "1100110011010101",
38450 => "1100110011010111",
38451 => "1100110011011010",
38452 => "1100110011011100",
38453 => "1100110011011111",
38454 => "1100110011100010",
38455 => "1100110011100100",
38456 => "1100110011100111",
38457 => "1100110011101001",
38458 => "1100110011101100",
38459 => "1100110011101110",
38460 => "1100110011110001",
38461 => "1100110011110011",
38462 => "1100110011110110",
38463 => "1100110011111001",
38464 => "1100110011111011",
38465 => "1100110011111110",
38466 => "1100110100000000",
38467 => "1100110100000011",
38468 => "1100110100000101",
38469 => "1100110100001000",
38470 => "1100110100001010",
38471 => "1100110100001101",
38472 => "1100110100010000",
38473 => "1100110100010010",
38474 => "1100110100010101",
38475 => "1100110100010111",
38476 => "1100110100011010",
38477 => "1100110100011100",
38478 => "1100110100011111",
38479 => "1100110100100001",
38480 => "1100110100100100",
38481 => "1100110100100110",
38482 => "1100110100101001",
38483 => "1100110100101100",
38484 => "1100110100101110",
38485 => "1100110100110001",
38486 => "1100110100110011",
38487 => "1100110100110110",
38488 => "1100110100111000",
38489 => "1100110100111011",
38490 => "1100110100111101",
38491 => "1100110101000000",
38492 => "1100110101000010",
38493 => "1100110101000101",
38494 => "1100110101001000",
38495 => "1100110101001010",
38496 => "1100110101001101",
38497 => "1100110101001111",
38498 => "1100110101010010",
38499 => "1100110101010100",
38500 => "1100110101010111",
38501 => "1100110101011001",
38502 => "1100110101011100",
38503 => "1100110101011110",
38504 => "1100110101100001",
38505 => "1100110101100100",
38506 => "1100110101100110",
38507 => "1100110101101001",
38508 => "1100110101101011",
38509 => "1100110101101110",
38510 => "1100110101110000",
38511 => "1100110101110011",
38512 => "1100110101110101",
38513 => "1100110101111000",
38514 => "1100110101111010",
38515 => "1100110101111101",
38516 => "1100110101111111",
38517 => "1100110110000010",
38518 => "1100110110000100",
38519 => "1100110110000111",
38520 => "1100110110001010",
38521 => "1100110110001100",
38522 => "1100110110001111",
38523 => "1100110110010001",
38524 => "1100110110010100",
38525 => "1100110110010110",
38526 => "1100110110011001",
38527 => "1100110110011011",
38528 => "1100110110011110",
38529 => "1100110110100000",
38530 => "1100110110100011",
38531 => "1100110110100101",
38532 => "1100110110101000",
38533 => "1100110110101010",
38534 => "1100110110101101",
38535 => "1100110110101111",
38536 => "1100110110110010",
38537 => "1100110110110101",
38538 => "1100110110110111",
38539 => "1100110110111010",
38540 => "1100110110111100",
38541 => "1100110110111111",
38542 => "1100110111000001",
38543 => "1100110111000100",
38544 => "1100110111000110",
38545 => "1100110111001001",
38546 => "1100110111001011",
38547 => "1100110111001110",
38548 => "1100110111010000",
38549 => "1100110111010011",
38550 => "1100110111010101",
38551 => "1100110111011000",
38552 => "1100110111011010",
38553 => "1100110111011101",
38554 => "1100110111011111",
38555 => "1100110111100010",
38556 => "1100110111100100",
38557 => "1100110111100111",
38558 => "1100110111101001",
38559 => "1100110111101100",
38560 => "1100110111101111",
38561 => "1100110111110001",
38562 => "1100110111110100",
38563 => "1100110111110110",
38564 => "1100110111111001",
38565 => "1100110111111011",
38566 => "1100110111111110",
38567 => "1100111000000000",
38568 => "1100111000000011",
38569 => "1100111000000101",
38570 => "1100111000001000",
38571 => "1100111000001010",
38572 => "1100111000001101",
38573 => "1100111000001111",
38574 => "1100111000010010",
38575 => "1100111000010100",
38576 => "1100111000010111",
38577 => "1100111000011001",
38578 => "1100111000011100",
38579 => "1100111000011110",
38580 => "1100111000100001",
38581 => "1100111000100011",
38582 => "1100111000100110",
38583 => "1100111000101000",
38584 => "1100111000101011",
38585 => "1100111000101101",
38586 => "1100111000110000",
38587 => "1100111000110010",
38588 => "1100111000110101",
38589 => "1100111000110111",
38590 => "1100111000111010",
38591 => "1100111000111100",
38592 => "1100111000111111",
38593 => "1100111001000001",
38594 => "1100111001000100",
38595 => "1100111001000110",
38596 => "1100111001001001",
38597 => "1100111001001011",
38598 => "1100111001001110",
38599 => "1100111001010000",
38600 => "1100111001010011",
38601 => "1100111001010101",
38602 => "1100111001011000",
38603 => "1100111001011010",
38604 => "1100111001011101",
38605 => "1100111001011111",
38606 => "1100111001100010",
38607 => "1100111001100100",
38608 => "1100111001100111",
38609 => "1100111001101001",
38610 => "1100111001101100",
38611 => "1100111001101110",
38612 => "1100111001110001",
38613 => "1100111001110011",
38614 => "1100111001110110",
38615 => "1100111001111000",
38616 => "1100111001111011",
38617 => "1100111001111101",
38618 => "1100111010000000",
38619 => "1100111010000010",
38620 => "1100111010000101",
38621 => "1100111010000111",
38622 => "1100111010001010",
38623 => "1100111010001100",
38624 => "1100111010001111",
38625 => "1100111010010001",
38626 => "1100111010010100",
38627 => "1100111010010110",
38628 => "1100111010011001",
38629 => "1100111010011011",
38630 => "1100111010011110",
38631 => "1100111010100000",
38632 => "1100111010100011",
38633 => "1100111010100101",
38634 => "1100111010101000",
38635 => "1100111010101010",
38636 => "1100111010101101",
38637 => "1100111010101111",
38638 => "1100111010110010",
38639 => "1100111010110100",
38640 => "1100111010110111",
38641 => "1100111010111001",
38642 => "1100111010111100",
38643 => "1100111010111110",
38644 => "1100111011000001",
38645 => "1100111011000011",
38646 => "1100111011000110",
38647 => "1100111011001000",
38648 => "1100111011001011",
38649 => "1100111011001101",
38650 => "1100111011010000",
38651 => "1100111011010010",
38652 => "1100111011010101",
38653 => "1100111011010111",
38654 => "1100111011011001",
38655 => "1100111011011100",
38656 => "1100111011011110",
38657 => "1100111011100001",
38658 => "1100111011100011",
38659 => "1100111011100110",
38660 => "1100111011101000",
38661 => "1100111011101011",
38662 => "1100111011101101",
38663 => "1100111011110000",
38664 => "1100111011110010",
38665 => "1100111011110101",
38666 => "1100111011110111",
38667 => "1100111011111010",
38668 => "1100111011111100",
38669 => "1100111011111111",
38670 => "1100111100000001",
38671 => "1100111100000100",
38672 => "1100111100000110",
38673 => "1100111100001001",
38674 => "1100111100001011",
38675 => "1100111100001110",
38676 => "1100111100010000",
38677 => "1100111100010010",
38678 => "1100111100010101",
38679 => "1100111100010111",
38680 => "1100111100011010",
38681 => "1100111100011100",
38682 => "1100111100011111",
38683 => "1100111100100001",
38684 => "1100111100100100",
38685 => "1100111100100110",
38686 => "1100111100101001",
38687 => "1100111100101011",
38688 => "1100111100101110",
38689 => "1100111100110000",
38690 => "1100111100110011",
38691 => "1100111100110101",
38692 => "1100111100111000",
38693 => "1100111100111010",
38694 => "1100111100111100",
38695 => "1100111100111111",
38696 => "1100111101000001",
38697 => "1100111101000100",
38698 => "1100111101000110",
38699 => "1100111101001001",
38700 => "1100111101001011",
38701 => "1100111101001110",
38702 => "1100111101010000",
38703 => "1100111101010011",
38704 => "1100111101010101",
38705 => "1100111101011000",
38706 => "1100111101011010",
38707 => "1100111101011101",
38708 => "1100111101011111",
38709 => "1100111101100001",
38710 => "1100111101100100",
38711 => "1100111101100110",
38712 => "1100111101101001",
38713 => "1100111101101011",
38714 => "1100111101101110",
38715 => "1100111101110000",
38716 => "1100111101110011",
38717 => "1100111101110101",
38718 => "1100111101111000",
38719 => "1100111101111010",
38720 => "1100111101111100",
38721 => "1100111101111111",
38722 => "1100111110000001",
38723 => "1100111110000100",
38724 => "1100111110000110",
38725 => "1100111110001001",
38726 => "1100111110001011",
38727 => "1100111110001110",
38728 => "1100111110010000",
38729 => "1100111110010011",
38730 => "1100111110010101",
38731 => "1100111110011000",
38732 => "1100111110011010",
38733 => "1100111110011100",
38734 => "1100111110011111",
38735 => "1100111110100001",
38736 => "1100111110100100",
38737 => "1100111110100110",
38738 => "1100111110101001",
38739 => "1100111110101011",
38740 => "1100111110101110",
38741 => "1100111110110000",
38742 => "1100111110110010",
38743 => "1100111110110101",
38744 => "1100111110110111",
38745 => "1100111110111010",
38746 => "1100111110111100",
38747 => "1100111110111111",
38748 => "1100111111000001",
38749 => "1100111111000100",
38750 => "1100111111000110",
38751 => "1100111111001001",
38752 => "1100111111001011",
38753 => "1100111111001101",
38754 => "1100111111010000",
38755 => "1100111111010010",
38756 => "1100111111010101",
38757 => "1100111111010111",
38758 => "1100111111011010",
38759 => "1100111111011100",
38760 => "1100111111011110",
38761 => "1100111111100001",
38762 => "1100111111100011",
38763 => "1100111111100110",
38764 => "1100111111101000",
38765 => "1100111111101011",
38766 => "1100111111101101",
38767 => "1100111111110000",
38768 => "1100111111110010",
38769 => "1100111111110100",
38770 => "1100111111110111",
38771 => "1100111111111001",
38772 => "1100111111111100",
38773 => "1100111111111110",
38774 => "1101000000000001",
38775 => "1101000000000011",
38776 => "1101000000000110",
38777 => "1101000000001000",
38778 => "1101000000001010",
38779 => "1101000000001101",
38780 => "1101000000001111",
38781 => "1101000000010010",
38782 => "1101000000010100",
38783 => "1101000000010111",
38784 => "1101000000011001",
38785 => "1101000000011011",
38786 => "1101000000011110",
38787 => "1101000000100000",
38788 => "1101000000100011",
38789 => "1101000000100101",
38790 => "1101000000101000",
38791 => "1101000000101010",
38792 => "1101000000101100",
38793 => "1101000000101111",
38794 => "1101000000110001",
38795 => "1101000000110100",
38796 => "1101000000110110",
38797 => "1101000000111001",
38798 => "1101000000111011",
38799 => "1101000000111101",
38800 => "1101000001000000",
38801 => "1101000001000010",
38802 => "1101000001000101",
38803 => "1101000001000111",
38804 => "1101000001001010",
38805 => "1101000001001100",
38806 => "1101000001001110",
38807 => "1101000001010001",
38808 => "1101000001010011",
38809 => "1101000001010110",
38810 => "1101000001011000",
38811 => "1101000001011011",
38812 => "1101000001011101",
38813 => "1101000001011111",
38814 => "1101000001100010",
38815 => "1101000001100100",
38816 => "1101000001100111",
38817 => "1101000001101001",
38818 => "1101000001101100",
38819 => "1101000001101110",
38820 => "1101000001110000",
38821 => "1101000001110011",
38822 => "1101000001110101",
38823 => "1101000001111000",
38824 => "1101000001111010",
38825 => "1101000001111100",
38826 => "1101000001111111",
38827 => "1101000010000001",
38828 => "1101000010000100",
38829 => "1101000010000110",
38830 => "1101000010001001",
38831 => "1101000010001011",
38832 => "1101000010001101",
38833 => "1101000010010000",
38834 => "1101000010010010",
38835 => "1101000010010101",
38836 => "1101000010010111",
38837 => "1101000010011001",
38838 => "1101000010011100",
38839 => "1101000010011110",
38840 => "1101000010100001",
38841 => "1101000010100011",
38842 => "1101000010100110",
38843 => "1101000010101000",
38844 => "1101000010101010",
38845 => "1101000010101101",
38846 => "1101000010101111",
38847 => "1101000010110010",
38848 => "1101000010110100",
38849 => "1101000010110110",
38850 => "1101000010111001",
38851 => "1101000010111011",
38852 => "1101000010111110",
38853 => "1101000011000000",
38854 => "1101000011000010",
38855 => "1101000011000101",
38856 => "1101000011000111",
38857 => "1101000011001010",
38858 => "1101000011001100",
38859 => "1101000011001110",
38860 => "1101000011010001",
38861 => "1101000011010011",
38862 => "1101000011010110",
38863 => "1101000011011000",
38864 => "1101000011011011",
38865 => "1101000011011101",
38866 => "1101000011011111",
38867 => "1101000011100010",
38868 => "1101000011100100",
38869 => "1101000011100111",
38870 => "1101000011101001",
38871 => "1101000011101011",
38872 => "1101000011101110",
38873 => "1101000011110000",
38874 => "1101000011110011",
38875 => "1101000011110101",
38876 => "1101000011110111",
38877 => "1101000011111010",
38878 => "1101000011111100",
38879 => "1101000011111111",
38880 => "1101000100000001",
38881 => "1101000100000011",
38882 => "1101000100000110",
38883 => "1101000100001000",
38884 => "1101000100001011",
38885 => "1101000100001101",
38886 => "1101000100001111",
38887 => "1101000100010010",
38888 => "1101000100010100",
38889 => "1101000100010110",
38890 => "1101000100011001",
38891 => "1101000100011011",
38892 => "1101000100011110",
38893 => "1101000100100000",
38894 => "1101000100100010",
38895 => "1101000100100101",
38896 => "1101000100100111",
38897 => "1101000100101010",
38898 => "1101000100101100",
38899 => "1101000100101110",
38900 => "1101000100110001",
38901 => "1101000100110011",
38902 => "1101000100110110",
38903 => "1101000100111000",
38904 => "1101000100111010",
38905 => "1101000100111101",
38906 => "1101000100111111",
38907 => "1101000101000010",
38908 => "1101000101000100",
38909 => "1101000101000110",
38910 => "1101000101001001",
38911 => "1101000101001011",
38912 => "1101000101001101",
38913 => "1101000101010000",
38914 => "1101000101010010",
38915 => "1101000101010101",
38916 => "1101000101010111",
38917 => "1101000101011001",
38918 => "1101000101011100",
38919 => "1101000101011110",
38920 => "1101000101100001",
38921 => "1101000101100011",
38922 => "1101000101100101",
38923 => "1101000101101000",
38924 => "1101000101101010",
38925 => "1101000101101100",
38926 => "1101000101101111",
38927 => "1101000101110001",
38928 => "1101000101110100",
38929 => "1101000101110110",
38930 => "1101000101111000",
38931 => "1101000101111011",
38932 => "1101000101111101",
38933 => "1101000110000000",
38934 => "1101000110000010",
38935 => "1101000110000100",
38936 => "1101000110000111",
38937 => "1101000110001001",
38938 => "1101000110001011",
38939 => "1101000110001110",
38940 => "1101000110010000",
38941 => "1101000110010011",
38942 => "1101000110010101",
38943 => "1101000110010111",
38944 => "1101000110011010",
38945 => "1101000110011100",
38946 => "1101000110011110",
38947 => "1101000110100001",
38948 => "1101000110100011",
38949 => "1101000110100110",
38950 => "1101000110101000",
38951 => "1101000110101010",
38952 => "1101000110101101",
38953 => "1101000110101111",
38954 => "1101000110110001",
38955 => "1101000110110100",
38956 => "1101000110110110",
38957 => "1101000110111000",
38958 => "1101000110111011",
38959 => "1101000110111101",
38960 => "1101000111000000",
38961 => "1101000111000010",
38962 => "1101000111000100",
38963 => "1101000111000111",
38964 => "1101000111001001",
38965 => "1101000111001011",
38966 => "1101000111001110",
38967 => "1101000111010000",
38968 => "1101000111010011",
38969 => "1101000111010101",
38970 => "1101000111010111",
38971 => "1101000111011010",
38972 => "1101000111011100",
38973 => "1101000111011110",
38974 => "1101000111100001",
38975 => "1101000111100011",
38976 => "1101000111100101",
38977 => "1101000111101000",
38978 => "1101000111101010",
38979 => "1101000111101101",
38980 => "1101000111101111",
38981 => "1101000111110001",
38982 => "1101000111110100",
38983 => "1101000111110110",
38984 => "1101000111111000",
38985 => "1101000111111011",
38986 => "1101000111111101",
38987 => "1101000111111111",
38988 => "1101001000000010",
38989 => "1101001000000100",
38990 => "1101001000000110",
38991 => "1101001000001001",
38992 => "1101001000001011",
38993 => "1101001000001110",
38994 => "1101001000010000",
38995 => "1101001000010010",
38996 => "1101001000010101",
38997 => "1101001000010111",
38998 => "1101001000011001",
38999 => "1101001000011100",
39000 => "1101001000011110",
39001 => "1101001000100000",
39002 => "1101001000100011",
39003 => "1101001000100101",
39004 => "1101001000100111",
39005 => "1101001000101010",
39006 => "1101001000101100",
39007 => "1101001000101110",
39008 => "1101001000110001",
39009 => "1101001000110011",
39010 => "1101001000110110",
39011 => "1101001000111000",
39012 => "1101001000111010",
39013 => "1101001000111101",
39014 => "1101001000111111",
39015 => "1101001001000001",
39016 => "1101001001000100",
39017 => "1101001001000110",
39018 => "1101001001001000",
39019 => "1101001001001011",
39020 => "1101001001001101",
39021 => "1101001001001111",
39022 => "1101001001010010",
39023 => "1101001001010100",
39024 => "1101001001010110",
39025 => "1101001001011001",
39026 => "1101001001011011",
39027 => "1101001001011101",
39028 => "1101001001100000",
39029 => "1101001001100010",
39030 => "1101001001100100",
39031 => "1101001001100111",
39032 => "1101001001101001",
39033 => "1101001001101011",
39034 => "1101001001101110",
39035 => "1101001001110000",
39036 => "1101001001110011",
39037 => "1101001001110101",
39038 => "1101001001110111",
39039 => "1101001001111010",
39040 => "1101001001111100",
39041 => "1101001001111110",
39042 => "1101001010000001",
39043 => "1101001010000011",
39044 => "1101001010000101",
39045 => "1101001010001000",
39046 => "1101001010001010",
39047 => "1101001010001100",
39048 => "1101001010001111",
39049 => "1101001010010001",
39050 => "1101001010010011",
39051 => "1101001010010110",
39052 => "1101001010011000",
39053 => "1101001010011010",
39054 => "1101001010011101",
39055 => "1101001010011111",
39056 => "1101001010100001",
39057 => "1101001010100100",
39058 => "1101001010100110",
39059 => "1101001010101000",
39060 => "1101001010101011",
39061 => "1101001010101101",
39062 => "1101001010101111",
39063 => "1101001010110010",
39064 => "1101001010110100",
39065 => "1101001010110110",
39066 => "1101001010111001",
39067 => "1101001010111011",
39068 => "1101001010111101",
39069 => "1101001011000000",
39070 => "1101001011000010",
39071 => "1101001011000100",
39072 => "1101001011000111",
39073 => "1101001011001001",
39074 => "1101001011001011",
39075 => "1101001011001110",
39076 => "1101001011010000",
39077 => "1101001011010010",
39078 => "1101001011010100",
39079 => "1101001011010111",
39080 => "1101001011011001",
39081 => "1101001011011011",
39082 => "1101001011011110",
39083 => "1101001011100000",
39084 => "1101001011100010",
39085 => "1101001011100101",
39086 => "1101001011100111",
39087 => "1101001011101001",
39088 => "1101001011101100",
39089 => "1101001011101110",
39090 => "1101001011110000",
39091 => "1101001011110011",
39092 => "1101001011110101",
39093 => "1101001011110111",
39094 => "1101001011111010",
39095 => "1101001011111100",
39096 => "1101001011111110",
39097 => "1101001100000001",
39098 => "1101001100000011",
39099 => "1101001100000101",
39100 => "1101001100001000",
39101 => "1101001100001010",
39102 => "1101001100001100",
39103 => "1101001100001111",
39104 => "1101001100010001",
39105 => "1101001100010011",
39106 => "1101001100010101",
39107 => "1101001100011000",
39108 => "1101001100011010",
39109 => "1101001100011100",
39110 => "1101001100011111",
39111 => "1101001100100001",
39112 => "1101001100100011",
39113 => "1101001100100110",
39114 => "1101001100101000",
39115 => "1101001100101010",
39116 => "1101001100101101",
39117 => "1101001100101111",
39118 => "1101001100110001",
39119 => "1101001100110100",
39120 => "1101001100110110",
39121 => "1101001100111000",
39122 => "1101001100111010",
39123 => "1101001100111101",
39124 => "1101001100111111",
39125 => "1101001101000001",
39126 => "1101001101000100",
39127 => "1101001101000110",
39128 => "1101001101001000",
39129 => "1101001101001011",
39130 => "1101001101001101",
39131 => "1101001101001111",
39132 => "1101001101010010",
39133 => "1101001101010100",
39134 => "1101001101010110",
39135 => "1101001101011000",
39136 => "1101001101011011",
39137 => "1101001101011101",
39138 => "1101001101011111",
39139 => "1101001101100010",
39140 => "1101001101100100",
39141 => "1101001101100110",
39142 => "1101001101101001",
39143 => "1101001101101011",
39144 => "1101001101101101",
39145 => "1101001101101111",
39146 => "1101001101110010",
39147 => "1101001101110100",
39148 => "1101001101110110",
39149 => "1101001101111001",
39150 => "1101001101111011",
39151 => "1101001101111101",
39152 => "1101001110000000",
39153 => "1101001110000010",
39154 => "1101001110000100",
39155 => "1101001110000110",
39156 => "1101001110001001",
39157 => "1101001110001011",
39158 => "1101001110001101",
39159 => "1101001110010000",
39160 => "1101001110010010",
39161 => "1101001110010100",
39162 => "1101001110010110",
39163 => "1101001110011001",
39164 => "1101001110011011",
39165 => "1101001110011101",
39166 => "1101001110100000",
39167 => "1101001110100010",
39168 => "1101001110100100",
39169 => "1101001110100111",
39170 => "1101001110101001",
39171 => "1101001110101011",
39172 => "1101001110101101",
39173 => "1101001110110000",
39174 => "1101001110110010",
39175 => "1101001110110100",
39176 => "1101001110110111",
39177 => "1101001110111001",
39178 => "1101001110111011",
39179 => "1101001110111101",
39180 => "1101001111000000",
39181 => "1101001111000010",
39182 => "1101001111000100",
39183 => "1101001111000111",
39184 => "1101001111001001",
39185 => "1101001111001011",
39186 => "1101001111001101",
39187 => "1101001111010000",
39188 => "1101001111010010",
39189 => "1101001111010100",
39190 => "1101001111010111",
39191 => "1101001111011001",
39192 => "1101001111011011",
39193 => "1101001111011101",
39194 => "1101001111100000",
39195 => "1101001111100010",
39196 => "1101001111100100",
39197 => "1101001111100111",
39198 => "1101001111101001",
39199 => "1101001111101011",
39200 => "1101001111101101",
39201 => "1101001111110000",
39202 => "1101001111110010",
39203 => "1101001111110100",
39204 => "1101001111110111",
39205 => "1101001111111001",
39206 => "1101001111111011",
39207 => "1101001111111101",
39208 => "1101010000000000",
39209 => "1101010000000010",
39210 => "1101010000000100",
39211 => "1101010000000110",
39212 => "1101010000001001",
39213 => "1101010000001011",
39214 => "1101010000001101",
39215 => "1101010000010000",
39216 => "1101010000010010",
39217 => "1101010000010100",
39218 => "1101010000010110",
39219 => "1101010000011001",
39220 => "1101010000011011",
39221 => "1101010000011101",
39222 => "1101010000011111",
39223 => "1101010000100010",
39224 => "1101010000100100",
39225 => "1101010000100110",
39226 => "1101010000101001",
39227 => "1101010000101011",
39228 => "1101010000101101",
39229 => "1101010000101111",
39230 => "1101010000110010",
39231 => "1101010000110100",
39232 => "1101010000110110",
39233 => "1101010000111000",
39234 => "1101010000111011",
39235 => "1101010000111101",
39236 => "1101010000111111",
39237 => "1101010001000010",
39238 => "1101010001000100",
39239 => "1101010001000110",
39240 => "1101010001001000",
39241 => "1101010001001011",
39242 => "1101010001001101",
39243 => "1101010001001111",
39244 => "1101010001010001",
39245 => "1101010001010100",
39246 => "1101010001010110",
39247 => "1101010001011000",
39248 => "1101010001011010",
39249 => "1101010001011101",
39250 => "1101010001011111",
39251 => "1101010001100001",
39252 => "1101010001100011",
39253 => "1101010001100110",
39254 => "1101010001101000",
39255 => "1101010001101010",
39256 => "1101010001101101",
39257 => "1101010001101111",
39258 => "1101010001110001",
39259 => "1101010001110011",
39260 => "1101010001110110",
39261 => "1101010001111000",
39262 => "1101010001111010",
39263 => "1101010001111100",
39264 => "1101010001111111",
39265 => "1101010010000001",
39266 => "1101010010000011",
39267 => "1101010010000101",
39268 => "1101010010001000",
39269 => "1101010010001010",
39270 => "1101010010001100",
39271 => "1101010010001110",
39272 => "1101010010010001",
39273 => "1101010010010011",
39274 => "1101010010010101",
39275 => "1101010010010111",
39276 => "1101010010011010",
39277 => "1101010010011100",
39278 => "1101010010011110",
39279 => "1101010010100000",
39280 => "1101010010100011",
39281 => "1101010010100101",
39282 => "1101010010100111",
39283 => "1101010010101001",
39284 => "1101010010101100",
39285 => "1101010010101110",
39286 => "1101010010110000",
39287 => "1101010010110010",
39288 => "1101010010110101",
39289 => "1101010010110111",
39290 => "1101010010111001",
39291 => "1101010010111011",
39292 => "1101010010111110",
39293 => "1101010011000000",
39294 => "1101010011000010",
39295 => "1101010011000100",
39296 => "1101010011000111",
39297 => "1101010011001001",
39298 => "1101010011001011",
39299 => "1101010011001101",
39300 => "1101010011010000",
39301 => "1101010011010010",
39302 => "1101010011010100",
39303 => "1101010011010110",
39304 => "1101010011011001",
39305 => "1101010011011011",
39306 => "1101010011011101",
39307 => "1101010011011111",
39308 => "1101010011100010",
39309 => "1101010011100100",
39310 => "1101010011100110",
39311 => "1101010011101000",
39312 => "1101010011101011",
39313 => "1101010011101101",
39314 => "1101010011101111",
39315 => "1101010011110001",
39316 => "1101010011110011",
39317 => "1101010011110110",
39318 => "1101010011111000",
39319 => "1101010011111010",
39320 => "1101010011111100",
39321 => "1101010011111111",
39322 => "1101010100000001",
39323 => "1101010100000011",
39324 => "1101010100000101",
39325 => "1101010100001000",
39326 => "1101010100001010",
39327 => "1101010100001100",
39328 => "1101010100001110",
39329 => "1101010100010001",
39330 => "1101010100010011",
39331 => "1101010100010101",
39332 => "1101010100010111",
39333 => "1101010100011001",
39334 => "1101010100011100",
39335 => "1101010100011110",
39336 => "1101010100100000",
39337 => "1101010100100010",
39338 => "1101010100100101",
39339 => "1101010100100111",
39340 => "1101010100101001",
39341 => "1101010100101011",
39342 => "1101010100101110",
39343 => "1101010100110000",
39344 => "1101010100110010",
39345 => "1101010100110100",
39346 => "1101010100110110",
39347 => "1101010100111001",
39348 => "1101010100111011",
39349 => "1101010100111101",
39350 => "1101010100111111",
39351 => "1101010101000010",
39352 => "1101010101000100",
39353 => "1101010101000110",
39354 => "1101010101001000",
39355 => "1101010101001010",
39356 => "1101010101001101",
39357 => "1101010101001111",
39358 => "1101010101010001",
39359 => "1101010101010011",
39360 => "1101010101010110",
39361 => "1101010101011000",
39362 => "1101010101011010",
39363 => "1101010101011100",
39364 => "1101010101011110",
39365 => "1101010101100001",
39366 => "1101010101100011",
39367 => "1101010101100101",
39368 => "1101010101100111",
39369 => "1101010101101010",
39370 => "1101010101101100",
39371 => "1101010101101110",
39372 => "1101010101110000",
39373 => "1101010101110010",
39374 => "1101010101110101",
39375 => "1101010101110111",
39376 => "1101010101111001",
39377 => "1101010101111011",
39378 => "1101010101111110",
39379 => "1101010110000000",
39380 => "1101010110000010",
39381 => "1101010110000100",
39382 => "1101010110000110",
39383 => "1101010110001001",
39384 => "1101010110001011",
39385 => "1101010110001101",
39386 => "1101010110001111",
39387 => "1101010110010001",
39388 => "1101010110010100",
39389 => "1101010110010110",
39390 => "1101010110011000",
39391 => "1101010110011010",
39392 => "1101010110011101",
39393 => "1101010110011111",
39394 => "1101010110100001",
39395 => "1101010110100011",
39396 => "1101010110100101",
39397 => "1101010110101000",
39398 => "1101010110101010",
39399 => "1101010110101100",
39400 => "1101010110101110",
39401 => "1101010110110000",
39402 => "1101010110110011",
39403 => "1101010110110101",
39404 => "1101010110110111",
39405 => "1101010110111001",
39406 => "1101010110111011",
39407 => "1101010110111110",
39408 => "1101010111000000",
39409 => "1101010111000010",
39410 => "1101010111000100",
39411 => "1101010111000110",
39412 => "1101010111001001",
39413 => "1101010111001011",
39414 => "1101010111001101",
39415 => "1101010111001111",
39416 => "1101010111010001",
39417 => "1101010111010100",
39418 => "1101010111010110",
39419 => "1101010111011000",
39420 => "1101010111011010",
39421 => "1101010111011100",
39422 => "1101010111011111",
39423 => "1101010111100001",
39424 => "1101010111100011",
39425 => "1101010111100101",
39426 => "1101010111100111",
39427 => "1101010111101010",
39428 => "1101010111101100",
39429 => "1101010111101110",
39430 => "1101010111110000",
39431 => "1101010111110010",
39432 => "1101010111110101",
39433 => "1101010111110111",
39434 => "1101010111111001",
39435 => "1101010111111011",
39436 => "1101010111111101",
39437 => "1101011000000000",
39438 => "1101011000000010",
39439 => "1101011000000100",
39440 => "1101011000000110",
39441 => "1101011000001000",
39442 => "1101011000001011",
39443 => "1101011000001101",
39444 => "1101011000001111",
39445 => "1101011000010001",
39446 => "1101011000010011",
39447 => "1101011000010110",
39448 => "1101011000011000",
39449 => "1101011000011010",
39450 => "1101011000011100",
39451 => "1101011000011110",
39452 => "1101011000100001",
39453 => "1101011000100011",
39454 => "1101011000100101",
39455 => "1101011000100111",
39456 => "1101011000101001",
39457 => "1101011000101011",
39458 => "1101011000101110",
39459 => "1101011000110000",
39460 => "1101011000110010",
39461 => "1101011000110100",
39462 => "1101011000110110",
39463 => "1101011000111001",
39464 => "1101011000111011",
39465 => "1101011000111101",
39466 => "1101011000111111",
39467 => "1101011001000001",
39468 => "1101011001000011",
39469 => "1101011001000110",
39470 => "1101011001001000",
39471 => "1101011001001010",
39472 => "1101011001001100",
39473 => "1101011001001110",
39474 => "1101011001010001",
39475 => "1101011001010011",
39476 => "1101011001010101",
39477 => "1101011001010111",
39478 => "1101011001011001",
39479 => "1101011001011011",
39480 => "1101011001011110",
39481 => "1101011001100000",
39482 => "1101011001100010",
39483 => "1101011001100100",
39484 => "1101011001100110",
39485 => "1101011001101001",
39486 => "1101011001101011",
39487 => "1101011001101101",
39488 => "1101011001101111",
39489 => "1101011001110001",
39490 => "1101011001110011",
39491 => "1101011001110110",
39492 => "1101011001111000",
39493 => "1101011001111010",
39494 => "1101011001111100",
39495 => "1101011001111110",
39496 => "1101011010000000",
39497 => "1101011010000011",
39498 => "1101011010000101",
39499 => "1101011010000111",
39500 => "1101011010001001",
39501 => "1101011010001011",
39502 => "1101011010001110",
39503 => "1101011010010000",
39504 => "1101011010010010",
39505 => "1101011010010100",
39506 => "1101011010010110",
39507 => "1101011010011000",
39508 => "1101011010011011",
39509 => "1101011010011101",
39510 => "1101011010011111",
39511 => "1101011010100001",
39512 => "1101011010100011",
39513 => "1101011010100101",
39514 => "1101011010101000",
39515 => "1101011010101010",
39516 => "1101011010101100",
39517 => "1101011010101110",
39518 => "1101011010110000",
39519 => "1101011010110010",
39520 => "1101011010110101",
39521 => "1101011010110111",
39522 => "1101011010111001",
39523 => "1101011010111011",
39524 => "1101011010111101",
39525 => "1101011010111111",
39526 => "1101011011000010",
39527 => "1101011011000100",
39528 => "1101011011000110",
39529 => "1101011011001000",
39530 => "1101011011001010",
39531 => "1101011011001100",
39532 => "1101011011001110",
39533 => "1101011011010001",
39534 => "1101011011010011",
39535 => "1101011011010101",
39536 => "1101011011010111",
39537 => "1101011011011001",
39538 => "1101011011011011",
39539 => "1101011011011110",
39540 => "1101011011100000",
39541 => "1101011011100010",
39542 => "1101011011100100",
39543 => "1101011011100110",
39544 => "1101011011101000",
39545 => "1101011011101011",
39546 => "1101011011101101",
39547 => "1101011011101111",
39548 => "1101011011110001",
39549 => "1101011011110011",
39550 => "1101011011110101",
39551 => "1101011011110111",
39552 => "1101011011111010",
39553 => "1101011011111100",
39554 => "1101011011111110",
39555 => "1101011100000000",
39556 => "1101011100000010",
39557 => "1101011100000100",
39558 => "1101011100000111",
39559 => "1101011100001001",
39560 => "1101011100001011",
39561 => "1101011100001101",
39562 => "1101011100001111",
39563 => "1101011100010001",
39564 => "1101011100010011",
39565 => "1101011100010110",
39566 => "1101011100011000",
39567 => "1101011100011010",
39568 => "1101011100011100",
39569 => "1101011100011110",
39570 => "1101011100100000",
39571 => "1101011100100010",
39572 => "1101011100100101",
39573 => "1101011100100111",
39574 => "1101011100101001",
39575 => "1101011100101011",
39576 => "1101011100101101",
39577 => "1101011100101111",
39578 => "1101011100110001",
39579 => "1101011100110100",
39580 => "1101011100110110",
39581 => "1101011100111000",
39582 => "1101011100111010",
39583 => "1101011100111100",
39584 => "1101011100111110",
39585 => "1101011101000000",
39586 => "1101011101000011",
39587 => "1101011101000101",
39588 => "1101011101000111",
39589 => "1101011101001001",
39590 => "1101011101001011",
39591 => "1101011101001101",
39592 => "1101011101001111",
39593 => "1101011101010010",
39594 => "1101011101010100",
39595 => "1101011101010110",
39596 => "1101011101011000",
39597 => "1101011101011010",
39598 => "1101011101011100",
39599 => "1101011101011110",
39600 => "1101011101100001",
39601 => "1101011101100011",
39602 => "1101011101100101",
39603 => "1101011101100111",
39604 => "1101011101101001",
39605 => "1101011101101011",
39606 => "1101011101101101",
39607 => "1101011101101111",
39608 => "1101011101110010",
39609 => "1101011101110100",
39610 => "1101011101110110",
39611 => "1101011101111000",
39612 => "1101011101111010",
39613 => "1101011101111100",
39614 => "1101011101111110",
39615 => "1101011110000001",
39616 => "1101011110000011",
39617 => "1101011110000101",
39618 => "1101011110000111",
39619 => "1101011110001001",
39620 => "1101011110001011",
39621 => "1101011110001101",
39622 => "1101011110001111",
39623 => "1101011110010010",
39624 => "1101011110010100",
39625 => "1101011110010110",
39626 => "1101011110011000",
39627 => "1101011110011010",
39628 => "1101011110011100",
39629 => "1101011110011110",
39630 => "1101011110100000",
39631 => "1101011110100011",
39632 => "1101011110100101",
39633 => "1101011110100111",
39634 => "1101011110101001",
39635 => "1101011110101011",
39636 => "1101011110101101",
39637 => "1101011110101111",
39638 => "1101011110110001",
39639 => "1101011110110100",
39640 => "1101011110110110",
39641 => "1101011110111000",
39642 => "1101011110111010",
39643 => "1101011110111100",
39644 => "1101011110111110",
39645 => "1101011111000000",
39646 => "1101011111000010",
39647 => "1101011111000101",
39648 => "1101011111000111",
39649 => "1101011111001001",
39650 => "1101011111001011",
39651 => "1101011111001101",
39652 => "1101011111001111",
39653 => "1101011111010001",
39654 => "1101011111010011",
39655 => "1101011111010101",
39656 => "1101011111011000",
39657 => "1101011111011010",
39658 => "1101011111011100",
39659 => "1101011111011110",
39660 => "1101011111100000",
39661 => "1101011111100010",
39662 => "1101011111100100",
39663 => "1101011111100110",
39664 => "1101011111101001",
39665 => "1101011111101011",
39666 => "1101011111101101",
39667 => "1101011111101111",
39668 => "1101011111110001",
39669 => "1101011111110011",
39670 => "1101011111110101",
39671 => "1101011111110111",
39672 => "1101011111111001",
39673 => "1101011111111100",
39674 => "1101011111111110",
39675 => "1101100000000000",
39676 => "1101100000000010",
39677 => "1101100000000100",
39678 => "1101100000000110",
39679 => "1101100000001000",
39680 => "1101100000001010",
39681 => "1101100000001100",
39682 => "1101100000001111",
39683 => "1101100000010001",
39684 => "1101100000010011",
39685 => "1101100000010101",
39686 => "1101100000010111",
39687 => "1101100000011001",
39688 => "1101100000011011",
39689 => "1101100000011101",
39690 => "1101100000011111",
39691 => "1101100000100001",
39692 => "1101100000100100",
39693 => "1101100000100110",
39694 => "1101100000101000",
39695 => "1101100000101010",
39696 => "1101100000101100",
39697 => "1101100000101110",
39698 => "1101100000110000",
39699 => "1101100000110010",
39700 => "1101100000110100",
39701 => "1101100000110110",
39702 => "1101100000111001",
39703 => "1101100000111011",
39704 => "1101100000111101",
39705 => "1101100000111111",
39706 => "1101100001000001",
39707 => "1101100001000011",
39708 => "1101100001000101",
39709 => "1101100001000111",
39710 => "1101100001001001",
39711 => "1101100001001011",
39712 => "1101100001001110",
39713 => "1101100001010000",
39714 => "1101100001010010",
39715 => "1101100001010100",
39716 => "1101100001010110",
39717 => "1101100001011000",
39718 => "1101100001011010",
39719 => "1101100001011100",
39720 => "1101100001011110",
39721 => "1101100001100000",
39722 => "1101100001100010",
39723 => "1101100001100101",
39724 => "1101100001100111",
39725 => "1101100001101001",
39726 => "1101100001101011",
39727 => "1101100001101101",
39728 => "1101100001101111",
39729 => "1101100001110001",
39730 => "1101100001110011",
39731 => "1101100001110101",
39732 => "1101100001110111",
39733 => "1101100001111001",
39734 => "1101100001111100",
39735 => "1101100001111110",
39736 => "1101100010000000",
39737 => "1101100010000010",
39738 => "1101100010000100",
39739 => "1101100010000110",
39740 => "1101100010001000",
39741 => "1101100010001010",
39742 => "1101100010001100",
39743 => "1101100010001110",
39744 => "1101100010010000",
39745 => "1101100010010011",
39746 => "1101100010010101",
39747 => "1101100010010111",
39748 => "1101100010011001",
39749 => "1101100010011011",
39750 => "1101100010011101",
39751 => "1101100010011111",
39752 => "1101100010100001",
39753 => "1101100010100011",
39754 => "1101100010100101",
39755 => "1101100010100111",
39756 => "1101100010101001",
39757 => "1101100010101100",
39758 => "1101100010101110",
39759 => "1101100010110000",
39760 => "1101100010110010",
39761 => "1101100010110100",
39762 => "1101100010110110",
39763 => "1101100010111000",
39764 => "1101100010111010",
39765 => "1101100010111100",
39766 => "1101100010111110",
39767 => "1101100011000000",
39768 => "1101100011000010",
39769 => "1101100011000100",
39770 => "1101100011000111",
39771 => "1101100011001001",
39772 => "1101100011001011",
39773 => "1101100011001101",
39774 => "1101100011001111",
39775 => "1101100011010001",
39776 => "1101100011010011",
39777 => "1101100011010101",
39778 => "1101100011010111",
39779 => "1101100011011001",
39780 => "1101100011011011",
39781 => "1101100011011101",
39782 => "1101100011011111",
39783 => "1101100011100001",
39784 => "1101100011100100",
39785 => "1101100011100110",
39786 => "1101100011101000",
39787 => "1101100011101010",
39788 => "1101100011101100",
39789 => "1101100011101110",
39790 => "1101100011110000",
39791 => "1101100011110010",
39792 => "1101100011110100",
39793 => "1101100011110110",
39794 => "1101100011111000",
39795 => "1101100011111010",
39796 => "1101100011111100",
39797 => "1101100011111110",
39798 => "1101100100000001",
39799 => "1101100100000011",
39800 => "1101100100000101",
39801 => "1101100100000111",
39802 => "1101100100001001",
39803 => "1101100100001011",
39804 => "1101100100001101",
39805 => "1101100100001111",
39806 => "1101100100010001",
39807 => "1101100100010011",
39808 => "1101100100010101",
39809 => "1101100100010111",
39810 => "1101100100011001",
39811 => "1101100100011011",
39812 => "1101100100011101",
39813 => "1101100100011111",
39814 => "1101100100100010",
39815 => "1101100100100100",
39816 => "1101100100100110",
39817 => "1101100100101000",
39818 => "1101100100101010",
39819 => "1101100100101100",
39820 => "1101100100101110",
39821 => "1101100100110000",
39822 => "1101100100110010",
39823 => "1101100100110100",
39824 => "1101100100110110",
39825 => "1101100100111000",
39826 => "1101100100111010",
39827 => "1101100100111100",
39828 => "1101100100111110",
39829 => "1101100101000000",
39830 => "1101100101000010",
39831 => "1101100101000101",
39832 => "1101100101000111",
39833 => "1101100101001001",
39834 => "1101100101001011",
39835 => "1101100101001101",
39836 => "1101100101001111",
39837 => "1101100101010001",
39838 => "1101100101010011",
39839 => "1101100101010101",
39840 => "1101100101010111",
39841 => "1101100101011001",
39842 => "1101100101011011",
39843 => "1101100101011101",
39844 => "1101100101011111",
39845 => "1101100101100001",
39846 => "1101100101100011",
39847 => "1101100101100101",
39848 => "1101100101100111",
39849 => "1101100101101001",
39850 => "1101100101101011",
39851 => "1101100101101110",
39852 => "1101100101110000",
39853 => "1101100101110010",
39854 => "1101100101110100",
39855 => "1101100101110110",
39856 => "1101100101111000",
39857 => "1101100101111010",
39858 => "1101100101111100",
39859 => "1101100101111110",
39860 => "1101100110000000",
39861 => "1101100110000010",
39862 => "1101100110000100",
39863 => "1101100110000110",
39864 => "1101100110001000",
39865 => "1101100110001010",
39866 => "1101100110001100",
39867 => "1101100110001110",
39868 => "1101100110010000",
39869 => "1101100110010010",
39870 => "1101100110010100",
39871 => "1101100110010110",
39872 => "1101100110011000",
39873 => "1101100110011010",
39874 => "1101100110011101",
39875 => "1101100110011111",
39876 => "1101100110100001",
39877 => "1101100110100011",
39878 => "1101100110100101",
39879 => "1101100110100111",
39880 => "1101100110101001",
39881 => "1101100110101011",
39882 => "1101100110101101",
39883 => "1101100110101111",
39884 => "1101100110110001",
39885 => "1101100110110011",
39886 => "1101100110110101",
39887 => "1101100110110111",
39888 => "1101100110111001",
39889 => "1101100110111011",
39890 => "1101100110111101",
39891 => "1101100110111111",
39892 => "1101100111000001",
39893 => "1101100111000011",
39894 => "1101100111000101",
39895 => "1101100111000111",
39896 => "1101100111001001",
39897 => "1101100111001011",
39898 => "1101100111001101",
39899 => "1101100111001111",
39900 => "1101100111010001",
39901 => "1101100111010011",
39902 => "1101100111010101",
39903 => "1101100111011000",
39904 => "1101100111011010",
39905 => "1101100111011100",
39906 => "1101100111011110",
39907 => "1101100111100000",
39908 => "1101100111100010",
39909 => "1101100111100100",
39910 => "1101100111100110",
39911 => "1101100111101000",
39912 => "1101100111101010",
39913 => "1101100111101100",
39914 => "1101100111101110",
39915 => "1101100111110000",
39916 => "1101100111110010",
39917 => "1101100111110100",
39918 => "1101100111110110",
39919 => "1101100111111000",
39920 => "1101100111111010",
39921 => "1101100111111100",
39922 => "1101100111111110",
39923 => "1101101000000000",
39924 => "1101101000000010",
39925 => "1101101000000100",
39926 => "1101101000000110",
39927 => "1101101000001000",
39928 => "1101101000001010",
39929 => "1101101000001100",
39930 => "1101101000001110",
39931 => "1101101000010000",
39932 => "1101101000010010",
39933 => "1101101000010100",
39934 => "1101101000010110",
39935 => "1101101000011000",
39936 => "1101101000011010",
39937 => "1101101000011100",
39938 => "1101101000011110",
39939 => "1101101000100000",
39940 => "1101101000100010",
39941 => "1101101000100100",
39942 => "1101101000100110",
39943 => "1101101000101000",
39944 => "1101101000101010",
39945 => "1101101000101100",
39946 => "1101101000101110",
39947 => "1101101000110000",
39948 => "1101101000110010",
39949 => "1101101000110101",
39950 => "1101101000110111",
39951 => "1101101000111001",
39952 => "1101101000111011",
39953 => "1101101000111101",
39954 => "1101101000111111",
39955 => "1101101001000001",
39956 => "1101101001000011",
39957 => "1101101001000101",
39958 => "1101101001000111",
39959 => "1101101001001001",
39960 => "1101101001001011",
39961 => "1101101001001101",
39962 => "1101101001001111",
39963 => "1101101001010001",
39964 => "1101101001010011",
39965 => "1101101001010101",
39966 => "1101101001010111",
39967 => "1101101001011001",
39968 => "1101101001011011",
39969 => "1101101001011101",
39970 => "1101101001011111",
39971 => "1101101001100001",
39972 => "1101101001100011",
39973 => "1101101001100101",
39974 => "1101101001100111",
39975 => "1101101001101001",
39976 => "1101101001101011",
39977 => "1101101001101101",
39978 => "1101101001101111",
39979 => "1101101001110001",
39980 => "1101101001110011",
39981 => "1101101001110101",
39982 => "1101101001110111",
39983 => "1101101001111001",
39984 => "1101101001111011",
39985 => "1101101001111101",
39986 => "1101101001111111",
39987 => "1101101010000001",
39988 => "1101101010000011",
39989 => "1101101010000101",
39990 => "1101101010000111",
39991 => "1101101010001001",
39992 => "1101101010001011",
39993 => "1101101010001101",
39994 => "1101101010001111",
39995 => "1101101010010001",
39996 => "1101101010010011",
39997 => "1101101010010101",
39998 => "1101101010010111",
39999 => "1101101010011001",
40000 => "1101101010011011",
40001 => "1101101010011101",
40002 => "1101101010011111",
40003 => "1101101010100001",
40004 => "1101101010100011",
40005 => "1101101010100101",
40006 => "1101101010100111",
40007 => "1101101010101001",
40008 => "1101101010101011",
40009 => "1101101010101101",
40010 => "1101101010101111",
40011 => "1101101010110001",
40012 => "1101101010110011",
40013 => "1101101010110101",
40014 => "1101101010110111",
40015 => "1101101010111001",
40016 => "1101101010111011",
40017 => "1101101010111101",
40018 => "1101101010111111",
40019 => "1101101011000001",
40020 => "1101101011000011",
40021 => "1101101011000101",
40022 => "1101101011000111",
40023 => "1101101011001001",
40024 => "1101101011001011",
40025 => "1101101011001101",
40026 => "1101101011001111",
40027 => "1101101011010001",
40028 => "1101101011010010",
40029 => "1101101011010100",
40030 => "1101101011010110",
40031 => "1101101011011000",
40032 => "1101101011011010",
40033 => "1101101011011100",
40034 => "1101101011011110",
40035 => "1101101011100000",
40036 => "1101101011100010",
40037 => "1101101011100100",
40038 => "1101101011100110",
40039 => "1101101011101000",
40040 => "1101101011101010",
40041 => "1101101011101100",
40042 => "1101101011101110",
40043 => "1101101011110000",
40044 => "1101101011110010",
40045 => "1101101011110100",
40046 => "1101101011110110",
40047 => "1101101011111000",
40048 => "1101101011111010",
40049 => "1101101011111100",
40050 => "1101101011111110",
40051 => "1101101100000000",
40052 => "1101101100000010",
40053 => "1101101100000100",
40054 => "1101101100000110",
40055 => "1101101100001000",
40056 => "1101101100001010",
40057 => "1101101100001100",
40058 => "1101101100001110",
40059 => "1101101100010000",
40060 => "1101101100010010",
40061 => "1101101100010100",
40062 => "1101101100010110",
40063 => "1101101100011000",
40064 => "1101101100011010",
40065 => "1101101100011100",
40066 => "1101101100011110",
40067 => "1101101100100000",
40068 => "1101101100100010",
40069 => "1101101100100100",
40070 => "1101101100100110",
40071 => "1101101100101000",
40072 => "1101101100101010",
40073 => "1101101100101100",
40074 => "1101101100101101",
40075 => "1101101100101111",
40076 => "1101101100110001",
40077 => "1101101100110011",
40078 => "1101101100110101",
40079 => "1101101100110111",
40080 => "1101101100111001",
40081 => "1101101100111011",
40082 => "1101101100111101",
40083 => "1101101100111111",
40084 => "1101101101000001",
40085 => "1101101101000011",
40086 => "1101101101000101",
40087 => "1101101101000111",
40088 => "1101101101001001",
40089 => "1101101101001011",
40090 => "1101101101001101",
40091 => "1101101101001111",
40092 => "1101101101010001",
40093 => "1101101101010011",
40094 => "1101101101010101",
40095 => "1101101101010111",
40096 => "1101101101011001",
40097 => "1101101101011011",
40098 => "1101101101011101",
40099 => "1101101101011111",
40100 => "1101101101100001",
40101 => "1101101101100011",
40102 => "1101101101100101",
40103 => "1101101101100110",
40104 => "1101101101101000",
40105 => "1101101101101010",
40106 => "1101101101101100",
40107 => "1101101101101110",
40108 => "1101101101110000",
40109 => "1101101101110010",
40110 => "1101101101110100",
40111 => "1101101101110110",
40112 => "1101101101111000",
40113 => "1101101101111010",
40114 => "1101101101111100",
40115 => "1101101101111110",
40116 => "1101101110000000",
40117 => "1101101110000010",
40118 => "1101101110000100",
40119 => "1101101110000110",
40120 => "1101101110001000",
40121 => "1101101110001010",
40122 => "1101101110001100",
40123 => "1101101110001110",
40124 => "1101101110010000",
40125 => "1101101110010010",
40126 => "1101101110010011",
40127 => "1101101110010101",
40128 => "1101101110010111",
40129 => "1101101110011001",
40130 => "1101101110011011",
40131 => "1101101110011101",
40132 => "1101101110011111",
40133 => "1101101110100001",
40134 => "1101101110100011",
40135 => "1101101110100101",
40136 => "1101101110100111",
40137 => "1101101110101001",
40138 => "1101101110101011",
40139 => "1101101110101101",
40140 => "1101101110101111",
40141 => "1101101110110001",
40142 => "1101101110110011",
40143 => "1101101110110101",
40144 => "1101101110110111",
40145 => "1101101110111001",
40146 => "1101101110111010",
40147 => "1101101110111100",
40148 => "1101101110111110",
40149 => "1101101111000000",
40150 => "1101101111000010",
40151 => "1101101111000100",
40152 => "1101101111000110",
40153 => "1101101111001000",
40154 => "1101101111001010",
40155 => "1101101111001100",
40156 => "1101101111001110",
40157 => "1101101111010000",
40158 => "1101101111010010",
40159 => "1101101111010100",
40160 => "1101101111010110",
40161 => "1101101111011000",
40162 => "1101101111011010",
40163 => "1101101111011011",
40164 => "1101101111011101",
40165 => "1101101111011111",
40166 => "1101101111100001",
40167 => "1101101111100011",
40168 => "1101101111100101",
40169 => "1101101111100111",
40170 => "1101101111101001",
40171 => "1101101111101011",
40172 => "1101101111101101",
40173 => "1101101111101111",
40174 => "1101101111110001",
40175 => "1101101111110011",
40176 => "1101101111110101",
40177 => "1101101111110111",
40178 => "1101101111111001",
40179 => "1101101111111010",
40180 => "1101101111111100",
40181 => "1101101111111110",
40182 => "1101110000000000",
40183 => "1101110000000010",
40184 => "1101110000000100",
40185 => "1101110000000110",
40186 => "1101110000001000",
40187 => "1101110000001010",
40188 => "1101110000001100",
40189 => "1101110000001110",
40190 => "1101110000010000",
40191 => "1101110000010010",
40192 => "1101110000010100",
40193 => "1101110000010110",
40194 => "1101110000010111",
40195 => "1101110000011001",
40196 => "1101110000011011",
40197 => "1101110000011101",
40198 => "1101110000011111",
40199 => "1101110000100001",
40200 => "1101110000100011",
40201 => "1101110000100101",
40202 => "1101110000100111",
40203 => "1101110000101001",
40204 => "1101110000101011",
40205 => "1101110000101101",
40206 => "1101110000101111",
40207 => "1101110000110001",
40208 => "1101110000110010",
40209 => "1101110000110100",
40210 => "1101110000110110",
40211 => "1101110000111000",
40212 => "1101110000111010",
40213 => "1101110000111100",
40214 => "1101110000111110",
40215 => "1101110001000000",
40216 => "1101110001000010",
40217 => "1101110001000100",
40218 => "1101110001000110",
40219 => "1101110001001000",
40220 => "1101110001001010",
40221 => "1101110001001011",
40222 => "1101110001001101",
40223 => "1101110001001111",
40224 => "1101110001010001",
40225 => "1101110001010011",
40226 => "1101110001010101",
40227 => "1101110001010111",
40228 => "1101110001011001",
40229 => "1101110001011011",
40230 => "1101110001011101",
40231 => "1101110001011111",
40232 => "1101110001100001",
40233 => "1101110001100010",
40234 => "1101110001100100",
40235 => "1101110001100110",
40236 => "1101110001101000",
40237 => "1101110001101010",
40238 => "1101110001101100",
40239 => "1101110001101110",
40240 => "1101110001110000",
40241 => "1101110001110010",
40242 => "1101110001110100",
40243 => "1101110001110110",
40244 => "1101110001111000",
40245 => "1101110001111001",
40246 => "1101110001111011",
40247 => "1101110001111101",
40248 => "1101110001111111",
40249 => "1101110010000001",
40250 => "1101110010000011",
40251 => "1101110010000101",
40252 => "1101110010000111",
40253 => "1101110010001001",
40254 => "1101110010001011",
40255 => "1101110010001101",
40256 => "1101110010001110",
40257 => "1101110010010000",
40258 => "1101110010010010",
40259 => "1101110010010100",
40260 => "1101110010010110",
40261 => "1101110010011000",
40262 => "1101110010011010",
40263 => "1101110010011100",
40264 => "1101110010011110",
40265 => "1101110010100000",
40266 => "1101110010100010",
40267 => "1101110010100011",
40268 => "1101110010100101",
40269 => "1101110010100111",
40270 => "1101110010101001",
40271 => "1101110010101011",
40272 => "1101110010101101",
40273 => "1101110010101111",
40274 => "1101110010110001",
40275 => "1101110010110011",
40276 => "1101110010110101",
40277 => "1101110010110110",
40278 => "1101110010111000",
40279 => "1101110010111010",
40280 => "1101110010111100",
40281 => "1101110010111110",
40282 => "1101110011000000",
40283 => "1101110011000010",
40284 => "1101110011000100",
40285 => "1101110011000110",
40286 => "1101110011001000",
40287 => "1101110011001001",
40288 => "1101110011001011",
40289 => "1101110011001101",
40290 => "1101110011001111",
40291 => "1101110011010001",
40292 => "1101110011010011",
40293 => "1101110011010101",
40294 => "1101110011010111",
40295 => "1101110011011001",
40296 => "1101110011011011",
40297 => "1101110011011100",
40298 => "1101110011011110",
40299 => "1101110011100000",
40300 => "1101110011100010",
40301 => "1101110011100100",
40302 => "1101110011100110",
40303 => "1101110011101000",
40304 => "1101110011101010",
40305 => "1101110011101100",
40306 => "1101110011101101",
40307 => "1101110011101111",
40308 => "1101110011110001",
40309 => "1101110011110011",
40310 => "1101110011110101",
40311 => "1101110011110111",
40312 => "1101110011111001",
40313 => "1101110011111011",
40314 => "1101110011111101",
40315 => "1101110011111110",
40316 => "1101110100000000",
40317 => "1101110100000010",
40318 => "1101110100000100",
40319 => "1101110100000110",
40320 => "1101110100001000",
40321 => "1101110100001010",
40322 => "1101110100001100",
40323 => "1101110100001110",
40324 => "1101110100001111",
40325 => "1101110100010001",
40326 => "1101110100010011",
40327 => "1101110100010101",
40328 => "1101110100010111",
40329 => "1101110100011001",
40330 => "1101110100011011",
40331 => "1101110100011101",
40332 => "1101110100011111",
40333 => "1101110100100000",
40334 => "1101110100100010",
40335 => "1101110100100100",
40336 => "1101110100100110",
40337 => "1101110100101000",
40338 => "1101110100101010",
40339 => "1101110100101100",
40340 => "1101110100101110",
40341 => "1101110100101111",
40342 => "1101110100110001",
40343 => "1101110100110011",
40344 => "1101110100110101",
40345 => "1101110100110111",
40346 => "1101110100111001",
40347 => "1101110100111011",
40348 => "1101110100111101",
40349 => "1101110100111110",
40350 => "1101110101000000",
40351 => "1101110101000010",
40352 => "1101110101000100",
40353 => "1101110101000110",
40354 => "1101110101001000",
40355 => "1101110101001010",
40356 => "1101110101001100",
40357 => "1101110101001101",
40358 => "1101110101001111",
40359 => "1101110101010001",
40360 => "1101110101010011",
40361 => "1101110101010101",
40362 => "1101110101010111",
40363 => "1101110101011001",
40364 => "1101110101011011",
40365 => "1101110101011100",
40366 => "1101110101011110",
40367 => "1101110101100000",
40368 => "1101110101100010",
40369 => "1101110101100100",
40370 => "1101110101100110",
40371 => "1101110101101000",
40372 => "1101110101101010",
40373 => "1101110101101011",
40374 => "1101110101101101",
40375 => "1101110101101111",
40376 => "1101110101110001",
40377 => "1101110101110011",
40378 => "1101110101110101",
40379 => "1101110101110111",
40380 => "1101110101111001",
40381 => "1101110101111010",
40382 => "1101110101111100",
40383 => "1101110101111110",
40384 => "1101110110000000",
40385 => "1101110110000010",
40386 => "1101110110000100",
40387 => "1101110110000110",
40388 => "1101110110000111",
40389 => "1101110110001001",
40390 => "1101110110001011",
40391 => "1101110110001101",
40392 => "1101110110001111",
40393 => "1101110110010001",
40394 => "1101110110010011",
40395 => "1101110110010100",
40396 => "1101110110010110",
40397 => "1101110110011000",
40398 => "1101110110011010",
40399 => "1101110110011100",
40400 => "1101110110011110",
40401 => "1101110110100000",
40402 => "1101110110100010",
40403 => "1101110110100011",
40404 => "1101110110100101",
40405 => "1101110110100111",
40406 => "1101110110101001",
40407 => "1101110110101011",
40408 => "1101110110101101",
40409 => "1101110110101111",
40410 => "1101110110110000",
40411 => "1101110110110010",
40412 => "1101110110110100",
40413 => "1101110110110110",
40414 => "1101110110111000",
40415 => "1101110110111010",
40416 => "1101110110111100",
40417 => "1101110110111101",
40418 => "1101110110111111",
40419 => "1101110111000001",
40420 => "1101110111000011",
40421 => "1101110111000101",
40422 => "1101110111000111",
40423 => "1101110111001000",
40424 => "1101110111001010",
40425 => "1101110111001100",
40426 => "1101110111001110",
40427 => "1101110111010000",
40428 => "1101110111010010",
40429 => "1101110111010100",
40430 => "1101110111010101",
40431 => "1101110111010111",
40432 => "1101110111011001",
40433 => "1101110111011011",
40434 => "1101110111011101",
40435 => "1101110111011111",
40436 => "1101110111100001",
40437 => "1101110111100010",
40438 => "1101110111100100",
40439 => "1101110111100110",
40440 => "1101110111101000",
40441 => "1101110111101010",
40442 => "1101110111101100",
40443 => "1101110111101101",
40444 => "1101110111101111",
40445 => "1101110111110001",
40446 => "1101110111110011",
40447 => "1101110111110101",
40448 => "1101110111110111",
40449 => "1101110111111001",
40450 => "1101110111111010",
40451 => "1101110111111100",
40452 => "1101110111111110",
40453 => "1101111000000000",
40454 => "1101111000000010",
40455 => "1101111000000100",
40456 => "1101111000000101",
40457 => "1101111000000111",
40458 => "1101111000001001",
40459 => "1101111000001011",
40460 => "1101111000001101",
40461 => "1101111000001111",
40462 => "1101111000010000",
40463 => "1101111000010010",
40464 => "1101111000010100",
40465 => "1101111000010110",
40466 => "1101111000011000",
40467 => "1101111000011010",
40468 => "1101111000011100",
40469 => "1101111000011101",
40470 => "1101111000011111",
40471 => "1101111000100001",
40472 => "1101111000100011",
40473 => "1101111000100101",
40474 => "1101111000100111",
40475 => "1101111000101000",
40476 => "1101111000101010",
40477 => "1101111000101100",
40478 => "1101111000101110",
40479 => "1101111000110000",
40480 => "1101111000110010",
40481 => "1101111000110011",
40482 => "1101111000110101",
40483 => "1101111000110111",
40484 => "1101111000111001",
40485 => "1101111000111011",
40486 => "1101111000111101",
40487 => "1101111000111110",
40488 => "1101111001000000",
40489 => "1101111001000010",
40490 => "1101111001000100",
40491 => "1101111001000110",
40492 => "1101111001001000",
40493 => "1101111001001001",
40494 => "1101111001001011",
40495 => "1101111001001101",
40496 => "1101111001001111",
40497 => "1101111001010001",
40498 => "1101111001010011",
40499 => "1101111001010100",
40500 => "1101111001010110",
40501 => "1101111001011000",
40502 => "1101111001011010",
40503 => "1101111001011100",
40504 => "1101111001011101",
40505 => "1101111001011111",
40506 => "1101111001100001",
40507 => "1101111001100011",
40508 => "1101111001100101",
40509 => "1101111001100111",
40510 => "1101111001101000",
40511 => "1101111001101010",
40512 => "1101111001101100",
40513 => "1101111001101110",
40514 => "1101111001110000",
40515 => "1101111001110010",
40516 => "1101111001110011",
40517 => "1101111001110101",
40518 => "1101111001110111",
40519 => "1101111001111001",
40520 => "1101111001111011",
40521 => "1101111001111100",
40522 => "1101111001111110",
40523 => "1101111010000000",
40524 => "1101111010000010",
40525 => "1101111010000100",
40526 => "1101111010000110",
40527 => "1101111010000111",
40528 => "1101111010001001",
40529 => "1101111010001011",
40530 => "1101111010001101",
40531 => "1101111010001111",
40532 => "1101111010010000",
40533 => "1101111010010010",
40534 => "1101111010010100",
40535 => "1101111010010110",
40536 => "1101111010011000",
40537 => "1101111010011010",
40538 => "1101111010011011",
40539 => "1101111010011101",
40540 => "1101111010011111",
40541 => "1101111010100001",
40542 => "1101111010100011",
40543 => "1101111010100100",
40544 => "1101111010100110",
40545 => "1101111010101000",
40546 => "1101111010101010",
40547 => "1101111010101100",
40548 => "1101111010101101",
40549 => "1101111010101111",
40550 => "1101111010110001",
40551 => "1101111010110011",
40552 => "1101111010110101",
40553 => "1101111010110111",
40554 => "1101111010111000",
40555 => "1101111010111010",
40556 => "1101111010111100",
40557 => "1101111010111110",
40558 => "1101111011000000",
40559 => "1101111011000001",
40560 => "1101111011000011",
40561 => "1101111011000101",
40562 => "1101111011000111",
40563 => "1101111011001001",
40564 => "1101111011001010",
40565 => "1101111011001100",
40566 => "1101111011001110",
40567 => "1101111011010000",
40568 => "1101111011010010",
40569 => "1101111011010011",
40570 => "1101111011010101",
40571 => "1101111011010111",
40572 => "1101111011011001",
40573 => "1101111011011011",
40574 => "1101111011011100",
40575 => "1101111011011110",
40576 => "1101111011100000",
40577 => "1101111011100010",
40578 => "1101111011100100",
40579 => "1101111011100101",
40580 => "1101111011100111",
40581 => "1101111011101001",
40582 => "1101111011101011",
40583 => "1101111011101101",
40584 => "1101111011101110",
40585 => "1101111011110000",
40586 => "1101111011110010",
40587 => "1101111011110100",
40588 => "1101111011110110",
40589 => "1101111011110111",
40590 => "1101111011111001",
40591 => "1101111011111011",
40592 => "1101111011111101",
40593 => "1101111011111111",
40594 => "1101111100000000",
40595 => "1101111100000010",
40596 => "1101111100000100",
40597 => "1101111100000110",
40598 => "1101111100001000",
40599 => "1101111100001001",
40600 => "1101111100001011",
40601 => "1101111100001101",
40602 => "1101111100001111",
40603 => "1101111100010001",
40604 => "1101111100010010",
40605 => "1101111100010100",
40606 => "1101111100010110",
40607 => "1101111100011000",
40608 => "1101111100011010",
40609 => "1101111100011011",
40610 => "1101111100011101",
40611 => "1101111100011111",
40612 => "1101111100100001",
40613 => "1101111100100011",
40614 => "1101111100100100",
40615 => "1101111100100110",
40616 => "1101111100101000",
40617 => "1101111100101010",
40618 => "1101111100101011",
40619 => "1101111100101101",
40620 => "1101111100101111",
40621 => "1101111100110001",
40622 => "1101111100110011",
40623 => "1101111100110100",
40624 => "1101111100110110",
40625 => "1101111100111000",
40626 => "1101111100111010",
40627 => "1101111100111100",
40628 => "1101111100111101",
40629 => "1101111100111111",
40630 => "1101111101000001",
40631 => "1101111101000011",
40632 => "1101111101000100",
40633 => "1101111101000110",
40634 => "1101111101001000",
40635 => "1101111101001010",
40636 => "1101111101001100",
40637 => "1101111101001101",
40638 => "1101111101001111",
40639 => "1101111101010001",
40640 => "1101111101010011",
40641 => "1101111101010101",
40642 => "1101111101010110",
40643 => "1101111101011000",
40644 => "1101111101011010",
40645 => "1101111101011100",
40646 => "1101111101011101",
40647 => "1101111101011111",
40648 => "1101111101100001",
40649 => "1101111101100011",
40650 => "1101111101100101",
40651 => "1101111101100110",
40652 => "1101111101101000",
40653 => "1101111101101010",
40654 => "1101111101101100",
40655 => "1101111101101101",
40656 => "1101111101101111",
40657 => "1101111101110001",
40658 => "1101111101110011",
40659 => "1101111101110101",
40660 => "1101111101110110",
40661 => "1101111101111000",
40662 => "1101111101111010",
40663 => "1101111101111100",
40664 => "1101111101111101",
40665 => "1101111101111111",
40666 => "1101111110000001",
40667 => "1101111110000011",
40668 => "1101111110000101",
40669 => "1101111110000110",
40670 => "1101111110001000",
40671 => "1101111110001010",
40672 => "1101111110001100",
40673 => "1101111110001101",
40674 => "1101111110001111",
40675 => "1101111110010001",
40676 => "1101111110010011",
40677 => "1101111110010100",
40678 => "1101111110010110",
40679 => "1101111110011000",
40680 => "1101111110011010",
40681 => "1101111110011100",
40682 => "1101111110011101",
40683 => "1101111110011111",
40684 => "1101111110100001",
40685 => "1101111110100011",
40686 => "1101111110100100",
40687 => "1101111110100110",
40688 => "1101111110101000",
40689 => "1101111110101010",
40690 => "1101111110101011",
40691 => "1101111110101101",
40692 => "1101111110101111",
40693 => "1101111110110001",
40694 => "1101111110110010",
40695 => "1101111110110100",
40696 => "1101111110110110",
40697 => "1101111110111000",
40698 => "1101111110111010",
40699 => "1101111110111011",
40700 => "1101111110111101",
40701 => "1101111110111111",
40702 => "1101111111000001",
40703 => "1101111111000010",
40704 => "1101111111000100",
40705 => "1101111111000110",
40706 => "1101111111001000",
40707 => "1101111111001001",
40708 => "1101111111001011",
40709 => "1101111111001101",
40710 => "1101111111001111",
40711 => "1101111111010000",
40712 => "1101111111010010",
40713 => "1101111111010100",
40714 => "1101111111010110",
40715 => "1101111111010111",
40716 => "1101111111011001",
40717 => "1101111111011011",
40718 => "1101111111011101",
40719 => "1101111111011110",
40720 => "1101111111100000",
40721 => "1101111111100010",
40722 => "1101111111100100",
40723 => "1101111111100110",
40724 => "1101111111100111",
40725 => "1101111111101001",
40726 => "1101111111101011",
40727 => "1101111111101101",
40728 => "1101111111101110",
40729 => "1101111111110000",
40730 => "1101111111110010",
40731 => "1101111111110100",
40732 => "1101111111110101",
40733 => "1101111111110111",
40734 => "1101111111111001",
40735 => "1101111111111011",
40736 => "1101111111111100",
40737 => "1101111111111110",
40738 => "1110000000000000",
40739 => "1110000000000010",
40740 => "1110000000000011",
40741 => "1110000000000101",
40742 => "1110000000000111",
40743 => "1110000000001001",
40744 => "1110000000001010",
40745 => "1110000000001100",
40746 => "1110000000001110",
40747 => "1110000000010000",
40748 => "1110000000010001",
40749 => "1110000000010011",
40750 => "1110000000010101",
40751 => "1110000000010111",
40752 => "1110000000011000",
40753 => "1110000000011010",
40754 => "1110000000011100",
40755 => "1110000000011110",
40756 => "1110000000011111",
40757 => "1110000000100001",
40758 => "1110000000100011",
40759 => "1110000000100100",
40760 => "1110000000100110",
40761 => "1110000000101000",
40762 => "1110000000101010",
40763 => "1110000000101011",
40764 => "1110000000101101",
40765 => "1110000000101111",
40766 => "1110000000110001",
40767 => "1110000000110010",
40768 => "1110000000110100",
40769 => "1110000000110110",
40770 => "1110000000111000",
40771 => "1110000000111001",
40772 => "1110000000111011",
40773 => "1110000000111101",
40774 => "1110000000111111",
40775 => "1110000001000000",
40776 => "1110000001000010",
40777 => "1110000001000100",
40778 => "1110000001000110",
40779 => "1110000001000111",
40780 => "1110000001001001",
40781 => "1110000001001011",
40782 => "1110000001001100",
40783 => "1110000001001110",
40784 => "1110000001010000",
40785 => "1110000001010010",
40786 => "1110000001010011",
40787 => "1110000001010101",
40788 => "1110000001010111",
40789 => "1110000001011001",
40790 => "1110000001011010",
40791 => "1110000001011100",
40792 => "1110000001011110",
40793 => "1110000001100000",
40794 => "1110000001100001",
40795 => "1110000001100011",
40796 => "1110000001100101",
40797 => "1110000001100110",
40798 => "1110000001101000",
40799 => "1110000001101010",
40800 => "1110000001101100",
40801 => "1110000001101101",
40802 => "1110000001101111",
40803 => "1110000001110001",
40804 => "1110000001110011",
40805 => "1110000001110100",
40806 => "1110000001110110",
40807 => "1110000001111000",
40808 => "1110000001111010",
40809 => "1110000001111011",
40810 => "1110000001111101",
40811 => "1110000001111111",
40812 => "1110000010000000",
40813 => "1110000010000010",
40814 => "1110000010000100",
40815 => "1110000010000110",
40816 => "1110000010000111",
40817 => "1110000010001001",
40818 => "1110000010001011",
40819 => "1110000010001101",
40820 => "1110000010001110",
40821 => "1110000010010000",
40822 => "1110000010010010",
40823 => "1110000010010011",
40824 => "1110000010010101",
40825 => "1110000010010111",
40826 => "1110000010011001",
40827 => "1110000010011010",
40828 => "1110000010011100",
40829 => "1110000010011110",
40830 => "1110000010011111",
40831 => "1110000010100001",
40832 => "1110000010100011",
40833 => "1110000010100101",
40834 => "1110000010100110",
40835 => "1110000010101000",
40836 => "1110000010101010",
40837 => "1110000010101011",
40838 => "1110000010101101",
40839 => "1110000010101111",
40840 => "1110000010110001",
40841 => "1110000010110010",
40842 => "1110000010110100",
40843 => "1110000010110110",
40844 => "1110000010111000",
40845 => "1110000010111001",
40846 => "1110000010111011",
40847 => "1110000010111101",
40848 => "1110000010111110",
40849 => "1110000011000000",
40850 => "1110000011000010",
40851 => "1110000011000100",
40852 => "1110000011000101",
40853 => "1110000011000111",
40854 => "1110000011001001",
40855 => "1110000011001010",
40856 => "1110000011001100",
40857 => "1110000011001110",
40858 => "1110000011010000",
40859 => "1110000011010001",
40860 => "1110000011010011",
40861 => "1110000011010101",
40862 => "1110000011010110",
40863 => "1110000011011000",
40864 => "1110000011011010",
40865 => "1110000011011011",
40866 => "1110000011011101",
40867 => "1110000011011111",
40868 => "1110000011100001",
40869 => "1110000011100010",
40870 => "1110000011100100",
40871 => "1110000011100110",
40872 => "1110000011100111",
40873 => "1110000011101001",
40874 => "1110000011101011",
40875 => "1110000011101101",
40876 => "1110000011101110",
40877 => "1110000011110000",
40878 => "1110000011110010",
40879 => "1110000011110011",
40880 => "1110000011110101",
40881 => "1110000011110111",
40882 => "1110000011111000",
40883 => "1110000011111010",
40884 => "1110000011111100",
40885 => "1110000011111110",
40886 => "1110000011111111",
40887 => "1110000100000001",
40888 => "1110000100000011",
40889 => "1110000100000100",
40890 => "1110000100000110",
40891 => "1110000100001000",
40892 => "1110000100001010",
40893 => "1110000100001011",
40894 => "1110000100001101",
40895 => "1110000100001111",
40896 => "1110000100010000",
40897 => "1110000100010010",
40898 => "1110000100010100",
40899 => "1110000100010101",
40900 => "1110000100010111",
40901 => "1110000100011001",
40902 => "1110000100011011",
40903 => "1110000100011100",
40904 => "1110000100011110",
40905 => "1110000100100000",
40906 => "1110000100100001",
40907 => "1110000100100011",
40908 => "1110000100100101",
40909 => "1110000100100110",
40910 => "1110000100101000",
40911 => "1110000100101010",
40912 => "1110000100101011",
40913 => "1110000100101101",
40914 => "1110000100101111",
40915 => "1110000100110001",
40916 => "1110000100110010",
40917 => "1110000100110100",
40918 => "1110000100110110",
40919 => "1110000100110111",
40920 => "1110000100111001",
40921 => "1110000100111011",
40922 => "1110000100111100",
40923 => "1110000100111110",
40924 => "1110000101000000",
40925 => "1110000101000001",
40926 => "1110000101000011",
40927 => "1110000101000101",
40928 => "1110000101000111",
40929 => "1110000101001000",
40930 => "1110000101001010",
40931 => "1110000101001100",
40932 => "1110000101001101",
40933 => "1110000101001111",
40934 => "1110000101010001",
40935 => "1110000101010010",
40936 => "1110000101010100",
40937 => "1110000101010110",
40938 => "1110000101010111",
40939 => "1110000101011001",
40940 => "1110000101011011",
40941 => "1110000101011100",
40942 => "1110000101011110",
40943 => "1110000101100000",
40944 => "1110000101100010",
40945 => "1110000101100011",
40946 => "1110000101100101",
40947 => "1110000101100111",
40948 => "1110000101101000",
40949 => "1110000101101010",
40950 => "1110000101101100",
40951 => "1110000101101101",
40952 => "1110000101101111",
40953 => "1110000101110001",
40954 => "1110000101110010",
40955 => "1110000101110100",
40956 => "1110000101110110",
40957 => "1110000101110111",
40958 => "1110000101111001",
40959 => "1110000101111011",
40960 => "1110000101111100",
40961 => "1110000101111110",
40962 => "1110000110000000",
40963 => "1110000110000010",
40964 => "1110000110000011",
40965 => "1110000110000101",
40966 => "1110000110000111",
40967 => "1110000110001000",
40968 => "1110000110001010",
40969 => "1110000110001100",
40970 => "1110000110001101",
40971 => "1110000110001111",
40972 => "1110000110010001",
40973 => "1110000110010010",
40974 => "1110000110010100",
40975 => "1110000110010110",
40976 => "1110000110010111",
40977 => "1110000110011001",
40978 => "1110000110011011",
40979 => "1110000110011100",
40980 => "1110000110011110",
40981 => "1110000110100000",
40982 => "1110000110100001",
40983 => "1110000110100011",
40984 => "1110000110100101",
40985 => "1110000110100110",
40986 => "1110000110101000",
40987 => "1110000110101010",
40988 => "1110000110101011",
40989 => "1110000110101101",
40990 => "1110000110101111",
40991 => "1110000110110000",
40992 => "1110000110110010",
40993 => "1110000110110100",
40994 => "1110000110110101",
40995 => "1110000110110111",
40996 => "1110000110111001",
40997 => "1110000110111010",
40998 => "1110000110111100",
40999 => "1110000110111110",
41000 => "1110000110111111",
41001 => "1110000111000001",
41002 => "1110000111000011",
41003 => "1110000111000100",
41004 => "1110000111000110",
41005 => "1110000111001000",
41006 => "1110000111001001",
41007 => "1110000111001011",
41008 => "1110000111001101",
41009 => "1110000111001110",
41010 => "1110000111010000",
41011 => "1110000111010010",
41012 => "1110000111010011",
41013 => "1110000111010101",
41014 => "1110000111010111",
41015 => "1110000111011000",
41016 => "1110000111011010",
41017 => "1110000111011100",
41018 => "1110000111011101",
41019 => "1110000111011111",
41020 => "1110000111100001",
41021 => "1110000111100010",
41022 => "1110000111100100",
41023 => "1110000111100110",
41024 => "1110000111100111",
41025 => "1110000111101001",
41026 => "1110000111101011",
41027 => "1110000111101100",
41028 => "1110000111101110",
41029 => "1110000111110000",
41030 => "1110000111110001",
41031 => "1110000111110011",
41032 => "1110000111110101",
41033 => "1110000111110110",
41034 => "1110000111111000",
41035 => "1110000111111010",
41036 => "1110000111111011",
41037 => "1110000111111101",
41038 => "1110000111111111",
41039 => "1110001000000000",
41040 => "1110001000000010",
41041 => "1110001000000100",
41042 => "1110001000000101",
41043 => "1110001000000111",
41044 => "1110001000001000",
41045 => "1110001000001010",
41046 => "1110001000001100",
41047 => "1110001000001101",
41048 => "1110001000001111",
41049 => "1110001000010001",
41050 => "1110001000010010",
41051 => "1110001000010100",
41052 => "1110001000010110",
41053 => "1110001000010111",
41054 => "1110001000011001",
41055 => "1110001000011011",
41056 => "1110001000011100",
41057 => "1110001000011110",
41058 => "1110001000100000",
41059 => "1110001000100001",
41060 => "1110001000100011",
41061 => "1110001000100101",
41062 => "1110001000100110",
41063 => "1110001000101000",
41064 => "1110001000101001",
41065 => "1110001000101011",
41066 => "1110001000101101",
41067 => "1110001000101110",
41068 => "1110001000110000",
41069 => "1110001000110010",
41070 => "1110001000110011",
41071 => "1110001000110101",
41072 => "1110001000110111",
41073 => "1110001000111000",
41074 => "1110001000111010",
41075 => "1110001000111100",
41076 => "1110001000111101",
41077 => "1110001000111111",
41078 => "1110001001000001",
41079 => "1110001001000010",
41080 => "1110001001000100",
41081 => "1110001001000101",
41082 => "1110001001000111",
41083 => "1110001001001001",
41084 => "1110001001001010",
41085 => "1110001001001100",
41086 => "1110001001001110",
41087 => "1110001001001111",
41088 => "1110001001010001",
41089 => "1110001001010011",
41090 => "1110001001010100",
41091 => "1110001001010110",
41092 => "1110001001010111",
41093 => "1110001001011001",
41094 => "1110001001011011",
41095 => "1110001001011100",
41096 => "1110001001011110",
41097 => "1110001001100000",
41098 => "1110001001100001",
41099 => "1110001001100011",
41100 => "1110001001100101",
41101 => "1110001001100110",
41102 => "1110001001101000",
41103 => "1110001001101001",
41104 => "1110001001101011",
41105 => "1110001001101101",
41106 => "1110001001101110",
41107 => "1110001001110000",
41108 => "1110001001110010",
41109 => "1110001001110011",
41110 => "1110001001110101",
41111 => "1110001001110111",
41112 => "1110001001111000",
41113 => "1110001001111010",
41114 => "1110001001111011",
41115 => "1110001001111101",
41116 => "1110001001111111",
41117 => "1110001010000000",
41118 => "1110001010000010",
41119 => "1110001010000100",
41120 => "1110001010000101",
41121 => "1110001010000111",
41122 => "1110001010001001",
41123 => "1110001010001010",
41124 => "1110001010001100",
41125 => "1110001010001101",
41126 => "1110001010001111",
41127 => "1110001010010001",
41128 => "1110001010010010",
41129 => "1110001010010100",
41130 => "1110001010010110",
41131 => "1110001010010111",
41132 => "1110001010011001",
41133 => "1110001010011010",
41134 => "1110001010011100",
41135 => "1110001010011110",
41136 => "1110001010011111",
41137 => "1110001010100001",
41138 => "1110001010100011",
41139 => "1110001010100100",
41140 => "1110001010100110",
41141 => "1110001010100111",
41142 => "1110001010101001",
41143 => "1110001010101011",
41144 => "1110001010101100",
41145 => "1110001010101110",
41146 => "1110001010110000",
41147 => "1110001010110001",
41148 => "1110001010110011",
41149 => "1110001010110100",
41150 => "1110001010110110",
41151 => "1110001010111000",
41152 => "1110001010111001",
41153 => "1110001010111011",
41154 => "1110001010111101",
41155 => "1110001010111110",
41156 => "1110001011000000",
41157 => "1110001011000001",
41158 => "1110001011000011",
41159 => "1110001011000101",
41160 => "1110001011000110",
41161 => "1110001011001000",
41162 => "1110001011001001",
41163 => "1110001011001011",
41164 => "1110001011001101",
41165 => "1110001011001110",
41166 => "1110001011010000",
41167 => "1110001011010010",
41168 => "1110001011010011",
41169 => "1110001011010101",
41170 => "1110001011010110",
41171 => "1110001011011000",
41172 => "1110001011011010",
41173 => "1110001011011011",
41174 => "1110001011011101",
41175 => "1110001011011110",
41176 => "1110001011100000",
41177 => "1110001011100010",
41178 => "1110001011100011",
41179 => "1110001011100101",
41180 => "1110001011100111",
41181 => "1110001011101000",
41182 => "1110001011101010",
41183 => "1110001011101011",
41184 => "1110001011101101",
41185 => "1110001011101111",
41186 => "1110001011110000",
41187 => "1110001011110010",
41188 => "1110001011110011",
41189 => "1110001011110101",
41190 => "1110001011110111",
41191 => "1110001011111000",
41192 => "1110001011111010",
41193 => "1110001011111011",
41194 => "1110001011111101",
41195 => "1110001011111111",
41196 => "1110001100000000",
41197 => "1110001100000010",
41198 => "1110001100000011",
41199 => "1110001100000101",
41200 => "1110001100000111",
41201 => "1110001100001000",
41202 => "1110001100001010",
41203 => "1110001100001100",
41204 => "1110001100001101",
41205 => "1110001100001111",
41206 => "1110001100010000",
41207 => "1110001100010010",
41208 => "1110001100010100",
41209 => "1110001100010101",
41210 => "1110001100010111",
41211 => "1110001100011000",
41212 => "1110001100011010",
41213 => "1110001100011100",
41214 => "1110001100011101",
41215 => "1110001100011111",
41216 => "1110001100100000",
41217 => "1110001100100010",
41218 => "1110001100100100",
41219 => "1110001100100101",
41220 => "1110001100100111",
41221 => "1110001100101000",
41222 => "1110001100101010",
41223 => "1110001100101100",
41224 => "1110001100101101",
41225 => "1110001100101111",
41226 => "1110001100110000",
41227 => "1110001100110010",
41228 => "1110001100110100",
41229 => "1110001100110101",
41230 => "1110001100110111",
41231 => "1110001100111000",
41232 => "1110001100111010",
41233 => "1110001100111100",
41234 => "1110001100111101",
41235 => "1110001100111111",
41236 => "1110001101000000",
41237 => "1110001101000010",
41238 => "1110001101000011",
41239 => "1110001101000101",
41240 => "1110001101000111",
41241 => "1110001101001000",
41242 => "1110001101001010",
41243 => "1110001101001011",
41244 => "1110001101001101",
41245 => "1110001101001111",
41246 => "1110001101010000",
41247 => "1110001101010010",
41248 => "1110001101010011",
41249 => "1110001101010101",
41250 => "1110001101010111",
41251 => "1110001101011000",
41252 => "1110001101011010",
41253 => "1110001101011011",
41254 => "1110001101011101",
41255 => "1110001101011111",
41256 => "1110001101100000",
41257 => "1110001101100010",
41258 => "1110001101100011",
41259 => "1110001101100101",
41260 => "1110001101100110",
41261 => "1110001101101000",
41262 => "1110001101101010",
41263 => "1110001101101011",
41264 => "1110001101101101",
41265 => "1110001101101110",
41266 => "1110001101110000",
41267 => "1110001101110010",
41268 => "1110001101110011",
41269 => "1110001101110101",
41270 => "1110001101110110",
41271 => "1110001101111000",
41272 => "1110001101111010",
41273 => "1110001101111011",
41274 => "1110001101111101",
41275 => "1110001101111110",
41276 => "1110001110000000",
41277 => "1110001110000001",
41278 => "1110001110000011",
41279 => "1110001110000101",
41280 => "1110001110000110",
41281 => "1110001110001000",
41282 => "1110001110001001",
41283 => "1110001110001011",
41284 => "1110001110001101",
41285 => "1110001110001110",
41286 => "1110001110010000",
41287 => "1110001110010001",
41288 => "1110001110010011",
41289 => "1110001110010100",
41290 => "1110001110010110",
41291 => "1110001110011000",
41292 => "1110001110011001",
41293 => "1110001110011011",
41294 => "1110001110011100",
41295 => "1110001110011110",
41296 => "1110001110011111",
41297 => "1110001110100001",
41298 => "1110001110100011",
41299 => "1110001110100100",
41300 => "1110001110100110",
41301 => "1110001110100111",
41302 => "1110001110101001",
41303 => "1110001110101010",
41304 => "1110001110101100",
41305 => "1110001110101110",
41306 => "1110001110101111",
41307 => "1110001110110001",
41308 => "1110001110110010",
41309 => "1110001110110100",
41310 => "1110001110110110",
41311 => "1110001110110111",
41312 => "1110001110111001",
41313 => "1110001110111010",
41314 => "1110001110111100",
41315 => "1110001110111101",
41316 => "1110001110111111",
41317 => "1110001111000001",
41318 => "1110001111000010",
41319 => "1110001111000100",
41320 => "1110001111000101",
41321 => "1110001111000111",
41322 => "1110001111001000",
41323 => "1110001111001010",
41324 => "1110001111001011",
41325 => "1110001111001101",
41326 => "1110001111001111",
41327 => "1110001111010000",
41328 => "1110001111010010",
41329 => "1110001111010011",
41330 => "1110001111010101",
41331 => "1110001111010110",
41332 => "1110001111011000",
41333 => "1110001111011010",
41334 => "1110001111011011",
41335 => "1110001111011101",
41336 => "1110001111011110",
41337 => "1110001111100000",
41338 => "1110001111100001",
41339 => "1110001111100011",
41340 => "1110001111100101",
41341 => "1110001111100110",
41342 => "1110001111101000",
41343 => "1110001111101001",
41344 => "1110001111101011",
41345 => "1110001111101100",
41346 => "1110001111101110",
41347 => "1110001111101111",
41348 => "1110001111110001",
41349 => "1110001111110011",
41350 => "1110001111110100",
41351 => "1110001111110110",
41352 => "1110001111110111",
41353 => "1110001111111001",
41354 => "1110001111111010",
41355 => "1110001111111100",
41356 => "1110001111111110",
41357 => "1110001111111111",
41358 => "1110010000000001",
41359 => "1110010000000010",
41360 => "1110010000000100",
41361 => "1110010000000101",
41362 => "1110010000000111",
41363 => "1110010000001000",
41364 => "1110010000001010",
41365 => "1110010000001100",
41366 => "1110010000001101",
41367 => "1110010000001111",
41368 => "1110010000010000",
41369 => "1110010000010010",
41370 => "1110010000010011",
41371 => "1110010000010101",
41372 => "1110010000010110",
41373 => "1110010000011000",
41374 => "1110010000011010",
41375 => "1110010000011011",
41376 => "1110010000011101",
41377 => "1110010000011110",
41378 => "1110010000100000",
41379 => "1110010000100001",
41380 => "1110010000100011",
41381 => "1110010000100100",
41382 => "1110010000100110",
41383 => "1110010000101000",
41384 => "1110010000101001",
41385 => "1110010000101011",
41386 => "1110010000101100",
41387 => "1110010000101110",
41388 => "1110010000101111",
41389 => "1110010000110001",
41390 => "1110010000110010",
41391 => "1110010000110100",
41392 => "1110010000110101",
41393 => "1110010000110111",
41394 => "1110010000111001",
41395 => "1110010000111010",
41396 => "1110010000111100",
41397 => "1110010000111101",
41398 => "1110010000111111",
41399 => "1110010001000000",
41400 => "1110010001000010",
41401 => "1110010001000011",
41402 => "1110010001000101",
41403 => "1110010001000110",
41404 => "1110010001001000",
41405 => "1110010001001010",
41406 => "1110010001001011",
41407 => "1110010001001101",
41408 => "1110010001001110",
41409 => "1110010001010000",
41410 => "1110010001010001",
41411 => "1110010001010011",
41412 => "1110010001010100",
41413 => "1110010001010110",
41414 => "1110010001010111",
41415 => "1110010001011001",
41416 => "1110010001011011",
41417 => "1110010001011100",
41418 => "1110010001011110",
41419 => "1110010001011111",
41420 => "1110010001100001",
41421 => "1110010001100010",
41422 => "1110010001100100",
41423 => "1110010001100101",
41424 => "1110010001100111",
41425 => "1110010001101000",
41426 => "1110010001101010",
41427 => "1110010001101011",
41428 => "1110010001101101",
41429 => "1110010001101111",
41430 => "1110010001110000",
41431 => "1110010001110010",
41432 => "1110010001110011",
41433 => "1110010001110101",
41434 => "1110010001110110",
41435 => "1110010001111000",
41436 => "1110010001111001",
41437 => "1110010001111011",
41438 => "1110010001111100",
41439 => "1110010001111110",
41440 => "1110010001111111",
41441 => "1110010010000001",
41442 => "1110010010000011",
41443 => "1110010010000100",
41444 => "1110010010000110",
41445 => "1110010010000111",
41446 => "1110010010001001",
41447 => "1110010010001010",
41448 => "1110010010001100",
41449 => "1110010010001101",
41450 => "1110010010001111",
41451 => "1110010010010000",
41452 => "1110010010010010",
41453 => "1110010010010011",
41454 => "1110010010010101",
41455 => "1110010010010110",
41456 => "1110010010011000",
41457 => "1110010010011001",
41458 => "1110010010011011",
41459 => "1110010010011101",
41460 => "1110010010011110",
41461 => "1110010010100000",
41462 => "1110010010100001",
41463 => "1110010010100011",
41464 => "1110010010100100",
41465 => "1110010010100110",
41466 => "1110010010100111",
41467 => "1110010010101001",
41468 => "1110010010101010",
41469 => "1110010010101100",
41470 => "1110010010101101",
41471 => "1110010010101111",
41472 => "1110010010110000",
41473 => "1110010010110010",
41474 => "1110010010110011",
41475 => "1110010010110101",
41476 => "1110010010110110",
41477 => "1110010010111000",
41478 => "1110010010111010",
41479 => "1110010010111011",
41480 => "1110010010111101",
41481 => "1110010010111110",
41482 => "1110010011000000",
41483 => "1110010011000001",
41484 => "1110010011000011",
41485 => "1110010011000100",
41486 => "1110010011000110",
41487 => "1110010011000111",
41488 => "1110010011001001",
41489 => "1110010011001010",
41490 => "1110010011001100",
41491 => "1110010011001101",
41492 => "1110010011001111",
41493 => "1110010011010000",
41494 => "1110010011010010",
41495 => "1110010011010011",
41496 => "1110010011010101",
41497 => "1110010011010110",
41498 => "1110010011011000",
41499 => "1110010011011001",
41500 => "1110010011011011",
41501 => "1110010011011100",
41502 => "1110010011011110",
41503 => "1110010011100000",
41504 => "1110010011100001",
41505 => "1110010011100011",
41506 => "1110010011100100",
41507 => "1110010011100110",
41508 => "1110010011100111",
41509 => "1110010011101001",
41510 => "1110010011101010",
41511 => "1110010011101100",
41512 => "1110010011101101",
41513 => "1110010011101111",
41514 => "1110010011110000",
41515 => "1110010011110010",
41516 => "1110010011110011",
41517 => "1110010011110101",
41518 => "1110010011110110",
41519 => "1110010011111000",
41520 => "1110010011111001",
41521 => "1110010011111011",
41522 => "1110010011111100",
41523 => "1110010011111110",
41524 => "1110010011111111",
41525 => "1110010100000001",
41526 => "1110010100000010",
41527 => "1110010100000100",
41528 => "1110010100000101",
41529 => "1110010100000111",
41530 => "1110010100001000",
41531 => "1110010100001010",
41532 => "1110010100001011",
41533 => "1110010100001101",
41534 => "1110010100001110",
41535 => "1110010100010000",
41536 => "1110010100010001",
41537 => "1110010100010011",
41538 => "1110010100010100",
41539 => "1110010100010110",
41540 => "1110010100010111",
41541 => "1110010100011001",
41542 => "1110010100011010",
41543 => "1110010100011100",
41544 => "1110010100011101",
41545 => "1110010100011111",
41546 => "1110010100100000",
41547 => "1110010100100010",
41548 => "1110010100100011",
41549 => "1110010100100101",
41550 => "1110010100100110",
41551 => "1110010100101000",
41552 => "1110010100101001",
41553 => "1110010100101011",
41554 => "1110010100101100",
41555 => "1110010100101110",
41556 => "1110010100101111",
41557 => "1110010100110001",
41558 => "1110010100110010",
41559 => "1110010100110100",
41560 => "1110010100110101",
41561 => "1110010100110111",
41562 => "1110010100111000",
41563 => "1110010100111010",
41564 => "1110010100111011",
41565 => "1110010100111101",
41566 => "1110010100111110",
41567 => "1110010101000000",
41568 => "1110010101000001",
41569 => "1110010101000011",
41570 => "1110010101000100",
41571 => "1110010101000110",
41572 => "1110010101000111",
41573 => "1110010101001001",
41574 => "1110010101001010",
41575 => "1110010101001100",
41576 => "1110010101001101",
41577 => "1110010101001111",
41578 => "1110010101010000",
41579 => "1110010101010010",
41580 => "1110010101010011",
41581 => "1110010101010101",
41582 => "1110010101010110",
41583 => "1110010101011000",
41584 => "1110010101011001",
41585 => "1110010101011011",
41586 => "1110010101011100",
41587 => "1110010101011110",
41588 => "1110010101011111",
41589 => "1110010101100001",
41590 => "1110010101100010",
41591 => "1110010101100100",
41592 => "1110010101100101",
41593 => "1110010101100111",
41594 => "1110010101101000",
41595 => "1110010101101010",
41596 => "1110010101101011",
41597 => "1110010101101101",
41598 => "1110010101101110",
41599 => "1110010101110000",
41600 => "1110010101110001",
41601 => "1110010101110011",
41602 => "1110010101110100",
41603 => "1110010101110110",
41604 => "1110010101110111",
41605 => "1110010101111001",
41606 => "1110010101111010",
41607 => "1110010101111100",
41608 => "1110010101111101",
41609 => "1110010101111111",
41610 => "1110010110000000",
41611 => "1110010110000010",
41612 => "1110010110000011",
41613 => "1110010110000100",
41614 => "1110010110000110",
41615 => "1110010110000111",
41616 => "1110010110001001",
41617 => "1110010110001010",
41618 => "1110010110001100",
41619 => "1110010110001101",
41620 => "1110010110001111",
41621 => "1110010110010000",
41622 => "1110010110010010",
41623 => "1110010110010011",
41624 => "1110010110010101",
41625 => "1110010110010110",
41626 => "1110010110011000",
41627 => "1110010110011001",
41628 => "1110010110011011",
41629 => "1110010110011100",
41630 => "1110010110011110",
41631 => "1110010110011111",
41632 => "1110010110100001",
41633 => "1110010110100010",
41634 => "1110010110100100",
41635 => "1110010110100101",
41636 => "1110010110100111",
41637 => "1110010110101000",
41638 => "1110010110101001",
41639 => "1110010110101011",
41640 => "1110010110101100",
41641 => "1110010110101110",
41642 => "1110010110101111",
41643 => "1110010110110001",
41644 => "1110010110110010",
41645 => "1110010110110100",
41646 => "1110010110110101",
41647 => "1110010110110111",
41648 => "1110010110111000",
41649 => "1110010110111010",
41650 => "1110010110111011",
41651 => "1110010110111101",
41652 => "1110010110111110",
41653 => "1110010111000000",
41654 => "1110010111000001",
41655 => "1110010111000011",
41656 => "1110010111000100",
41657 => "1110010111000110",
41658 => "1110010111000111",
41659 => "1110010111001000",
41660 => "1110010111001010",
41661 => "1110010111001011",
41662 => "1110010111001101",
41663 => "1110010111001110",
41664 => "1110010111010000",
41665 => "1110010111010001",
41666 => "1110010111010011",
41667 => "1110010111010100",
41668 => "1110010111010110",
41669 => "1110010111010111",
41670 => "1110010111011001",
41671 => "1110010111011010",
41672 => "1110010111011100",
41673 => "1110010111011101",
41674 => "1110010111011110",
41675 => "1110010111100000",
41676 => "1110010111100001",
41677 => "1110010111100011",
41678 => "1110010111100100",
41679 => "1110010111100110",
41680 => "1110010111100111",
41681 => "1110010111101001",
41682 => "1110010111101010",
41683 => "1110010111101100",
41684 => "1110010111101101",
41685 => "1110010111101111",
41686 => "1110010111110000",
41687 => "1110010111110010",
41688 => "1110010111110011",
41689 => "1110010111110100",
41690 => "1110010111110110",
41691 => "1110010111110111",
41692 => "1110010111111001",
41693 => "1110010111111010",
41694 => "1110010111111100",
41695 => "1110010111111101",
41696 => "1110010111111111",
41697 => "1110011000000000",
41698 => "1110011000000010",
41699 => "1110011000000011",
41700 => "1110011000000101",
41701 => "1110011000000110",
41702 => "1110011000000111",
41703 => "1110011000001001",
41704 => "1110011000001010",
41705 => "1110011000001100",
41706 => "1110011000001101",
41707 => "1110011000001111",
41708 => "1110011000010000",
41709 => "1110011000010010",
41710 => "1110011000010011",
41711 => "1110011000010101",
41712 => "1110011000010110",
41713 => "1110011000010111",
41714 => "1110011000011001",
41715 => "1110011000011010",
41716 => "1110011000011100",
41717 => "1110011000011101",
41718 => "1110011000011111",
41719 => "1110011000100000",
41720 => "1110011000100010",
41721 => "1110011000100011",
41722 => "1110011000100101",
41723 => "1110011000100110",
41724 => "1110011000100111",
41725 => "1110011000101001",
41726 => "1110011000101010",
41727 => "1110011000101100",
41728 => "1110011000101101",
41729 => "1110011000101111",
41730 => "1110011000110000",
41731 => "1110011000110010",
41732 => "1110011000110011",
41733 => "1110011000110100",
41734 => "1110011000110110",
41735 => "1110011000110111",
41736 => "1110011000111001",
41737 => "1110011000111010",
41738 => "1110011000111100",
41739 => "1110011000111101",
41740 => "1110011000111111",
41741 => "1110011001000000",
41742 => "1110011001000010",
41743 => "1110011001000011",
41744 => "1110011001000100",
41745 => "1110011001000110",
41746 => "1110011001000111",
41747 => "1110011001001001",
41748 => "1110011001001010",
41749 => "1110011001001100",
41750 => "1110011001001101",
41751 => "1110011001001111",
41752 => "1110011001010000",
41753 => "1110011001010001",
41754 => "1110011001010011",
41755 => "1110011001010100",
41756 => "1110011001010110",
41757 => "1110011001010111",
41758 => "1110011001011001",
41759 => "1110011001011010",
41760 => "1110011001011100",
41761 => "1110011001011101",
41762 => "1110011001011110",
41763 => "1110011001100000",
41764 => "1110011001100001",
41765 => "1110011001100011",
41766 => "1110011001100100",
41767 => "1110011001100110",
41768 => "1110011001100111",
41769 => "1110011001101000",
41770 => "1110011001101010",
41771 => "1110011001101011",
41772 => "1110011001101101",
41773 => "1110011001101110",
41774 => "1110011001110000",
41775 => "1110011001110001",
41776 => "1110011001110011",
41777 => "1110011001110100",
41778 => "1110011001110101",
41779 => "1110011001110111",
41780 => "1110011001111000",
41781 => "1110011001111010",
41782 => "1110011001111011",
41783 => "1110011001111101",
41784 => "1110011001111110",
41785 => "1110011001111111",
41786 => "1110011010000001",
41787 => "1110011010000010",
41788 => "1110011010000100",
41789 => "1110011010000101",
41790 => "1110011010000111",
41791 => "1110011010001000",
41792 => "1110011010001010",
41793 => "1110011010001011",
41794 => "1110011010001100",
41795 => "1110011010001110",
41796 => "1110011010001111",
41797 => "1110011010010001",
41798 => "1110011010010010",
41799 => "1110011010010100",
41800 => "1110011010010101",
41801 => "1110011010010110",
41802 => "1110011010011000",
41803 => "1110011010011001",
41804 => "1110011010011011",
41805 => "1110011010011100",
41806 => "1110011010011110",
41807 => "1110011010011111",
41808 => "1110011010100000",
41809 => "1110011010100010",
41810 => "1110011010100011",
41811 => "1110011010100101",
41812 => "1110011010100110",
41813 => "1110011010101000",
41814 => "1110011010101001",
41815 => "1110011010101010",
41816 => "1110011010101100",
41817 => "1110011010101101",
41818 => "1110011010101111",
41819 => "1110011010110000",
41820 => "1110011010110010",
41821 => "1110011010110011",
41822 => "1110011010110100",
41823 => "1110011010110110",
41824 => "1110011010110111",
41825 => "1110011010111001",
41826 => "1110011010111010",
41827 => "1110011010111100",
41828 => "1110011010111101",
41829 => "1110011010111110",
41830 => "1110011011000000",
41831 => "1110011011000001",
41832 => "1110011011000011",
41833 => "1110011011000100",
41834 => "1110011011000101",
41835 => "1110011011000111",
41836 => "1110011011001000",
41837 => "1110011011001010",
41838 => "1110011011001011",
41839 => "1110011011001101",
41840 => "1110011011001110",
41841 => "1110011011001111",
41842 => "1110011011010001",
41843 => "1110011011010010",
41844 => "1110011011010100",
41845 => "1110011011010101",
41846 => "1110011011010111",
41847 => "1110011011011000",
41848 => "1110011011011001",
41849 => "1110011011011011",
41850 => "1110011011011100",
41851 => "1110011011011110",
41852 => "1110011011011111",
41853 => "1110011011100000",
41854 => "1110011011100010",
41855 => "1110011011100011",
41856 => "1110011011100101",
41857 => "1110011011100110",
41858 => "1110011011101000",
41859 => "1110011011101001",
41860 => "1110011011101010",
41861 => "1110011011101100",
41862 => "1110011011101101",
41863 => "1110011011101111",
41864 => "1110011011110000",
41865 => "1110011011110001",
41866 => "1110011011110011",
41867 => "1110011011110100",
41868 => "1110011011110110",
41869 => "1110011011110111",
41870 => "1110011011111000",
41871 => "1110011011111010",
41872 => "1110011011111011",
41873 => "1110011011111101",
41874 => "1110011011111110",
41875 => "1110011100000000",
41876 => "1110011100000001",
41877 => "1110011100000010",
41878 => "1110011100000100",
41879 => "1110011100000101",
41880 => "1110011100000111",
41881 => "1110011100001000",
41882 => "1110011100001001",
41883 => "1110011100001011",
41884 => "1110011100001100",
41885 => "1110011100001110",
41886 => "1110011100001111",
41887 => "1110011100010000",
41888 => "1110011100010010",
41889 => "1110011100010011",
41890 => "1110011100010101",
41891 => "1110011100010110",
41892 => "1110011100010111",
41893 => "1110011100011001",
41894 => "1110011100011010",
41895 => "1110011100011100",
41896 => "1110011100011101",
41897 => "1110011100011110",
41898 => "1110011100100000",
41899 => "1110011100100001",
41900 => "1110011100100011",
41901 => "1110011100100100",
41902 => "1110011100100101",
41903 => "1110011100100111",
41904 => "1110011100101000",
41905 => "1110011100101010",
41906 => "1110011100101011",
41907 => "1110011100101100",
41908 => "1110011100101110",
41909 => "1110011100101111",
41910 => "1110011100110001",
41911 => "1110011100110010",
41912 => "1110011100110011",
41913 => "1110011100110101",
41914 => "1110011100110110",
41915 => "1110011100111000",
41916 => "1110011100111001",
41917 => "1110011100111010",
41918 => "1110011100111100",
41919 => "1110011100111101",
41920 => "1110011100111111",
41921 => "1110011101000000",
41922 => "1110011101000001",
41923 => "1110011101000011",
41924 => "1110011101000100",
41925 => "1110011101000110",
41926 => "1110011101000111",
41927 => "1110011101001000",
41928 => "1110011101001010",
41929 => "1110011101001011",
41930 => "1110011101001101",
41931 => "1110011101001110",
41932 => "1110011101001111",
41933 => "1110011101010001",
41934 => "1110011101010010",
41935 => "1110011101010100",
41936 => "1110011101010101",
41937 => "1110011101010110",
41938 => "1110011101011000",
41939 => "1110011101011001",
41940 => "1110011101011011",
41941 => "1110011101011100",
41942 => "1110011101011101",
41943 => "1110011101011111",
41944 => "1110011101100000",
41945 => "1110011101100010",
41946 => "1110011101100011",
41947 => "1110011101100100",
41948 => "1110011101100110",
41949 => "1110011101100111",
41950 => "1110011101101000",
41951 => "1110011101101010",
41952 => "1110011101101011",
41953 => "1110011101101101",
41954 => "1110011101101110",
41955 => "1110011101101111",
41956 => "1110011101110001",
41957 => "1110011101110010",
41958 => "1110011101110100",
41959 => "1110011101110101",
41960 => "1110011101110110",
41961 => "1110011101111000",
41962 => "1110011101111001",
41963 => "1110011101111011",
41964 => "1110011101111100",
41965 => "1110011101111101",
41966 => "1110011101111111",
41967 => "1110011110000000",
41968 => "1110011110000001",
41969 => "1110011110000011",
41970 => "1110011110000100",
41971 => "1110011110000110",
41972 => "1110011110000111",
41973 => "1110011110001000",
41974 => "1110011110001010",
41975 => "1110011110001011",
41976 => "1110011110001101",
41977 => "1110011110001110",
41978 => "1110011110001111",
41979 => "1110011110010001",
41980 => "1110011110010010",
41981 => "1110011110010011",
41982 => "1110011110010101",
41983 => "1110011110010110",
41984 => "1110011110011000",
41985 => "1110011110011001",
41986 => "1110011110011010",
41987 => "1110011110011100",
41988 => "1110011110011101",
41989 => "1110011110011110",
41990 => "1110011110100000",
41991 => "1110011110100001",
41992 => "1110011110100011",
41993 => "1110011110100100",
41994 => "1110011110100101",
41995 => "1110011110100111",
41996 => "1110011110101000",
41997 => "1110011110101001",
41998 => "1110011110101011",
41999 => "1110011110101100",
42000 => "1110011110101110",
42001 => "1110011110101111",
42002 => "1110011110110000",
42003 => "1110011110110010",
42004 => "1110011110110011",
42005 => "1110011110110100",
42006 => "1110011110110110",
42007 => "1110011110110111",
42008 => "1110011110111001",
42009 => "1110011110111010",
42010 => "1110011110111011",
42011 => "1110011110111101",
42012 => "1110011110111110",
42013 => "1110011110111111",
42014 => "1110011111000001",
42015 => "1110011111000010",
42016 => "1110011111000100",
42017 => "1110011111000101",
42018 => "1110011111000110",
42019 => "1110011111001000",
42020 => "1110011111001001",
42021 => "1110011111001010",
42022 => "1110011111001100",
42023 => "1110011111001101",
42024 => "1110011111001111",
42025 => "1110011111010000",
42026 => "1110011111010001",
42027 => "1110011111010011",
42028 => "1110011111010100",
42029 => "1110011111010101",
42030 => "1110011111010111",
42031 => "1110011111011000",
42032 => "1110011111011001",
42033 => "1110011111011011",
42034 => "1110011111011100",
42035 => "1110011111011110",
42036 => "1110011111011111",
42037 => "1110011111100000",
42038 => "1110011111100010",
42039 => "1110011111100011",
42040 => "1110011111100100",
42041 => "1110011111100110",
42042 => "1110011111100111",
42043 => "1110011111101001",
42044 => "1110011111101010",
42045 => "1110011111101011",
42046 => "1110011111101101",
42047 => "1110011111101110",
42048 => "1110011111101111",
42049 => "1110011111110001",
42050 => "1110011111110010",
42051 => "1110011111110011",
42052 => "1110011111110101",
42053 => "1110011111110110",
42054 => "1110011111110111",
42055 => "1110011111111001",
42056 => "1110011111111010",
42057 => "1110011111111100",
42058 => "1110011111111101",
42059 => "1110011111111110",
42060 => "1110100000000000",
42061 => "1110100000000001",
42062 => "1110100000000010",
42063 => "1110100000000100",
42064 => "1110100000000101",
42065 => "1110100000000110",
42066 => "1110100000001000",
42067 => "1110100000001001",
42068 => "1110100000001011",
42069 => "1110100000001100",
42070 => "1110100000001101",
42071 => "1110100000001111",
42072 => "1110100000010000",
42073 => "1110100000010001",
42074 => "1110100000010011",
42075 => "1110100000010100",
42076 => "1110100000010101",
42077 => "1110100000010111",
42078 => "1110100000011000",
42079 => "1110100000011001",
42080 => "1110100000011011",
42081 => "1110100000011100",
42082 => "1110100000011101",
42083 => "1110100000011111",
42084 => "1110100000100000",
42085 => "1110100000100010",
42086 => "1110100000100011",
42087 => "1110100000100100",
42088 => "1110100000100110",
42089 => "1110100000100111",
42090 => "1110100000101000",
42091 => "1110100000101010",
42092 => "1110100000101011",
42093 => "1110100000101100",
42094 => "1110100000101110",
42095 => "1110100000101111",
42096 => "1110100000110000",
42097 => "1110100000110010",
42098 => "1110100000110011",
42099 => "1110100000110100",
42100 => "1110100000110110",
42101 => "1110100000110111",
42102 => "1110100000111001",
42103 => "1110100000111010",
42104 => "1110100000111011",
42105 => "1110100000111101",
42106 => "1110100000111110",
42107 => "1110100000111111",
42108 => "1110100001000001",
42109 => "1110100001000010",
42110 => "1110100001000011",
42111 => "1110100001000101",
42112 => "1110100001000110",
42113 => "1110100001000111",
42114 => "1110100001001001",
42115 => "1110100001001010",
42116 => "1110100001001011",
42117 => "1110100001001101",
42118 => "1110100001001110",
42119 => "1110100001001111",
42120 => "1110100001010001",
42121 => "1110100001010010",
42122 => "1110100001010011",
42123 => "1110100001010101",
42124 => "1110100001010110",
42125 => "1110100001010111",
42126 => "1110100001011001",
42127 => "1110100001011010",
42128 => "1110100001011011",
42129 => "1110100001011101",
42130 => "1110100001011110",
42131 => "1110100001011111",
42132 => "1110100001100001",
42133 => "1110100001100010",
42134 => "1110100001100100",
42135 => "1110100001100101",
42136 => "1110100001100110",
42137 => "1110100001101000",
42138 => "1110100001101001",
42139 => "1110100001101010",
42140 => "1110100001101100",
42141 => "1110100001101101",
42142 => "1110100001101110",
42143 => "1110100001110000",
42144 => "1110100001110001",
42145 => "1110100001110010",
42146 => "1110100001110100",
42147 => "1110100001110101",
42148 => "1110100001110110",
42149 => "1110100001111000",
42150 => "1110100001111001",
42151 => "1110100001111010",
42152 => "1110100001111100",
42153 => "1110100001111101",
42154 => "1110100001111110",
42155 => "1110100010000000",
42156 => "1110100010000001",
42157 => "1110100010000010",
42158 => "1110100010000100",
42159 => "1110100010000101",
42160 => "1110100010000110",
42161 => "1110100010001000",
42162 => "1110100010001001",
42163 => "1110100010001010",
42164 => "1110100010001100",
42165 => "1110100010001101",
42166 => "1110100010001110",
42167 => "1110100010010000",
42168 => "1110100010010001",
42169 => "1110100010010010",
42170 => "1110100010010100",
42171 => "1110100010010101",
42172 => "1110100010010110",
42173 => "1110100010011000",
42174 => "1110100010011001",
42175 => "1110100010011010",
42176 => "1110100010011100",
42177 => "1110100010011101",
42178 => "1110100010011110",
42179 => "1110100010100000",
42180 => "1110100010100001",
42181 => "1110100010100010",
42182 => "1110100010100100",
42183 => "1110100010100101",
42184 => "1110100010100110",
42185 => "1110100010100111",
42186 => "1110100010101001",
42187 => "1110100010101010",
42188 => "1110100010101011",
42189 => "1110100010101101",
42190 => "1110100010101110",
42191 => "1110100010101111",
42192 => "1110100010110001",
42193 => "1110100010110010",
42194 => "1110100010110011",
42195 => "1110100010110101",
42196 => "1110100010110110",
42197 => "1110100010110111",
42198 => "1110100010111001",
42199 => "1110100010111010",
42200 => "1110100010111011",
42201 => "1110100010111101",
42202 => "1110100010111110",
42203 => "1110100010111111",
42204 => "1110100011000001",
42205 => "1110100011000010",
42206 => "1110100011000011",
42207 => "1110100011000101",
42208 => "1110100011000110",
42209 => "1110100011000111",
42210 => "1110100011001001",
42211 => "1110100011001010",
42212 => "1110100011001011",
42213 => "1110100011001101",
42214 => "1110100011001110",
42215 => "1110100011001111",
42216 => "1110100011010000",
42217 => "1110100011010010",
42218 => "1110100011010011",
42219 => "1110100011010100",
42220 => "1110100011010110",
42221 => "1110100011010111",
42222 => "1110100011011000",
42223 => "1110100011011010",
42224 => "1110100011011011",
42225 => "1110100011011100",
42226 => "1110100011011110",
42227 => "1110100011011111",
42228 => "1110100011100000",
42229 => "1110100011100010",
42230 => "1110100011100011",
42231 => "1110100011100100",
42232 => "1110100011100110",
42233 => "1110100011100111",
42234 => "1110100011101000",
42235 => "1110100011101001",
42236 => "1110100011101011",
42237 => "1110100011101100",
42238 => "1110100011101101",
42239 => "1110100011101111",
42240 => "1110100011110000",
42241 => "1110100011110001",
42242 => "1110100011110011",
42243 => "1110100011110100",
42244 => "1110100011110101",
42245 => "1110100011110111",
42246 => "1110100011111000",
42247 => "1110100011111001",
42248 => "1110100011111010",
42249 => "1110100011111100",
42250 => "1110100011111101",
42251 => "1110100011111110",
42252 => "1110100100000000",
42253 => "1110100100000001",
42254 => "1110100100000010",
42255 => "1110100100000100",
42256 => "1110100100000101",
42257 => "1110100100000110",
42258 => "1110100100001000",
42259 => "1110100100001001",
42260 => "1110100100001010",
42261 => "1110100100001011",
42262 => "1110100100001101",
42263 => "1110100100001110",
42264 => "1110100100001111",
42265 => "1110100100010001",
42266 => "1110100100010010",
42267 => "1110100100010011",
42268 => "1110100100010101",
42269 => "1110100100010110",
42270 => "1110100100010111",
42271 => "1110100100011001",
42272 => "1110100100011010",
42273 => "1110100100011011",
42274 => "1110100100011100",
42275 => "1110100100011110",
42276 => "1110100100011111",
42277 => "1110100100100000",
42278 => "1110100100100010",
42279 => "1110100100100011",
42280 => "1110100100100100",
42281 => "1110100100100110",
42282 => "1110100100100111",
42283 => "1110100100101000",
42284 => "1110100100101001",
42285 => "1110100100101011",
42286 => "1110100100101100",
42287 => "1110100100101101",
42288 => "1110100100101111",
42289 => "1110100100110000",
42290 => "1110100100110001",
42291 => "1110100100110011",
42292 => "1110100100110100",
42293 => "1110100100110101",
42294 => "1110100100110110",
42295 => "1110100100111000",
42296 => "1110100100111001",
42297 => "1110100100111010",
42298 => "1110100100111100",
42299 => "1110100100111101",
42300 => "1110100100111110",
42301 => "1110100101000000",
42302 => "1110100101000001",
42303 => "1110100101000010",
42304 => "1110100101000011",
42305 => "1110100101000101",
42306 => "1110100101000110",
42307 => "1110100101000111",
42308 => "1110100101001001",
42309 => "1110100101001010",
42310 => "1110100101001011",
42311 => "1110100101001100",
42312 => "1110100101001110",
42313 => "1110100101001111",
42314 => "1110100101010000",
42315 => "1110100101010010",
42316 => "1110100101010011",
42317 => "1110100101010100",
42318 => "1110100101010110",
42319 => "1110100101010111",
42320 => "1110100101011000",
42321 => "1110100101011001",
42322 => "1110100101011011",
42323 => "1110100101011100",
42324 => "1110100101011101",
42325 => "1110100101011111",
42326 => "1110100101100000",
42327 => "1110100101100001",
42328 => "1110100101100010",
42329 => "1110100101100100",
42330 => "1110100101100101",
42331 => "1110100101100110",
42332 => "1110100101101000",
42333 => "1110100101101001",
42334 => "1110100101101010",
42335 => "1110100101101011",
42336 => "1110100101101101",
42337 => "1110100101101110",
42338 => "1110100101101111",
42339 => "1110100101110001",
42340 => "1110100101110010",
42341 => "1110100101110011",
42342 => "1110100101110100",
42343 => "1110100101110110",
42344 => "1110100101110111",
42345 => "1110100101111000",
42346 => "1110100101111010",
42347 => "1110100101111011",
42348 => "1110100101111100",
42349 => "1110100101111101",
42350 => "1110100101111111",
42351 => "1110100110000000",
42352 => "1110100110000001",
42353 => "1110100110000011",
42354 => "1110100110000100",
42355 => "1110100110000101",
42356 => "1110100110000110",
42357 => "1110100110001000",
42358 => "1110100110001001",
42359 => "1110100110001010",
42360 => "1110100110001100",
42361 => "1110100110001101",
42362 => "1110100110001110",
42363 => "1110100110001111",
42364 => "1110100110010001",
42365 => "1110100110010010",
42366 => "1110100110010011",
42367 => "1110100110010100",
42368 => "1110100110010110",
42369 => "1110100110010111",
42370 => "1110100110011000",
42371 => "1110100110011010",
42372 => "1110100110011011",
42373 => "1110100110011100",
42374 => "1110100110011101",
42375 => "1110100110011111",
42376 => "1110100110100000",
42377 => "1110100110100001",
42378 => "1110100110100011",
42379 => "1110100110100100",
42380 => "1110100110100101",
42381 => "1110100110100110",
42382 => "1110100110101000",
42383 => "1110100110101001",
42384 => "1110100110101010",
42385 => "1110100110101011",
42386 => "1110100110101101",
42387 => "1110100110101110",
42388 => "1110100110101111",
42389 => "1110100110110001",
42390 => "1110100110110010",
42391 => "1110100110110011",
42392 => "1110100110110100",
42393 => "1110100110110110",
42394 => "1110100110110111",
42395 => "1110100110111000",
42396 => "1110100110111001",
42397 => "1110100110111011",
42398 => "1110100110111100",
42399 => "1110100110111101",
42400 => "1110100110111111",
42401 => "1110100111000000",
42402 => "1110100111000001",
42403 => "1110100111000010",
42404 => "1110100111000100",
42405 => "1110100111000101",
42406 => "1110100111000110",
42407 => "1110100111000111",
42408 => "1110100111001001",
42409 => "1110100111001010",
42410 => "1110100111001011",
42411 => "1110100111001100",
42412 => "1110100111001110",
42413 => "1110100111001111",
42414 => "1110100111010000",
42415 => "1110100111010010",
42416 => "1110100111010011",
42417 => "1110100111010100",
42418 => "1110100111010101",
42419 => "1110100111010111",
42420 => "1110100111011000",
42421 => "1110100111011001",
42422 => "1110100111011010",
42423 => "1110100111011100",
42424 => "1110100111011101",
42425 => "1110100111011110",
42426 => "1110100111011111",
42427 => "1110100111100001",
42428 => "1110100111100010",
42429 => "1110100111100011",
42430 => "1110100111100100",
42431 => "1110100111100110",
42432 => "1110100111100111",
42433 => "1110100111101000",
42434 => "1110100111101010",
42435 => "1110100111101011",
42436 => "1110100111101100",
42437 => "1110100111101101",
42438 => "1110100111101111",
42439 => "1110100111110000",
42440 => "1110100111110001",
42441 => "1110100111110010",
42442 => "1110100111110100",
42443 => "1110100111110101",
42444 => "1110100111110110",
42445 => "1110100111110111",
42446 => "1110100111111001",
42447 => "1110100111111010",
42448 => "1110100111111011",
42449 => "1110100111111100",
42450 => "1110100111111110",
42451 => "1110100111111111",
42452 => "1110101000000000",
42453 => "1110101000000001",
42454 => "1110101000000011",
42455 => "1110101000000100",
42456 => "1110101000000101",
42457 => "1110101000000110",
42458 => "1110101000001000",
42459 => "1110101000001001",
42460 => "1110101000001010",
42461 => "1110101000001100",
42462 => "1110101000001101",
42463 => "1110101000001110",
42464 => "1110101000001111",
42465 => "1110101000010001",
42466 => "1110101000010010",
42467 => "1110101000010011",
42468 => "1110101000010100",
42469 => "1110101000010110",
42470 => "1110101000010111",
42471 => "1110101000011000",
42472 => "1110101000011001",
42473 => "1110101000011011",
42474 => "1110101000011100",
42475 => "1110101000011101",
42476 => "1110101000011110",
42477 => "1110101000100000",
42478 => "1110101000100001",
42479 => "1110101000100010",
42480 => "1110101000100011",
42481 => "1110101000100101",
42482 => "1110101000100110",
42483 => "1110101000100111",
42484 => "1110101000101000",
42485 => "1110101000101010",
42486 => "1110101000101011",
42487 => "1110101000101100",
42488 => "1110101000101101",
42489 => "1110101000101111",
42490 => "1110101000110000",
42491 => "1110101000110001",
42492 => "1110101000110010",
42493 => "1110101000110100",
42494 => "1110101000110101",
42495 => "1110101000110110",
42496 => "1110101000110111",
42497 => "1110101000111001",
42498 => "1110101000111010",
42499 => "1110101000111011",
42500 => "1110101000111100",
42501 => "1110101000111101",
42502 => "1110101000111111",
42503 => "1110101001000000",
42504 => "1110101001000001",
42505 => "1110101001000010",
42506 => "1110101001000100",
42507 => "1110101001000101",
42508 => "1110101001000110",
42509 => "1110101001000111",
42510 => "1110101001001001",
42511 => "1110101001001010",
42512 => "1110101001001011",
42513 => "1110101001001100",
42514 => "1110101001001110",
42515 => "1110101001001111",
42516 => "1110101001010000",
42517 => "1110101001010001",
42518 => "1110101001010011",
42519 => "1110101001010100",
42520 => "1110101001010101",
42521 => "1110101001010110",
42522 => "1110101001011000",
42523 => "1110101001011001",
42524 => "1110101001011010",
42525 => "1110101001011011",
42526 => "1110101001011101",
42527 => "1110101001011110",
42528 => "1110101001011111",
42529 => "1110101001100000",
42530 => "1110101001100001",
42531 => "1110101001100011",
42532 => "1110101001100100",
42533 => "1110101001100101",
42534 => "1110101001100110",
42535 => "1110101001101000",
42536 => "1110101001101001",
42537 => "1110101001101010",
42538 => "1110101001101011",
42539 => "1110101001101101",
42540 => "1110101001101110",
42541 => "1110101001101111",
42542 => "1110101001110000",
42543 => "1110101001110010",
42544 => "1110101001110011",
42545 => "1110101001110100",
42546 => "1110101001110101",
42547 => "1110101001110110",
42548 => "1110101001111000",
42549 => "1110101001111001",
42550 => "1110101001111010",
42551 => "1110101001111011",
42552 => "1110101001111101",
42553 => "1110101001111110",
42554 => "1110101001111111",
42555 => "1110101010000000",
42556 => "1110101010000010",
42557 => "1110101010000011",
42558 => "1110101010000100",
42559 => "1110101010000101",
42560 => "1110101010000110",
42561 => "1110101010001000",
42562 => "1110101010001001",
42563 => "1110101010001010",
42564 => "1110101010001011",
42565 => "1110101010001101",
42566 => "1110101010001110",
42567 => "1110101010001111",
42568 => "1110101010010000",
42569 => "1110101010010010",
42570 => "1110101010010011",
42571 => "1110101010010100",
42572 => "1110101010010101",
42573 => "1110101010010110",
42574 => "1110101010011000",
42575 => "1110101010011001",
42576 => "1110101010011010",
42577 => "1110101010011011",
42578 => "1110101010011101",
42579 => "1110101010011110",
42580 => "1110101010011111",
42581 => "1110101010100000",
42582 => "1110101010100001",
42583 => "1110101010100011",
42584 => "1110101010100100",
42585 => "1110101010100101",
42586 => "1110101010100110",
42587 => "1110101010101000",
42588 => "1110101010101001",
42589 => "1110101010101010",
42590 => "1110101010101011",
42591 => "1110101010101100",
42592 => "1110101010101110",
42593 => "1110101010101111",
42594 => "1110101010110000",
42595 => "1110101010110001",
42596 => "1110101010110011",
42597 => "1110101010110100",
42598 => "1110101010110101",
42599 => "1110101010110110",
42600 => "1110101010110111",
42601 => "1110101010111001",
42602 => "1110101010111010",
42603 => "1110101010111011",
42604 => "1110101010111100",
42605 => "1110101010111110",
42606 => "1110101010111111",
42607 => "1110101011000000",
42608 => "1110101011000001",
42609 => "1110101011000010",
42610 => "1110101011000100",
42611 => "1110101011000101",
42612 => "1110101011000110",
42613 => "1110101011000111",
42614 => "1110101011001000",
42615 => "1110101011001010",
42616 => "1110101011001011",
42617 => "1110101011001100",
42618 => "1110101011001101",
42619 => "1110101011001111",
42620 => "1110101011010000",
42621 => "1110101011010001",
42622 => "1110101011010010",
42623 => "1110101011010011",
42624 => "1110101011010101",
42625 => "1110101011010110",
42626 => "1110101011010111",
42627 => "1110101011011000",
42628 => "1110101011011001",
42629 => "1110101011011011",
42630 => "1110101011011100",
42631 => "1110101011011101",
42632 => "1110101011011110",
42633 => "1110101011100000",
42634 => "1110101011100001",
42635 => "1110101011100010",
42636 => "1110101011100011",
42637 => "1110101011100100",
42638 => "1110101011100110",
42639 => "1110101011100111",
42640 => "1110101011101000",
42641 => "1110101011101001",
42642 => "1110101011101010",
42643 => "1110101011101100",
42644 => "1110101011101101",
42645 => "1110101011101110",
42646 => "1110101011101111",
42647 => "1110101011110000",
42648 => "1110101011110010",
42649 => "1110101011110011",
42650 => "1110101011110100",
42651 => "1110101011110101",
42652 => "1110101011110111",
42653 => "1110101011111000",
42654 => "1110101011111001",
42655 => "1110101011111010",
42656 => "1110101011111011",
42657 => "1110101011111101",
42658 => "1110101011111110",
42659 => "1110101011111111",
42660 => "1110101100000000",
42661 => "1110101100000001",
42662 => "1110101100000011",
42663 => "1110101100000100",
42664 => "1110101100000101",
42665 => "1110101100000110",
42666 => "1110101100000111",
42667 => "1110101100001001",
42668 => "1110101100001010",
42669 => "1110101100001011",
42670 => "1110101100001100",
42671 => "1110101100001101",
42672 => "1110101100001111",
42673 => "1110101100010000",
42674 => "1110101100010001",
42675 => "1110101100010010",
42676 => "1110101100010011",
42677 => "1110101100010101",
42678 => "1110101100010110",
42679 => "1110101100010111",
42680 => "1110101100011000",
42681 => "1110101100011001",
42682 => "1110101100011011",
42683 => "1110101100011100",
42684 => "1110101100011101",
42685 => "1110101100011110",
42686 => "1110101100011111",
42687 => "1110101100100001",
42688 => "1110101100100010",
42689 => "1110101100100011",
42690 => "1110101100100100",
42691 => "1110101100100101",
42692 => "1110101100100111",
42693 => "1110101100101000",
42694 => "1110101100101001",
42695 => "1110101100101010",
42696 => "1110101100101011",
42697 => "1110101100101101",
42698 => "1110101100101110",
42699 => "1110101100101111",
42700 => "1110101100110000",
42701 => "1110101100110001",
42702 => "1110101100110011",
42703 => "1110101100110100",
42704 => "1110101100110101",
42705 => "1110101100110110",
42706 => "1110101100110111",
42707 => "1110101100111001",
42708 => "1110101100111010",
42709 => "1110101100111011",
42710 => "1110101100111100",
42711 => "1110101100111101",
42712 => "1110101100111110",
42713 => "1110101101000000",
42714 => "1110101101000001",
42715 => "1110101101000010",
42716 => "1110101101000011",
42717 => "1110101101000100",
42718 => "1110101101000110",
42719 => "1110101101000111",
42720 => "1110101101001000",
42721 => "1110101101001001",
42722 => "1110101101001010",
42723 => "1110101101001100",
42724 => "1110101101001101",
42725 => "1110101101001110",
42726 => "1110101101001111",
42727 => "1110101101010000",
42728 => "1110101101010010",
42729 => "1110101101010011",
42730 => "1110101101010100",
42731 => "1110101101010101",
42732 => "1110101101010110",
42733 => "1110101101010111",
42734 => "1110101101011001",
42735 => "1110101101011010",
42736 => "1110101101011011",
42737 => "1110101101011100",
42738 => "1110101101011101",
42739 => "1110101101011111",
42740 => "1110101101100000",
42741 => "1110101101100001",
42742 => "1110101101100010",
42743 => "1110101101100011",
42744 => "1110101101100100",
42745 => "1110101101100110",
42746 => "1110101101100111",
42747 => "1110101101101000",
42748 => "1110101101101001",
42749 => "1110101101101010",
42750 => "1110101101101100",
42751 => "1110101101101101",
42752 => "1110101101101110",
42753 => "1110101101101111",
42754 => "1110101101110000",
42755 => "1110101101110010",
42756 => "1110101101110011",
42757 => "1110101101110100",
42758 => "1110101101110101",
42759 => "1110101101110110",
42760 => "1110101101110111",
42761 => "1110101101111001",
42762 => "1110101101111010",
42763 => "1110101101111011",
42764 => "1110101101111100",
42765 => "1110101101111101",
42766 => "1110101101111110",
42767 => "1110101110000000",
42768 => "1110101110000001",
42769 => "1110101110000010",
42770 => "1110101110000011",
42771 => "1110101110000100",
42772 => "1110101110000110",
42773 => "1110101110000111",
42774 => "1110101110001000",
42775 => "1110101110001001",
42776 => "1110101110001010",
42777 => "1110101110001011",
42778 => "1110101110001101",
42779 => "1110101110001110",
42780 => "1110101110001111",
42781 => "1110101110010000",
42782 => "1110101110010001",
42783 => "1110101110010010",
42784 => "1110101110010100",
42785 => "1110101110010101",
42786 => "1110101110010110",
42787 => "1110101110010111",
42788 => "1110101110011000",
42789 => "1110101110011010",
42790 => "1110101110011011",
42791 => "1110101110011100",
42792 => "1110101110011101",
42793 => "1110101110011110",
42794 => "1110101110011111",
42795 => "1110101110100001",
42796 => "1110101110100010",
42797 => "1110101110100011",
42798 => "1110101110100100",
42799 => "1110101110100101",
42800 => "1110101110100110",
42801 => "1110101110101000",
42802 => "1110101110101001",
42803 => "1110101110101010",
42804 => "1110101110101011",
42805 => "1110101110101100",
42806 => "1110101110101101",
42807 => "1110101110101111",
42808 => "1110101110110000",
42809 => "1110101110110001",
42810 => "1110101110110010",
42811 => "1110101110110011",
42812 => "1110101110110100",
42813 => "1110101110110110",
42814 => "1110101110110111",
42815 => "1110101110111000",
42816 => "1110101110111001",
42817 => "1110101110111010",
42818 => "1110101110111011",
42819 => "1110101110111101",
42820 => "1110101110111110",
42821 => "1110101110111111",
42822 => "1110101111000000",
42823 => "1110101111000001",
42824 => "1110101111000010",
42825 => "1110101111000100",
42826 => "1110101111000101",
42827 => "1110101111000110",
42828 => "1110101111000111",
42829 => "1110101111001000",
42830 => "1110101111001001",
42831 => "1110101111001011",
42832 => "1110101111001100",
42833 => "1110101111001101",
42834 => "1110101111001110",
42835 => "1110101111001111",
42836 => "1110101111010000",
42837 => "1110101111010010",
42838 => "1110101111010011",
42839 => "1110101111010100",
42840 => "1110101111010101",
42841 => "1110101111010110",
42842 => "1110101111010111",
42843 => "1110101111011001",
42844 => "1110101111011010",
42845 => "1110101111011011",
42846 => "1110101111011100",
42847 => "1110101111011101",
42848 => "1110101111011110",
42849 => "1110101111100000",
42850 => "1110101111100001",
42851 => "1110101111100010",
42852 => "1110101111100011",
42853 => "1110101111100100",
42854 => "1110101111100101",
42855 => "1110101111100110",
42856 => "1110101111101000",
42857 => "1110101111101001",
42858 => "1110101111101010",
42859 => "1110101111101011",
42860 => "1110101111101100",
42861 => "1110101111101101",
42862 => "1110101111101111",
42863 => "1110101111110000",
42864 => "1110101111110001",
42865 => "1110101111110010",
42866 => "1110101111110011",
42867 => "1110101111110100",
42868 => "1110101111110101",
42869 => "1110101111110111",
42870 => "1110101111111000",
42871 => "1110101111111001",
42872 => "1110101111111010",
42873 => "1110101111111011",
42874 => "1110101111111100",
42875 => "1110101111111110",
42876 => "1110101111111111",
42877 => "1110110000000000",
42878 => "1110110000000001",
42879 => "1110110000000010",
42880 => "1110110000000011",
42881 => "1110110000000100",
42882 => "1110110000000110",
42883 => "1110110000000111",
42884 => "1110110000001000",
42885 => "1110110000001001",
42886 => "1110110000001010",
42887 => "1110110000001011",
42888 => "1110110000001101",
42889 => "1110110000001110",
42890 => "1110110000001111",
42891 => "1110110000010000",
42892 => "1110110000010001",
42893 => "1110110000010010",
42894 => "1110110000010011",
42895 => "1110110000010101",
42896 => "1110110000010110",
42897 => "1110110000010111",
42898 => "1110110000011000",
42899 => "1110110000011001",
42900 => "1110110000011010",
42901 => "1110110000011011",
42902 => "1110110000011101",
42903 => "1110110000011110",
42904 => "1110110000011111",
42905 => "1110110000100000",
42906 => "1110110000100001",
42907 => "1110110000100010",
42908 => "1110110000100011",
42909 => "1110110000100101",
42910 => "1110110000100110",
42911 => "1110110000100111",
42912 => "1110110000101000",
42913 => "1110110000101001",
42914 => "1110110000101010",
42915 => "1110110000101011",
42916 => "1110110000101101",
42917 => "1110110000101110",
42918 => "1110110000101111",
42919 => "1110110000110000",
42920 => "1110110000110001",
42921 => "1110110000110010",
42922 => "1110110000110011",
42923 => "1110110000110101",
42924 => "1110110000110110",
42925 => "1110110000110111",
42926 => "1110110000111000",
42927 => "1110110000111001",
42928 => "1110110000111010",
42929 => "1110110000111011",
42930 => "1110110000111101",
42931 => "1110110000111110",
42932 => "1110110000111111",
42933 => "1110110001000000",
42934 => "1110110001000001",
42935 => "1110110001000010",
42936 => "1110110001000011",
42937 => "1110110001000101",
42938 => "1110110001000110",
42939 => "1110110001000111",
42940 => "1110110001001000",
42941 => "1110110001001001",
42942 => "1110110001001010",
42943 => "1110110001001011",
42944 => "1110110001001101",
42945 => "1110110001001110",
42946 => "1110110001001111",
42947 => "1110110001010000",
42948 => "1110110001010001",
42949 => "1110110001010010",
42950 => "1110110001010011",
42951 => "1110110001010100",
42952 => "1110110001010110",
42953 => "1110110001010111",
42954 => "1110110001011000",
42955 => "1110110001011001",
42956 => "1110110001011010",
42957 => "1110110001011011",
42958 => "1110110001011100",
42959 => "1110110001011110",
42960 => "1110110001011111",
42961 => "1110110001100000",
42962 => "1110110001100001",
42963 => "1110110001100010",
42964 => "1110110001100011",
42965 => "1110110001100100",
42966 => "1110110001100101",
42967 => "1110110001100111",
42968 => "1110110001101000",
42969 => "1110110001101001",
42970 => "1110110001101010",
42971 => "1110110001101011",
42972 => "1110110001101100",
42973 => "1110110001101101",
42974 => "1110110001101111",
42975 => "1110110001110000",
42976 => "1110110001110001",
42977 => "1110110001110010",
42978 => "1110110001110011",
42979 => "1110110001110100",
42980 => "1110110001110101",
42981 => "1110110001110110",
42982 => "1110110001111000",
42983 => "1110110001111001",
42984 => "1110110001111010",
42985 => "1110110001111011",
42986 => "1110110001111100",
42987 => "1110110001111101",
42988 => "1110110001111110",
42989 => "1110110001111111",
42990 => "1110110010000001",
42991 => "1110110010000010",
42992 => "1110110010000011",
42993 => "1110110010000100",
42994 => "1110110010000101",
42995 => "1110110010000110",
42996 => "1110110010000111",
42997 => "1110110010001000",
42998 => "1110110010001010",
42999 => "1110110010001011",
43000 => "1110110010001100",
43001 => "1110110010001101",
43002 => "1110110010001110",
43003 => "1110110010001111",
43004 => "1110110010010000",
43005 => "1110110010010001",
43006 => "1110110010010011",
43007 => "1110110010010100",
43008 => "1110110010010101",
43009 => "1110110010010110",
43010 => "1110110010010111",
43011 => "1110110010011000",
43012 => "1110110010011001",
43013 => "1110110010011010",
43014 => "1110110010011100",
43015 => "1110110010011101",
43016 => "1110110010011110",
43017 => "1110110010011111",
43018 => "1110110010100000",
43019 => "1110110010100001",
43020 => "1110110010100010",
43021 => "1110110010100011",
43022 => "1110110010100100",
43023 => "1110110010100110",
43024 => "1110110010100111",
43025 => "1110110010101000",
43026 => "1110110010101001",
43027 => "1110110010101010",
43028 => "1110110010101011",
43029 => "1110110010101100",
43030 => "1110110010101101",
43031 => "1110110010101111",
43032 => "1110110010110000",
43033 => "1110110010110001",
43034 => "1110110010110010",
43035 => "1110110010110011",
43036 => "1110110010110100",
43037 => "1110110010110101",
43038 => "1110110010110110",
43039 => "1110110010110111",
43040 => "1110110010111001",
43041 => "1110110010111010",
43042 => "1110110010111011",
43043 => "1110110010111100",
43044 => "1110110010111101",
43045 => "1110110010111110",
43046 => "1110110010111111",
43047 => "1110110011000000",
43048 => "1110110011000001",
43049 => "1110110011000011",
43050 => "1110110011000100",
43051 => "1110110011000101",
43052 => "1110110011000110",
43053 => "1110110011000111",
43054 => "1110110011001000",
43055 => "1110110011001001",
43056 => "1110110011001010",
43057 => "1110110011001011",
43058 => "1110110011001101",
43059 => "1110110011001110",
43060 => "1110110011001111",
43061 => "1110110011010000",
43062 => "1110110011010001",
43063 => "1110110011010010",
43064 => "1110110011010011",
43065 => "1110110011010100",
43066 => "1110110011010101",
43067 => "1110110011010111",
43068 => "1110110011011000",
43069 => "1110110011011001",
43070 => "1110110011011010",
43071 => "1110110011011011",
43072 => "1110110011011100",
43073 => "1110110011011101",
43074 => "1110110011011110",
43075 => "1110110011011111",
43076 => "1110110011100001",
43077 => "1110110011100010",
43078 => "1110110011100011",
43079 => "1110110011100100",
43080 => "1110110011100101",
43081 => "1110110011100110",
43082 => "1110110011100111",
43083 => "1110110011101000",
43084 => "1110110011101001",
43085 => "1110110011101010",
43086 => "1110110011101100",
43087 => "1110110011101101",
43088 => "1110110011101110",
43089 => "1110110011101111",
43090 => "1110110011110000",
43091 => "1110110011110001",
43092 => "1110110011110010",
43093 => "1110110011110011",
43094 => "1110110011110100",
43095 => "1110110011110101",
43096 => "1110110011110111",
43097 => "1110110011111000",
43098 => "1110110011111001",
43099 => "1110110011111010",
43100 => "1110110011111011",
43101 => "1110110011111100",
43102 => "1110110011111101",
43103 => "1110110011111110",
43104 => "1110110011111111",
43105 => "1110110100000000",
43106 => "1110110100000010",
43107 => "1110110100000011",
43108 => "1110110100000100",
43109 => "1110110100000101",
43110 => "1110110100000110",
43111 => "1110110100000111",
43112 => "1110110100001000",
43113 => "1110110100001001",
43114 => "1110110100001010",
43115 => "1110110100001011",
43116 => "1110110100001101",
43117 => "1110110100001110",
43118 => "1110110100001111",
43119 => "1110110100010000",
43120 => "1110110100010001",
43121 => "1110110100010010",
43122 => "1110110100010011",
43123 => "1110110100010100",
43124 => "1110110100010101",
43125 => "1110110100010110",
43126 => "1110110100011000",
43127 => "1110110100011001",
43128 => "1110110100011010",
43129 => "1110110100011011",
43130 => "1110110100011100",
43131 => "1110110100011101",
43132 => "1110110100011110",
43133 => "1110110100011111",
43134 => "1110110100100000",
43135 => "1110110100100001",
43136 => "1110110100100010",
43137 => "1110110100100100",
43138 => "1110110100100101",
43139 => "1110110100100110",
43140 => "1110110100100111",
43141 => "1110110100101000",
43142 => "1110110100101001",
43143 => "1110110100101010",
43144 => "1110110100101011",
43145 => "1110110100101100",
43146 => "1110110100101101",
43147 => "1110110100101110",
43148 => "1110110100110000",
43149 => "1110110100110001",
43150 => "1110110100110010",
43151 => "1110110100110011",
43152 => "1110110100110100",
43153 => "1110110100110101",
43154 => "1110110100110110",
43155 => "1110110100110111",
43156 => "1110110100111000",
43157 => "1110110100111001",
43158 => "1110110100111010",
43159 => "1110110100111100",
43160 => "1110110100111101",
43161 => "1110110100111110",
43162 => "1110110100111111",
43163 => "1110110101000000",
43164 => "1110110101000001",
43165 => "1110110101000010",
43166 => "1110110101000011",
43167 => "1110110101000100",
43168 => "1110110101000101",
43169 => "1110110101000110",
43170 => "1110110101000111",
43171 => "1110110101001001",
43172 => "1110110101001010",
43173 => "1110110101001011",
43174 => "1110110101001100",
43175 => "1110110101001101",
43176 => "1110110101001110",
43177 => "1110110101001111",
43178 => "1110110101010000",
43179 => "1110110101010001",
43180 => "1110110101010010",
43181 => "1110110101010011",
43182 => "1110110101010100",
43183 => "1110110101010110",
43184 => "1110110101010111",
43185 => "1110110101011000",
43186 => "1110110101011001",
43187 => "1110110101011010",
43188 => "1110110101011011",
43189 => "1110110101011100",
43190 => "1110110101011101",
43191 => "1110110101011110",
43192 => "1110110101011111",
43193 => "1110110101100000",
43194 => "1110110101100001",
43195 => "1110110101100011",
43196 => "1110110101100100",
43197 => "1110110101100101",
43198 => "1110110101100110",
43199 => "1110110101100111",
43200 => "1110110101101000",
43201 => "1110110101101001",
43202 => "1110110101101010",
43203 => "1110110101101011",
43204 => "1110110101101100",
43205 => "1110110101101101",
43206 => "1110110101101110",
43207 => "1110110101101111",
43208 => "1110110101110001",
43209 => "1110110101110010",
43210 => "1110110101110011",
43211 => "1110110101110100",
43212 => "1110110101110101",
43213 => "1110110101110110",
43214 => "1110110101110111",
43215 => "1110110101111000",
43216 => "1110110101111001",
43217 => "1110110101111010",
43218 => "1110110101111011",
43219 => "1110110101111100",
43220 => "1110110101111101",
43221 => "1110110101111110",
43222 => "1110110110000000",
43223 => "1110110110000001",
43224 => "1110110110000010",
43225 => "1110110110000011",
43226 => "1110110110000100",
43227 => "1110110110000101",
43228 => "1110110110000110",
43229 => "1110110110000111",
43230 => "1110110110001000",
43231 => "1110110110001001",
43232 => "1110110110001010",
43233 => "1110110110001011",
43234 => "1110110110001100",
43235 => "1110110110001101",
43236 => "1110110110001111",
43237 => "1110110110010000",
43238 => "1110110110010001",
43239 => "1110110110010010",
43240 => "1110110110010011",
43241 => "1110110110010100",
43242 => "1110110110010101",
43243 => "1110110110010110",
43244 => "1110110110010111",
43245 => "1110110110011000",
43246 => "1110110110011001",
43247 => "1110110110011010",
43248 => "1110110110011011",
43249 => "1110110110011100",
43250 => "1110110110011101",
43251 => "1110110110011111",
43252 => "1110110110100000",
43253 => "1110110110100001",
43254 => "1110110110100010",
43255 => "1110110110100011",
43256 => "1110110110100100",
43257 => "1110110110100101",
43258 => "1110110110100110",
43259 => "1110110110100111",
43260 => "1110110110101000",
43261 => "1110110110101001",
43262 => "1110110110101010",
43263 => "1110110110101011",
43264 => "1110110110101100",
43265 => "1110110110101101",
43266 => "1110110110101111",
43267 => "1110110110110000",
43268 => "1110110110110001",
43269 => "1110110110110010",
43270 => "1110110110110011",
43271 => "1110110110110100",
43272 => "1110110110110101",
43273 => "1110110110110110",
43274 => "1110110110110111",
43275 => "1110110110111000",
43276 => "1110110110111001",
43277 => "1110110110111010",
43278 => "1110110110111011",
43279 => "1110110110111100",
43280 => "1110110110111101",
43281 => "1110110110111110",
43282 => "1110110111000000",
43283 => "1110110111000001",
43284 => "1110110111000010",
43285 => "1110110111000011",
43286 => "1110110111000100",
43287 => "1110110111000101",
43288 => "1110110111000110",
43289 => "1110110111000111",
43290 => "1110110111001000",
43291 => "1110110111001001",
43292 => "1110110111001010",
43293 => "1110110111001011",
43294 => "1110110111001100",
43295 => "1110110111001101",
43296 => "1110110111001110",
43297 => "1110110111001111",
43298 => "1110110111010000",
43299 => "1110110111010001",
43300 => "1110110111010011",
43301 => "1110110111010100",
43302 => "1110110111010101",
43303 => "1110110111010110",
43304 => "1110110111010111",
43305 => "1110110111011000",
43306 => "1110110111011001",
43307 => "1110110111011010",
43308 => "1110110111011011",
43309 => "1110110111011100",
43310 => "1110110111011101",
43311 => "1110110111011110",
43312 => "1110110111011111",
43313 => "1110110111100000",
43314 => "1110110111100001",
43315 => "1110110111100010",
43316 => "1110110111100011",
43317 => "1110110111100100",
43318 => "1110110111100101",
43319 => "1110110111100111",
43320 => "1110110111101000",
43321 => "1110110111101001",
43322 => "1110110111101010",
43323 => "1110110111101011",
43324 => "1110110111101100",
43325 => "1110110111101101",
43326 => "1110110111101110",
43327 => "1110110111101111",
43328 => "1110110111110000",
43329 => "1110110111110001",
43330 => "1110110111110010",
43331 => "1110110111110011",
43332 => "1110110111110100",
43333 => "1110110111110101",
43334 => "1110110111110110",
43335 => "1110110111110111",
43336 => "1110110111111000",
43337 => "1110110111111001",
43338 => "1110110111111010",
43339 => "1110110111111100",
43340 => "1110110111111101",
43341 => "1110110111111110",
43342 => "1110110111111111",
43343 => "1110111000000000",
43344 => "1110111000000001",
43345 => "1110111000000010",
43346 => "1110111000000011",
43347 => "1110111000000100",
43348 => "1110111000000101",
43349 => "1110111000000110",
43350 => "1110111000000111",
43351 => "1110111000001000",
43352 => "1110111000001001",
43353 => "1110111000001010",
43354 => "1110111000001011",
43355 => "1110111000001100",
43356 => "1110111000001101",
43357 => "1110111000001110",
43358 => "1110111000001111",
43359 => "1110111000010000",
43360 => "1110111000010001",
43361 => "1110111000010011",
43362 => "1110111000010100",
43363 => "1110111000010101",
43364 => "1110111000010110",
43365 => "1110111000010111",
43366 => "1110111000011000",
43367 => "1110111000011001",
43368 => "1110111000011010",
43369 => "1110111000011011",
43370 => "1110111000011100",
43371 => "1110111000011101",
43372 => "1110111000011110",
43373 => "1110111000011111",
43374 => "1110111000100000",
43375 => "1110111000100001",
43376 => "1110111000100010",
43377 => "1110111000100011",
43378 => "1110111000100100",
43379 => "1110111000100101",
43380 => "1110111000100110",
43381 => "1110111000100111",
43382 => "1110111000101000",
43383 => "1110111000101001",
43384 => "1110111000101010",
43385 => "1110111000101011",
43386 => "1110111000101100",
43387 => "1110111000101110",
43388 => "1110111000101111",
43389 => "1110111000110000",
43390 => "1110111000110001",
43391 => "1110111000110010",
43392 => "1110111000110011",
43393 => "1110111000110100",
43394 => "1110111000110101",
43395 => "1110111000110110",
43396 => "1110111000110111",
43397 => "1110111000111000",
43398 => "1110111000111001",
43399 => "1110111000111010",
43400 => "1110111000111011",
43401 => "1110111000111100",
43402 => "1110111000111101",
43403 => "1110111000111110",
43404 => "1110111000111111",
43405 => "1110111001000000",
43406 => "1110111001000001",
43407 => "1110111001000010",
43408 => "1110111001000011",
43409 => "1110111001000100",
43410 => "1110111001000101",
43411 => "1110111001000110",
43412 => "1110111001000111",
43413 => "1110111001001000",
43414 => "1110111001001001",
43415 => "1110111001001010",
43416 => "1110111001001011",
43417 => "1110111001001101",
43418 => "1110111001001110",
43419 => "1110111001001111",
43420 => "1110111001010000",
43421 => "1110111001010001",
43422 => "1110111001010010",
43423 => "1110111001010011",
43424 => "1110111001010100",
43425 => "1110111001010101",
43426 => "1110111001010110",
43427 => "1110111001010111",
43428 => "1110111001011000",
43429 => "1110111001011001",
43430 => "1110111001011010",
43431 => "1110111001011011",
43432 => "1110111001011100",
43433 => "1110111001011101",
43434 => "1110111001011110",
43435 => "1110111001011111",
43436 => "1110111001100000",
43437 => "1110111001100001",
43438 => "1110111001100010",
43439 => "1110111001100011",
43440 => "1110111001100100",
43441 => "1110111001100101",
43442 => "1110111001100110",
43443 => "1110111001100111",
43444 => "1110111001101000",
43445 => "1110111001101001",
43446 => "1110111001101010",
43447 => "1110111001101011",
43448 => "1110111001101100",
43449 => "1110111001101101",
43450 => "1110111001101110",
43451 => "1110111001101111",
43452 => "1110111001110000",
43453 => "1110111001110001",
43454 => "1110111001110010",
43455 => "1110111001110011",
43456 => "1110111001110101",
43457 => "1110111001110110",
43458 => "1110111001110111",
43459 => "1110111001111000",
43460 => "1110111001111001",
43461 => "1110111001111010",
43462 => "1110111001111011",
43463 => "1110111001111100",
43464 => "1110111001111101",
43465 => "1110111001111110",
43466 => "1110111001111111",
43467 => "1110111010000000",
43468 => "1110111010000001",
43469 => "1110111010000010",
43470 => "1110111010000011",
43471 => "1110111010000100",
43472 => "1110111010000101",
43473 => "1110111010000110",
43474 => "1110111010000111",
43475 => "1110111010001000",
43476 => "1110111010001001",
43477 => "1110111010001010",
43478 => "1110111010001011",
43479 => "1110111010001100",
43480 => "1110111010001101",
43481 => "1110111010001110",
43482 => "1110111010001111",
43483 => "1110111010010000",
43484 => "1110111010010001",
43485 => "1110111010010010",
43486 => "1110111010010011",
43487 => "1110111010010100",
43488 => "1110111010010101",
43489 => "1110111010010110",
43490 => "1110111010010111",
43491 => "1110111010011000",
43492 => "1110111010011001",
43493 => "1110111010011010",
43494 => "1110111010011011",
43495 => "1110111010011100",
43496 => "1110111010011101",
43497 => "1110111010011110",
43498 => "1110111010011111",
43499 => "1110111010100000",
43500 => "1110111010100001",
43501 => "1110111010100010",
43502 => "1110111010100011",
43503 => "1110111010100100",
43504 => "1110111010100101",
43505 => "1110111010100110",
43506 => "1110111010100111",
43507 => "1110111010101000",
43508 => "1110111010101001",
43509 => "1110111010101010",
43510 => "1110111010101011",
43511 => "1110111010101100",
43512 => "1110111010101101",
43513 => "1110111010101110",
43514 => "1110111010101111",
43515 => "1110111010110000",
43516 => "1110111010110001",
43517 => "1110111010110010",
43518 => "1110111010110011",
43519 => "1110111010110100",
43520 => "1110111010110101",
43521 => "1110111010110110",
43522 => "1110111010110111",
43523 => "1110111010111000",
43524 => "1110111010111001",
43525 => "1110111010111010",
43526 => "1110111010111011",
43527 => "1110111010111100",
43528 => "1110111010111101",
43529 => "1110111010111110",
43530 => "1110111010111111",
43531 => "1110111011000001",
43532 => "1110111011000010",
43533 => "1110111011000011",
43534 => "1110111011000100",
43535 => "1110111011000101",
43536 => "1110111011000110",
43537 => "1110111011000111",
43538 => "1110111011001000",
43539 => "1110111011001001",
43540 => "1110111011001010",
43541 => "1110111011001011",
43542 => "1110111011001100",
43543 => "1110111011001101",
43544 => "1110111011001110",
43545 => "1110111011001111",
43546 => "1110111011010000",
43547 => "1110111011010001",
43548 => "1110111011010010",
43549 => "1110111011010011",
43550 => "1110111011010100",
43551 => "1110111011010101",
43552 => "1110111011010110",
43553 => "1110111011010111",
43554 => "1110111011011000",
43555 => "1110111011011001",
43556 => "1110111011011010",
43557 => "1110111011011011",
43558 => "1110111011011100",
43559 => "1110111011011101",
43560 => "1110111011011110",
43561 => "1110111011011111",
43562 => "1110111011100000",
43563 => "1110111011100001",
43564 => "1110111011100010",
43565 => "1110111011100011",
43566 => "1110111011100100",
43567 => "1110111011100101",
43568 => "1110111011100110",
43569 => "1110111011100111",
43570 => "1110111011101000",
43571 => "1110111011101001",
43572 => "1110111011101010",
43573 => "1110111011101011",
43574 => "1110111011101100",
43575 => "1110111011101101",
43576 => "1110111011101110",
43577 => "1110111011101111",
43578 => "1110111011110000",
43579 => "1110111011110001",
43580 => "1110111011110010",
43581 => "1110111011110010",
43582 => "1110111011110011",
43583 => "1110111011110100",
43584 => "1110111011110101",
43585 => "1110111011110110",
43586 => "1110111011110111",
43587 => "1110111011111000",
43588 => "1110111011111001",
43589 => "1110111011111010",
43590 => "1110111011111011",
43591 => "1110111011111100",
43592 => "1110111011111101",
43593 => "1110111011111110",
43594 => "1110111011111111",
43595 => "1110111100000000",
43596 => "1110111100000001",
43597 => "1110111100000010",
43598 => "1110111100000011",
43599 => "1110111100000100",
43600 => "1110111100000101",
43601 => "1110111100000110",
43602 => "1110111100000111",
43603 => "1110111100001000",
43604 => "1110111100001001",
43605 => "1110111100001010",
43606 => "1110111100001011",
43607 => "1110111100001100",
43608 => "1110111100001101",
43609 => "1110111100001110",
43610 => "1110111100001111",
43611 => "1110111100010000",
43612 => "1110111100010001",
43613 => "1110111100010010",
43614 => "1110111100010011",
43615 => "1110111100010100",
43616 => "1110111100010101",
43617 => "1110111100010110",
43618 => "1110111100010111",
43619 => "1110111100011000",
43620 => "1110111100011001",
43621 => "1110111100011010",
43622 => "1110111100011011",
43623 => "1110111100011100",
43624 => "1110111100011101",
43625 => "1110111100011110",
43626 => "1110111100011111",
43627 => "1110111100100000",
43628 => "1110111100100001",
43629 => "1110111100100010",
43630 => "1110111100100011",
43631 => "1110111100100100",
43632 => "1110111100100101",
43633 => "1110111100100110",
43634 => "1110111100100111",
43635 => "1110111100101000",
43636 => "1110111100101001",
43637 => "1110111100101010",
43638 => "1110111100101011",
43639 => "1110111100101100",
43640 => "1110111100101101",
43641 => "1110111100101110",
43642 => "1110111100101111",
43643 => "1110111100110000",
43644 => "1110111100110001",
43645 => "1110111100110010",
43646 => "1110111100110011",
43647 => "1110111100110100",
43648 => "1110111100110101",
43649 => "1110111100110110",
43650 => "1110111100110111",
43651 => "1110111100111000",
43652 => "1110111100111001",
43653 => "1110111100111010",
43654 => "1110111100111011",
43655 => "1110111100111100",
43656 => "1110111100111101",
43657 => "1110111100111101",
43658 => "1110111100111110",
43659 => "1110111100111111",
43660 => "1110111101000000",
43661 => "1110111101000001",
43662 => "1110111101000010",
43663 => "1110111101000011",
43664 => "1110111101000100",
43665 => "1110111101000101",
43666 => "1110111101000110",
43667 => "1110111101000111",
43668 => "1110111101001000",
43669 => "1110111101001001",
43670 => "1110111101001010",
43671 => "1110111101001011",
43672 => "1110111101001100",
43673 => "1110111101001101",
43674 => "1110111101001110",
43675 => "1110111101001111",
43676 => "1110111101010000",
43677 => "1110111101010001",
43678 => "1110111101010010",
43679 => "1110111101010011",
43680 => "1110111101010100",
43681 => "1110111101010101",
43682 => "1110111101010110",
43683 => "1110111101010111",
43684 => "1110111101011000",
43685 => "1110111101011001",
43686 => "1110111101011010",
43687 => "1110111101011011",
43688 => "1110111101011100",
43689 => "1110111101011101",
43690 => "1110111101011110",
43691 => "1110111101011111",
43692 => "1110111101100000",
43693 => "1110111101100001",
43694 => "1110111101100010",
43695 => "1110111101100011",
43696 => "1110111101100100",
43697 => "1110111101100100",
43698 => "1110111101100101",
43699 => "1110111101100110",
43700 => "1110111101100111",
43701 => "1110111101101000",
43702 => "1110111101101001",
43703 => "1110111101101010",
43704 => "1110111101101011",
43705 => "1110111101101100",
43706 => "1110111101101101",
43707 => "1110111101101110",
43708 => "1110111101101111",
43709 => "1110111101110000",
43710 => "1110111101110001",
43711 => "1110111101110010",
43712 => "1110111101110011",
43713 => "1110111101110100",
43714 => "1110111101110101",
43715 => "1110111101110110",
43716 => "1110111101110111",
43717 => "1110111101111000",
43718 => "1110111101111001",
43719 => "1110111101111010",
43720 => "1110111101111011",
43721 => "1110111101111100",
43722 => "1110111101111101",
43723 => "1110111101111110",
43724 => "1110111101111111",
43725 => "1110111110000000",
43726 => "1110111110000001",
43727 => "1110111110000010",
43728 => "1110111110000010",
43729 => "1110111110000011",
43730 => "1110111110000100",
43731 => "1110111110000101",
43732 => "1110111110000110",
43733 => "1110111110000111",
43734 => "1110111110001000",
43735 => "1110111110001001",
43736 => "1110111110001010",
43737 => "1110111110001011",
43738 => "1110111110001100",
43739 => "1110111110001101",
43740 => "1110111110001110",
43741 => "1110111110001111",
43742 => "1110111110010000",
43743 => "1110111110010001",
43744 => "1110111110010010",
43745 => "1110111110010011",
43746 => "1110111110010100",
43747 => "1110111110010101",
43748 => "1110111110010110",
43749 => "1110111110010111",
43750 => "1110111110011000",
43751 => "1110111110011001",
43752 => "1110111110011010",
43753 => "1110111110011011",
43754 => "1110111110011011",
43755 => "1110111110011100",
43756 => "1110111110011101",
43757 => "1110111110011110",
43758 => "1110111110011111",
43759 => "1110111110100000",
43760 => "1110111110100001",
43761 => "1110111110100010",
43762 => "1110111110100011",
43763 => "1110111110100100",
43764 => "1110111110100101",
43765 => "1110111110100110",
43766 => "1110111110100111",
43767 => "1110111110101000",
43768 => "1110111110101001",
43769 => "1110111110101010",
43770 => "1110111110101011",
43771 => "1110111110101100",
43772 => "1110111110101101",
43773 => "1110111110101110",
43774 => "1110111110101111",
43775 => "1110111110110000",
43776 => "1110111110110001",
43777 => "1110111110110001",
43778 => "1110111110110010",
43779 => "1110111110110011",
43780 => "1110111110110100",
43781 => "1110111110110101",
43782 => "1110111110110110",
43783 => "1110111110110111",
43784 => "1110111110111000",
43785 => "1110111110111001",
43786 => "1110111110111010",
43787 => "1110111110111011",
43788 => "1110111110111100",
43789 => "1110111110111101",
43790 => "1110111110111110",
43791 => "1110111110111111",
43792 => "1110111111000000",
43793 => "1110111111000001",
43794 => "1110111111000010",
43795 => "1110111111000011",
43796 => "1110111111000100",
43797 => "1110111111000101",
43798 => "1110111111000101",
43799 => "1110111111000110",
43800 => "1110111111000111",
43801 => "1110111111001000",
43802 => "1110111111001001",
43803 => "1110111111001010",
43804 => "1110111111001011",
43805 => "1110111111001100",
43806 => "1110111111001101",
43807 => "1110111111001110",
43808 => "1110111111001111",
43809 => "1110111111010000",
43810 => "1110111111010001",
43811 => "1110111111010010",
43812 => "1110111111010011",
43813 => "1110111111010100",
43814 => "1110111111010101",
43815 => "1110111111010110",
43816 => "1110111111010111",
43817 => "1110111111010111",
43818 => "1110111111011000",
43819 => "1110111111011001",
43820 => "1110111111011010",
43821 => "1110111111011011",
43822 => "1110111111011100",
43823 => "1110111111011101",
43824 => "1110111111011110",
43825 => "1110111111011111",
43826 => "1110111111100000",
43827 => "1110111111100001",
43828 => "1110111111100010",
43829 => "1110111111100011",
43830 => "1110111111100100",
43831 => "1110111111100101",
43832 => "1110111111100110",
43833 => "1110111111100111",
43834 => "1110111111101000",
43835 => "1110111111101000",
43836 => "1110111111101001",
43837 => "1110111111101010",
43838 => "1110111111101011",
43839 => "1110111111101100",
43840 => "1110111111101101",
43841 => "1110111111101110",
43842 => "1110111111101111",
43843 => "1110111111110000",
43844 => "1110111111110001",
43845 => "1110111111110010",
43846 => "1110111111110011",
43847 => "1110111111110100",
43848 => "1110111111110101",
43849 => "1110111111110110",
43850 => "1110111111110111",
43851 => "1110111111111000",
43852 => "1110111111111000",
43853 => "1110111111111001",
43854 => "1110111111111010",
43855 => "1110111111111011",
43856 => "1110111111111100",
43857 => "1110111111111101",
43858 => "1110111111111110",
43859 => "1110111111111111",
43860 => "1111000000000000",
43861 => "1111000000000001",
43862 => "1111000000000010",
43863 => "1111000000000011",
43864 => "1111000000000100",
43865 => "1111000000000101",
43866 => "1111000000000110",
43867 => "1111000000000111",
43868 => "1111000000000111",
43869 => "1111000000001000",
43870 => "1111000000001001",
43871 => "1111000000001010",
43872 => "1111000000001011",
43873 => "1111000000001100",
43874 => "1111000000001101",
43875 => "1111000000001110",
43876 => "1111000000001111",
43877 => "1111000000010000",
43878 => "1111000000010001",
43879 => "1111000000010010",
43880 => "1111000000010011",
43881 => "1111000000010100",
43882 => "1111000000010101",
43883 => "1111000000010101",
43884 => "1111000000010110",
43885 => "1111000000010111",
43886 => "1111000000011000",
43887 => "1111000000011001",
43888 => "1111000000011010",
43889 => "1111000000011011",
43890 => "1111000000011100",
43891 => "1111000000011101",
43892 => "1111000000011110",
43893 => "1111000000011111",
43894 => "1111000000100000",
43895 => "1111000000100001",
43896 => "1111000000100010",
43897 => "1111000000100011",
43898 => "1111000000100011",
43899 => "1111000000100100",
43900 => "1111000000100101",
43901 => "1111000000100110",
43902 => "1111000000100111",
43903 => "1111000000101000",
43904 => "1111000000101001",
43905 => "1111000000101010",
43906 => "1111000000101011",
43907 => "1111000000101100",
43908 => "1111000000101101",
43909 => "1111000000101110",
43910 => "1111000000101111",
43911 => "1111000000110000",
43912 => "1111000000110000",
43913 => "1111000000110001",
43914 => "1111000000110010",
43915 => "1111000000110011",
43916 => "1111000000110100",
43917 => "1111000000110101",
43918 => "1111000000110110",
43919 => "1111000000110111",
43920 => "1111000000111000",
43921 => "1111000000111001",
43922 => "1111000000111010",
43923 => "1111000000111011",
43924 => "1111000000111100",
43925 => "1111000000111100",
43926 => "1111000000111101",
43927 => "1111000000111110",
43928 => "1111000000111111",
43929 => "1111000001000000",
43930 => "1111000001000001",
43931 => "1111000001000010",
43932 => "1111000001000011",
43933 => "1111000001000100",
43934 => "1111000001000101",
43935 => "1111000001000110",
43936 => "1111000001000111",
43937 => "1111000001001000",
43938 => "1111000001001000",
43939 => "1111000001001001",
43940 => "1111000001001010",
43941 => "1111000001001011",
43942 => "1111000001001100",
43943 => "1111000001001101",
43944 => "1111000001001110",
43945 => "1111000001001111",
43946 => "1111000001010000",
43947 => "1111000001010001",
43948 => "1111000001010010",
43949 => "1111000001010011",
43950 => "1111000001010100",
43951 => "1111000001010100",
43952 => "1111000001010101",
43953 => "1111000001010110",
43954 => "1111000001010111",
43955 => "1111000001011000",
43956 => "1111000001011001",
43957 => "1111000001011010",
43958 => "1111000001011011",
43959 => "1111000001011100",
43960 => "1111000001011101",
43961 => "1111000001011110",
43962 => "1111000001011111",
43963 => "1111000001011111",
43964 => "1111000001100000",
43965 => "1111000001100001",
43966 => "1111000001100010",
43967 => "1111000001100011",
43968 => "1111000001100100",
43969 => "1111000001100101",
43970 => "1111000001100110",
43971 => "1111000001100111",
43972 => "1111000001101000",
43973 => "1111000001101001",
43974 => "1111000001101010",
43975 => "1111000001101010",
43976 => "1111000001101011",
43977 => "1111000001101100",
43978 => "1111000001101101",
43979 => "1111000001101110",
43980 => "1111000001101111",
43981 => "1111000001110000",
43982 => "1111000001110001",
43983 => "1111000001110010",
43984 => "1111000001110011",
43985 => "1111000001110100",
43986 => "1111000001110101",
43987 => "1111000001110101",
43988 => "1111000001110110",
43989 => "1111000001110111",
43990 => "1111000001111000",
43991 => "1111000001111001",
43992 => "1111000001111010",
43993 => "1111000001111011",
43994 => "1111000001111100",
43995 => "1111000001111101",
43996 => "1111000001111110",
43997 => "1111000001111111",
43998 => "1111000001111111",
43999 => "1111000010000000",
44000 => "1111000010000001",
44001 => "1111000010000010",
44002 => "1111000010000011",
44003 => "1111000010000100",
44004 => "1111000010000101",
44005 => "1111000010000110",
44006 => "1111000010000111",
44007 => "1111000010001000",
44008 => "1111000010001001",
44009 => "1111000010001001",
44010 => "1111000010001010",
44011 => "1111000010001011",
44012 => "1111000010001100",
44013 => "1111000010001101",
44014 => "1111000010001110",
44015 => "1111000010001111",
44016 => "1111000010010000",
44017 => "1111000010010001",
44018 => "1111000010010010",
44019 => "1111000010010011",
44020 => "1111000010010011",
44021 => "1111000010010100",
44022 => "1111000010010101",
44023 => "1111000010010110",
44024 => "1111000010010111",
44025 => "1111000010011000",
44026 => "1111000010011001",
44027 => "1111000010011010",
44028 => "1111000010011011",
44029 => "1111000010011100",
44030 => "1111000010011100",
44031 => "1111000010011101",
44032 => "1111000010011110",
44033 => "1111000010011111",
44034 => "1111000010100000",
44035 => "1111000010100001",
44036 => "1111000010100010",
44037 => "1111000010100011",
44038 => "1111000010100100",
44039 => "1111000010100101",
44040 => "1111000010100101",
44041 => "1111000010100110",
44042 => "1111000010100111",
44043 => "1111000010101000",
44044 => "1111000010101001",
44045 => "1111000010101010",
44046 => "1111000010101011",
44047 => "1111000010101100",
44048 => "1111000010101101",
44049 => "1111000010101110",
44050 => "1111000010101111",
44051 => "1111000010101111",
44052 => "1111000010110000",
44053 => "1111000010110001",
44054 => "1111000010110010",
44055 => "1111000010110011",
44056 => "1111000010110100",
44057 => "1111000010110101",
44058 => "1111000010110110",
44059 => "1111000010110111",
44060 => "1111000010110111",
44061 => "1111000010111000",
44062 => "1111000010111001",
44063 => "1111000010111010",
44064 => "1111000010111011",
44065 => "1111000010111100",
44066 => "1111000010111101",
44067 => "1111000010111110",
44068 => "1111000010111111",
44069 => "1111000011000000",
44070 => "1111000011000000",
44071 => "1111000011000001",
44072 => "1111000011000010",
44073 => "1111000011000011",
44074 => "1111000011000100",
44075 => "1111000011000101",
44076 => "1111000011000110",
44077 => "1111000011000111",
44078 => "1111000011001000",
44079 => "1111000011001001",
44080 => "1111000011001001",
44081 => "1111000011001010",
44082 => "1111000011001011",
44083 => "1111000011001100",
44084 => "1111000011001101",
44085 => "1111000011001110",
44086 => "1111000011001111",
44087 => "1111000011010000",
44088 => "1111000011010001",
44089 => "1111000011010001",
44090 => "1111000011010010",
44091 => "1111000011010011",
44092 => "1111000011010100",
44093 => "1111000011010101",
44094 => "1111000011010110",
44095 => "1111000011010111",
44096 => "1111000011011000",
44097 => "1111000011011001",
44098 => "1111000011011001",
44099 => "1111000011011010",
44100 => "1111000011011011",
44101 => "1111000011011100",
44102 => "1111000011011101",
44103 => "1111000011011110",
44104 => "1111000011011111",
44105 => "1111000011100000",
44106 => "1111000011100001",
44107 => "1111000011100001",
44108 => "1111000011100010",
44109 => "1111000011100011",
44110 => "1111000011100100",
44111 => "1111000011100101",
44112 => "1111000011100110",
44113 => "1111000011100111",
44114 => "1111000011101000",
44115 => "1111000011101001",
44116 => "1111000011101001",
44117 => "1111000011101010",
44118 => "1111000011101011",
44119 => "1111000011101100",
44120 => "1111000011101101",
44121 => "1111000011101110",
44122 => "1111000011101111",
44123 => "1111000011110000",
44124 => "1111000011110001",
44125 => "1111000011110001",
44126 => "1111000011110010",
44127 => "1111000011110011",
44128 => "1111000011110100",
44129 => "1111000011110101",
44130 => "1111000011110110",
44131 => "1111000011110111",
44132 => "1111000011111000",
44133 => "1111000011111001",
44134 => "1111000011111001",
44135 => "1111000011111010",
44136 => "1111000011111011",
44137 => "1111000011111100",
44138 => "1111000011111101",
44139 => "1111000011111110",
44140 => "1111000011111111",
44141 => "1111000100000000",
44142 => "1111000100000000",
44143 => "1111000100000001",
44144 => "1111000100000010",
44145 => "1111000100000011",
44146 => "1111000100000100",
44147 => "1111000100000101",
44148 => "1111000100000110",
44149 => "1111000100000111",
44150 => "1111000100001000",
44151 => "1111000100001000",
44152 => "1111000100001001",
44153 => "1111000100001010",
44154 => "1111000100001011",
44155 => "1111000100001100",
44156 => "1111000100001101",
44157 => "1111000100001110",
44158 => "1111000100001111",
44159 => "1111000100001111",
44160 => "1111000100010000",
44161 => "1111000100010001",
44162 => "1111000100010010",
44163 => "1111000100010011",
44164 => "1111000100010100",
44165 => "1111000100010101",
44166 => "1111000100010110",
44167 => "1111000100010110",
44168 => "1111000100010111",
44169 => "1111000100011000",
44170 => "1111000100011001",
44171 => "1111000100011010",
44172 => "1111000100011011",
44173 => "1111000100011100",
44174 => "1111000100011101",
44175 => "1111000100011110",
44176 => "1111000100011110",
44177 => "1111000100011111",
44178 => "1111000100100000",
44179 => "1111000100100001",
44180 => "1111000100100010",
44181 => "1111000100100011",
44182 => "1111000100100100",
44183 => "1111000100100101",
44184 => "1111000100100101",
44185 => "1111000100100110",
44186 => "1111000100100111",
44187 => "1111000100101000",
44188 => "1111000100101001",
44189 => "1111000100101010",
44190 => "1111000100101011",
44191 => "1111000100101011",
44192 => "1111000100101100",
44193 => "1111000100101101",
44194 => "1111000100101110",
44195 => "1111000100101111",
44196 => "1111000100110000",
44197 => "1111000100110001",
44198 => "1111000100110010",
44199 => "1111000100110010",
44200 => "1111000100110011",
44201 => "1111000100110100",
44202 => "1111000100110101",
44203 => "1111000100110110",
44204 => "1111000100110111",
44205 => "1111000100111000",
44206 => "1111000100111001",
44207 => "1111000100111001",
44208 => "1111000100111010",
44209 => "1111000100111011",
44210 => "1111000100111100",
44211 => "1111000100111101",
44212 => "1111000100111110",
44213 => "1111000100111111",
44214 => "1111000101000000",
44215 => "1111000101000000",
44216 => "1111000101000001",
44217 => "1111000101000010",
44218 => "1111000101000011",
44219 => "1111000101000100",
44220 => "1111000101000101",
44221 => "1111000101000110",
44222 => "1111000101000110",
44223 => "1111000101000111",
44224 => "1111000101001000",
44225 => "1111000101001001",
44226 => "1111000101001010",
44227 => "1111000101001011",
44228 => "1111000101001100",
44229 => "1111000101001101",
44230 => "1111000101001101",
44231 => "1111000101001110",
44232 => "1111000101001111",
44233 => "1111000101010000",
44234 => "1111000101010001",
44235 => "1111000101010010",
44236 => "1111000101010011",
44237 => "1111000101010011",
44238 => "1111000101010100",
44239 => "1111000101010101",
44240 => "1111000101010110",
44241 => "1111000101010111",
44242 => "1111000101011000",
44243 => "1111000101011001",
44244 => "1111000101011010",
44245 => "1111000101011010",
44246 => "1111000101011011",
44247 => "1111000101011100",
44248 => "1111000101011101",
44249 => "1111000101011110",
44250 => "1111000101011111",
44251 => "1111000101100000",
44252 => "1111000101100000",
44253 => "1111000101100001",
44254 => "1111000101100010",
44255 => "1111000101100011",
44256 => "1111000101100100",
44257 => "1111000101100101",
44258 => "1111000101100110",
44259 => "1111000101100110",
44260 => "1111000101100111",
44261 => "1111000101101000",
44262 => "1111000101101001",
44263 => "1111000101101010",
44264 => "1111000101101011",
44265 => "1111000101101100",
44266 => "1111000101101100",
44267 => "1111000101101101",
44268 => "1111000101101110",
44269 => "1111000101101111",
44270 => "1111000101110000",
44271 => "1111000101110001",
44272 => "1111000101110010",
44273 => "1111000101110010",
44274 => "1111000101110011",
44275 => "1111000101110100",
44276 => "1111000101110101",
44277 => "1111000101110110",
44278 => "1111000101110111",
44279 => "1111000101111000",
44280 => "1111000101111000",
44281 => "1111000101111001",
44282 => "1111000101111010",
44283 => "1111000101111011",
44284 => "1111000101111100",
44285 => "1111000101111101",
44286 => "1111000101111110",
44287 => "1111000101111110",
44288 => "1111000101111111",
44289 => "1111000110000000",
44290 => "1111000110000001",
44291 => "1111000110000010",
44292 => "1111000110000011",
44293 => "1111000110000100",
44294 => "1111000110000100",
44295 => "1111000110000101",
44296 => "1111000110000110",
44297 => "1111000110000111",
44298 => "1111000110001000",
44299 => "1111000110001001",
44300 => "1111000110001010",
44301 => "1111000110001010",
44302 => "1111000110001011",
44303 => "1111000110001100",
44304 => "1111000110001101",
44305 => "1111000110001110",
44306 => "1111000110001111",
44307 => "1111000110010000",
44308 => "1111000110010000",
44309 => "1111000110010001",
44310 => "1111000110010010",
44311 => "1111000110010011",
44312 => "1111000110010100",
44313 => "1111000110010101",
44314 => "1111000110010101",
44315 => "1111000110010110",
44316 => "1111000110010111",
44317 => "1111000110011000",
44318 => "1111000110011001",
44319 => "1111000110011010",
44320 => "1111000110011011",
44321 => "1111000110011011",
44322 => "1111000110011100",
44323 => "1111000110011101",
44324 => "1111000110011110",
44325 => "1111000110011111",
44326 => "1111000110100000",
44327 => "1111000110100001",
44328 => "1111000110100001",
44329 => "1111000110100010",
44330 => "1111000110100011",
44331 => "1111000110100100",
44332 => "1111000110100101",
44333 => "1111000110100110",
44334 => "1111000110100110",
44335 => "1111000110100111",
44336 => "1111000110101000",
44337 => "1111000110101001",
44338 => "1111000110101010",
44339 => "1111000110101011",
44340 => "1111000110101100",
44341 => "1111000110101100",
44342 => "1111000110101101",
44343 => "1111000110101110",
44344 => "1111000110101111",
44345 => "1111000110110000",
44346 => "1111000110110001",
44347 => "1111000110110001",
44348 => "1111000110110010",
44349 => "1111000110110011",
44350 => "1111000110110100",
44351 => "1111000110110101",
44352 => "1111000110110110",
44353 => "1111000110110110",
44354 => "1111000110110111",
44355 => "1111000110111000",
44356 => "1111000110111001",
44357 => "1111000110111010",
44358 => "1111000110111011",
44359 => "1111000110111100",
44360 => "1111000110111100",
44361 => "1111000110111101",
44362 => "1111000110111110",
44363 => "1111000110111111",
44364 => "1111000111000000",
44365 => "1111000111000001",
44366 => "1111000111000001",
44367 => "1111000111000010",
44368 => "1111000111000011",
44369 => "1111000111000100",
44370 => "1111000111000101",
44371 => "1111000111000110",
44372 => "1111000111000110",
44373 => "1111000111000111",
44374 => "1111000111001000",
44375 => "1111000111001001",
44376 => "1111000111001010",
44377 => "1111000111001011",
44378 => "1111000111001100",
44379 => "1111000111001100",
44380 => "1111000111001101",
44381 => "1111000111001110",
44382 => "1111000111001111",
44383 => "1111000111010000",
44384 => "1111000111010001",
44385 => "1111000111010001",
44386 => "1111000111010010",
44387 => "1111000111010011",
44388 => "1111000111010100",
44389 => "1111000111010101",
44390 => "1111000111010110",
44391 => "1111000111010110",
44392 => "1111000111010111",
44393 => "1111000111011000",
44394 => "1111000111011001",
44395 => "1111000111011010",
44396 => "1111000111011011",
44397 => "1111000111011011",
44398 => "1111000111011100",
44399 => "1111000111011101",
44400 => "1111000111011110",
44401 => "1111000111011111",
44402 => "1111000111100000",
44403 => "1111000111100000",
44404 => "1111000111100001",
44405 => "1111000111100010",
44406 => "1111000111100011",
44407 => "1111000111100100",
44408 => "1111000111100101",
44409 => "1111000111100101",
44410 => "1111000111100110",
44411 => "1111000111100111",
44412 => "1111000111101000",
44413 => "1111000111101001",
44414 => "1111000111101010",
44415 => "1111000111101010",
44416 => "1111000111101011",
44417 => "1111000111101100",
44418 => "1111000111101101",
44419 => "1111000111101110",
44420 => "1111000111101111",
44421 => "1111000111101111",
44422 => "1111000111110000",
44423 => "1111000111110001",
44424 => "1111000111110010",
44425 => "1111000111110011",
44426 => "1111000111110100",
44427 => "1111000111110100",
44428 => "1111000111110101",
44429 => "1111000111110110",
44430 => "1111000111110111",
44431 => "1111000111111000",
44432 => "1111000111111001",
44433 => "1111000111111001",
44434 => "1111000111111010",
44435 => "1111000111111011",
44436 => "1111000111111100",
44437 => "1111000111111101",
44438 => "1111000111111101",
44439 => "1111000111111110",
44440 => "1111000111111111",
44441 => "1111001000000000",
44442 => "1111001000000001",
44443 => "1111001000000010",
44444 => "1111001000000010",
44445 => "1111001000000011",
44446 => "1111001000000100",
44447 => "1111001000000101",
44448 => "1111001000000110",
44449 => "1111001000000111",
44450 => "1111001000000111",
44451 => "1111001000001000",
44452 => "1111001000001001",
44453 => "1111001000001010",
44454 => "1111001000001011",
44455 => "1111001000001100",
44456 => "1111001000001100",
44457 => "1111001000001101",
44458 => "1111001000001110",
44459 => "1111001000001111",
44460 => "1111001000010000",
44461 => "1111001000010000",
44462 => "1111001000010001",
44463 => "1111001000010010",
44464 => "1111001000010011",
44465 => "1111001000010100",
44466 => "1111001000010101",
44467 => "1111001000010101",
44468 => "1111001000010110",
44469 => "1111001000010111",
44470 => "1111001000011000",
44471 => "1111001000011001",
44472 => "1111001000011010",
44473 => "1111001000011010",
44474 => "1111001000011011",
44475 => "1111001000011100",
44476 => "1111001000011101",
44477 => "1111001000011110",
44478 => "1111001000011110",
44479 => "1111001000011111",
44480 => "1111001000100000",
44481 => "1111001000100001",
44482 => "1111001000100010",
44483 => "1111001000100011",
44484 => "1111001000100011",
44485 => "1111001000100100",
44486 => "1111001000100101",
44487 => "1111001000100110",
44488 => "1111001000100111",
44489 => "1111001000100111",
44490 => "1111001000101000",
44491 => "1111001000101001",
44492 => "1111001000101010",
44493 => "1111001000101011",
44494 => "1111001000101100",
44495 => "1111001000101100",
44496 => "1111001000101101",
44497 => "1111001000101110",
44498 => "1111001000101111",
44499 => "1111001000110000",
44500 => "1111001000110000",
44501 => "1111001000110001",
44502 => "1111001000110010",
44503 => "1111001000110011",
44504 => "1111001000110100",
44505 => "1111001000110101",
44506 => "1111001000110101",
44507 => "1111001000110110",
44508 => "1111001000110111",
44509 => "1111001000111000",
44510 => "1111001000111001",
44511 => "1111001000111001",
44512 => "1111001000111010",
44513 => "1111001000111011",
44514 => "1111001000111100",
44515 => "1111001000111101",
44516 => "1111001000111101",
44517 => "1111001000111110",
44518 => "1111001000111111",
44519 => "1111001001000000",
44520 => "1111001001000001",
44521 => "1111001001000010",
44522 => "1111001001000010",
44523 => "1111001001000011",
44524 => "1111001001000100",
44525 => "1111001001000101",
44526 => "1111001001000110",
44527 => "1111001001000110",
44528 => "1111001001000111",
44529 => "1111001001001000",
44530 => "1111001001001001",
44531 => "1111001001001010",
44532 => "1111001001001010",
44533 => "1111001001001011",
44534 => "1111001001001100",
44535 => "1111001001001101",
44536 => "1111001001001110",
44537 => "1111001001001111",
44538 => "1111001001001111",
44539 => "1111001001010000",
44540 => "1111001001010001",
44541 => "1111001001010010",
44542 => "1111001001010011",
44543 => "1111001001010011",
44544 => "1111001001010100",
44545 => "1111001001010101",
44546 => "1111001001010110",
44547 => "1111001001010111",
44548 => "1111001001010111",
44549 => "1111001001011000",
44550 => "1111001001011001",
44551 => "1111001001011010",
44552 => "1111001001011011",
44553 => "1111001001011011",
44554 => "1111001001011100",
44555 => "1111001001011101",
44556 => "1111001001011110",
44557 => "1111001001011111",
44558 => "1111001001100000",
44559 => "1111001001100000",
44560 => "1111001001100001",
44561 => "1111001001100010",
44562 => "1111001001100011",
44563 => "1111001001100100",
44564 => "1111001001100100",
44565 => "1111001001100101",
44566 => "1111001001100110",
44567 => "1111001001100111",
44568 => "1111001001101000",
44569 => "1111001001101000",
44570 => "1111001001101001",
44571 => "1111001001101010",
44572 => "1111001001101011",
44573 => "1111001001101100",
44574 => "1111001001101100",
44575 => "1111001001101101",
44576 => "1111001001101110",
44577 => "1111001001101111",
44578 => "1111001001110000",
44579 => "1111001001110000",
44580 => "1111001001110001",
44581 => "1111001001110010",
44582 => "1111001001110011",
44583 => "1111001001110100",
44584 => "1111001001110100",
44585 => "1111001001110101",
44586 => "1111001001110110",
44587 => "1111001001110111",
44588 => "1111001001111000",
44589 => "1111001001111000",
44590 => "1111001001111001",
44591 => "1111001001111010",
44592 => "1111001001111011",
44593 => "1111001001111100",
44594 => "1111001001111100",
44595 => "1111001001111101",
44596 => "1111001001111110",
44597 => "1111001001111111",
44598 => "1111001010000000",
44599 => "1111001010000000",
44600 => "1111001010000001",
44601 => "1111001010000010",
44602 => "1111001010000011",
44603 => "1111001010000100",
44604 => "1111001010000100",
44605 => "1111001010000101",
44606 => "1111001010000110",
44607 => "1111001010000111",
44608 => "1111001010001000",
44609 => "1111001010001000",
44610 => "1111001010001001",
44611 => "1111001010001010",
44612 => "1111001010001011",
44613 => "1111001010001100",
44614 => "1111001010001100",
44615 => "1111001010001101",
44616 => "1111001010001110",
44617 => "1111001010001111",
44618 => "1111001010010000",
44619 => "1111001010010000",
44620 => "1111001010010001",
44621 => "1111001010010010",
44622 => "1111001010010011",
44623 => "1111001010010100",
44624 => "1111001010010100",
44625 => "1111001010010101",
44626 => "1111001010010110",
44627 => "1111001010010111",
44628 => "1111001010011000",
44629 => "1111001010011000",
44630 => "1111001010011001",
44631 => "1111001010011010",
44632 => "1111001010011011",
44633 => "1111001010011011",
44634 => "1111001010011100",
44635 => "1111001010011101",
44636 => "1111001010011110",
44637 => "1111001010011111",
44638 => "1111001010011111",
44639 => "1111001010100000",
44640 => "1111001010100001",
44641 => "1111001010100010",
44642 => "1111001010100011",
44643 => "1111001010100011",
44644 => "1111001010100100",
44645 => "1111001010100101",
44646 => "1111001010100110",
44647 => "1111001010100111",
44648 => "1111001010100111",
44649 => "1111001010101000",
44650 => "1111001010101001",
44651 => "1111001010101010",
44652 => "1111001010101011",
44653 => "1111001010101011",
44654 => "1111001010101100",
44655 => "1111001010101101",
44656 => "1111001010101110",
44657 => "1111001010101110",
44658 => "1111001010101111",
44659 => "1111001010110000",
44660 => "1111001010110001",
44661 => "1111001010110010",
44662 => "1111001010110010",
44663 => "1111001010110011",
44664 => "1111001010110100",
44665 => "1111001010110101",
44666 => "1111001010110110",
44667 => "1111001010110110",
44668 => "1111001010110111",
44669 => "1111001010111000",
44670 => "1111001010111001",
44671 => "1111001010111010",
44672 => "1111001010111010",
44673 => "1111001010111011",
44674 => "1111001010111100",
44675 => "1111001010111101",
44676 => "1111001010111101",
44677 => "1111001010111110",
44678 => "1111001010111111",
44679 => "1111001011000000",
44680 => "1111001011000001",
44681 => "1111001011000001",
44682 => "1111001011000010",
44683 => "1111001011000011",
44684 => "1111001011000100",
44685 => "1111001011000101",
44686 => "1111001011000101",
44687 => "1111001011000110",
44688 => "1111001011000111",
44689 => "1111001011001000",
44690 => "1111001011001000",
44691 => "1111001011001001",
44692 => "1111001011001010",
44693 => "1111001011001011",
44694 => "1111001011001100",
44695 => "1111001011001100",
44696 => "1111001011001101",
44697 => "1111001011001110",
44698 => "1111001011001111",
44699 => "1111001011001111",
44700 => "1111001011010000",
44701 => "1111001011010001",
44702 => "1111001011010010",
44703 => "1111001011010011",
44704 => "1111001011010011",
44705 => "1111001011010100",
44706 => "1111001011010101",
44707 => "1111001011010110",
44708 => "1111001011010110",
44709 => "1111001011010111",
44710 => "1111001011011000",
44711 => "1111001011011001",
44712 => "1111001011011010",
44713 => "1111001011011010",
44714 => "1111001011011011",
44715 => "1111001011011100",
44716 => "1111001011011101",
44717 => "1111001011011110",
44718 => "1111001011011110",
44719 => "1111001011011111",
44720 => "1111001011100000",
44721 => "1111001011100001",
44722 => "1111001011100001",
44723 => "1111001011100010",
44724 => "1111001011100011",
44725 => "1111001011100100",
44726 => "1111001011100101",
44727 => "1111001011100101",
44728 => "1111001011100110",
44729 => "1111001011100111",
44730 => "1111001011101000",
44731 => "1111001011101000",
44732 => "1111001011101001",
44733 => "1111001011101010",
44734 => "1111001011101011",
44735 => "1111001011101011",
44736 => "1111001011101100",
44737 => "1111001011101101",
44738 => "1111001011101110",
44739 => "1111001011101111",
44740 => "1111001011101111",
44741 => "1111001011110000",
44742 => "1111001011110001",
44743 => "1111001011110010",
44744 => "1111001011110010",
44745 => "1111001011110011",
44746 => "1111001011110100",
44747 => "1111001011110101",
44748 => "1111001011110110",
44749 => "1111001011110110",
44750 => "1111001011110111",
44751 => "1111001011111000",
44752 => "1111001011111001",
44753 => "1111001011111001",
44754 => "1111001011111010",
44755 => "1111001011111011",
44756 => "1111001011111100",
44757 => "1111001011111101",
44758 => "1111001011111101",
44759 => "1111001011111110",
44760 => "1111001011111111",
44761 => "1111001100000000",
44762 => "1111001100000000",
44763 => "1111001100000001",
44764 => "1111001100000010",
44765 => "1111001100000011",
44766 => "1111001100000011",
44767 => "1111001100000100",
44768 => "1111001100000101",
44769 => "1111001100000110",
44770 => "1111001100000111",
44771 => "1111001100000111",
44772 => "1111001100001000",
44773 => "1111001100001001",
44774 => "1111001100001010",
44775 => "1111001100001010",
44776 => "1111001100001011",
44777 => "1111001100001100",
44778 => "1111001100001101",
44779 => "1111001100001101",
44780 => "1111001100001110",
44781 => "1111001100001111",
44782 => "1111001100010000",
44783 => "1111001100010001",
44784 => "1111001100010001",
44785 => "1111001100010010",
44786 => "1111001100010011",
44787 => "1111001100010100",
44788 => "1111001100010100",
44789 => "1111001100010101",
44790 => "1111001100010110",
44791 => "1111001100010111",
44792 => "1111001100010111",
44793 => "1111001100011000",
44794 => "1111001100011001",
44795 => "1111001100011010",
44796 => "1111001100011010",
44797 => "1111001100011011",
44798 => "1111001100011100",
44799 => "1111001100011101",
44800 => "1111001100011110",
44801 => "1111001100011110",
44802 => "1111001100011111",
44803 => "1111001100100000",
44804 => "1111001100100001",
44805 => "1111001100100001",
44806 => "1111001100100010",
44807 => "1111001100100011",
44808 => "1111001100100100",
44809 => "1111001100100100",
44810 => "1111001100100101",
44811 => "1111001100100110",
44812 => "1111001100100111",
44813 => "1111001100100111",
44814 => "1111001100101000",
44815 => "1111001100101001",
44816 => "1111001100101010",
44817 => "1111001100101011",
44818 => "1111001100101011",
44819 => "1111001100101100",
44820 => "1111001100101101",
44821 => "1111001100101110",
44822 => "1111001100101110",
44823 => "1111001100101111",
44824 => "1111001100110000",
44825 => "1111001100110001",
44826 => "1111001100110001",
44827 => "1111001100110010",
44828 => "1111001100110011",
44829 => "1111001100110100",
44830 => "1111001100110100",
44831 => "1111001100110101",
44832 => "1111001100110110",
44833 => "1111001100110111",
44834 => "1111001100110111",
44835 => "1111001100111000",
44836 => "1111001100111001",
44837 => "1111001100111010",
44838 => "1111001100111010",
44839 => "1111001100111011",
44840 => "1111001100111100",
44841 => "1111001100111101",
44842 => "1111001100111110",
44843 => "1111001100111110",
44844 => "1111001100111111",
44845 => "1111001101000000",
44846 => "1111001101000001",
44847 => "1111001101000001",
44848 => "1111001101000010",
44849 => "1111001101000011",
44850 => "1111001101000100",
44851 => "1111001101000100",
44852 => "1111001101000101",
44853 => "1111001101000110",
44854 => "1111001101000111",
44855 => "1111001101000111",
44856 => "1111001101001000",
44857 => "1111001101001001",
44858 => "1111001101001010",
44859 => "1111001101001010",
44860 => "1111001101001011",
44861 => "1111001101001100",
44862 => "1111001101001101",
44863 => "1111001101001101",
44864 => "1111001101001110",
44865 => "1111001101001111",
44866 => "1111001101010000",
44867 => "1111001101010000",
44868 => "1111001101010001",
44869 => "1111001101010010",
44870 => "1111001101010011",
44871 => "1111001101010011",
44872 => "1111001101010100",
44873 => "1111001101010101",
44874 => "1111001101010110",
44875 => "1111001101010110",
44876 => "1111001101010111",
44877 => "1111001101011000",
44878 => "1111001101011001",
44879 => "1111001101011001",
44880 => "1111001101011010",
44881 => "1111001101011011",
44882 => "1111001101011100",
44883 => "1111001101011100",
44884 => "1111001101011101",
44885 => "1111001101011110",
44886 => "1111001101011111",
44887 => "1111001101011111",
44888 => "1111001101100000",
44889 => "1111001101100001",
44890 => "1111001101100010",
44891 => "1111001101100010",
44892 => "1111001101100011",
44893 => "1111001101100100",
44894 => "1111001101100101",
44895 => "1111001101100101",
44896 => "1111001101100110",
44897 => "1111001101100111",
44898 => "1111001101101000",
44899 => "1111001101101000",
44900 => "1111001101101001",
44901 => "1111001101101010",
44902 => "1111001101101011",
44903 => "1111001101101011",
44904 => "1111001101101100",
44905 => "1111001101101101",
44906 => "1111001101101110",
44907 => "1111001101101110",
44908 => "1111001101101111",
44909 => "1111001101110000",
44910 => "1111001101110001",
44911 => "1111001101110001",
44912 => "1111001101110010",
44913 => "1111001101110011",
44914 => "1111001101110100",
44915 => "1111001101110100",
44916 => "1111001101110101",
44917 => "1111001101110110",
44918 => "1111001101110111",
44919 => "1111001101110111",
44920 => "1111001101111000",
44921 => "1111001101111001",
44922 => "1111001101111010",
44923 => "1111001101111010",
44924 => "1111001101111011",
44925 => "1111001101111100",
44926 => "1111001101111101",
44927 => "1111001101111101",
44928 => "1111001101111110",
44929 => "1111001101111111",
44930 => "1111001110000000",
44931 => "1111001110000000",
44932 => "1111001110000001",
44933 => "1111001110000010",
44934 => "1111001110000011",
44935 => "1111001110000011",
44936 => "1111001110000100",
44937 => "1111001110000101",
44938 => "1111001110000101",
44939 => "1111001110000110",
44940 => "1111001110000111",
44941 => "1111001110001000",
44942 => "1111001110001000",
44943 => "1111001110001001",
44944 => "1111001110001010",
44945 => "1111001110001011",
44946 => "1111001110001011",
44947 => "1111001110001100",
44948 => "1111001110001101",
44949 => "1111001110001110",
44950 => "1111001110001110",
44951 => "1111001110001111",
44952 => "1111001110010000",
44953 => "1111001110010001",
44954 => "1111001110010001",
44955 => "1111001110010010",
44956 => "1111001110010011",
44957 => "1111001110010100",
44958 => "1111001110010100",
44959 => "1111001110010101",
44960 => "1111001110010110",
44961 => "1111001110010111",
44962 => "1111001110010111",
44963 => "1111001110011000",
44964 => "1111001110011001",
44965 => "1111001110011001",
44966 => "1111001110011010",
44967 => "1111001110011011",
44968 => "1111001110011100",
44969 => "1111001110011100",
44970 => "1111001110011101",
44971 => "1111001110011110",
44972 => "1111001110011111",
44973 => "1111001110011111",
44974 => "1111001110100000",
44975 => "1111001110100001",
44976 => "1111001110100010",
44977 => "1111001110100010",
44978 => "1111001110100011",
44979 => "1111001110100100",
44980 => "1111001110100101",
44981 => "1111001110100101",
44982 => "1111001110100110",
44983 => "1111001110100111",
44984 => "1111001110100111",
44985 => "1111001110101000",
44986 => "1111001110101001",
44987 => "1111001110101010",
44988 => "1111001110101010",
44989 => "1111001110101011",
44990 => "1111001110101100",
44991 => "1111001110101101",
44992 => "1111001110101101",
44993 => "1111001110101110",
44994 => "1111001110101111",
44995 => "1111001110110000",
44996 => "1111001110110000",
44997 => "1111001110110001",
44998 => "1111001110110010",
44999 => "1111001110110010",
45000 => "1111001110110011",
45001 => "1111001110110100",
45002 => "1111001110110101",
45003 => "1111001110110101",
45004 => "1111001110110110",
45005 => "1111001110110111",
45006 => "1111001110111000",
45007 => "1111001110111000",
45008 => "1111001110111001",
45009 => "1111001110111010",
45010 => "1111001110111010",
45011 => "1111001110111011",
45012 => "1111001110111100",
45013 => "1111001110111101",
45014 => "1111001110111101",
45015 => "1111001110111110",
45016 => "1111001110111111",
45017 => "1111001111000000",
45018 => "1111001111000000",
45019 => "1111001111000001",
45020 => "1111001111000010",
45021 => "1111001111000011",
45022 => "1111001111000011",
45023 => "1111001111000100",
45024 => "1111001111000101",
45025 => "1111001111000101",
45026 => "1111001111000110",
45027 => "1111001111000111",
45028 => "1111001111001000",
45029 => "1111001111001000",
45030 => "1111001111001001",
45031 => "1111001111001010",
45032 => "1111001111001011",
45033 => "1111001111001011",
45034 => "1111001111001100",
45035 => "1111001111001101",
45036 => "1111001111001101",
45037 => "1111001111001110",
45038 => "1111001111001111",
45039 => "1111001111010000",
45040 => "1111001111010000",
45041 => "1111001111010001",
45042 => "1111001111010010",
45043 => "1111001111010010",
45044 => "1111001111010011",
45045 => "1111001111010100",
45046 => "1111001111010101",
45047 => "1111001111010101",
45048 => "1111001111010110",
45049 => "1111001111010111",
45050 => "1111001111011000",
45051 => "1111001111011000",
45052 => "1111001111011001",
45053 => "1111001111011010",
45054 => "1111001111011010",
45055 => "1111001111011011",
45056 => "1111001111011100",
45057 => "1111001111011101",
45058 => "1111001111011101",
45059 => "1111001111011110",
45060 => "1111001111011111",
45061 => "1111001111100000",
45062 => "1111001111100000",
45063 => "1111001111100001",
45064 => "1111001111100010",
45065 => "1111001111100010",
45066 => "1111001111100011",
45067 => "1111001111100100",
45068 => "1111001111100101",
45069 => "1111001111100101",
45070 => "1111001111100110",
45071 => "1111001111100111",
45072 => "1111001111100111",
45073 => "1111001111101000",
45074 => "1111001111101001",
45075 => "1111001111101010",
45076 => "1111001111101010",
45077 => "1111001111101011",
45078 => "1111001111101100",
45079 => "1111001111101100",
45080 => "1111001111101101",
45081 => "1111001111101110",
45082 => "1111001111101111",
45083 => "1111001111101111",
45084 => "1111001111110000",
45085 => "1111001111110001",
45086 => "1111001111110010",
45087 => "1111001111110010",
45088 => "1111001111110011",
45089 => "1111001111110100",
45090 => "1111001111110100",
45091 => "1111001111110101",
45092 => "1111001111110110",
45093 => "1111001111110111",
45094 => "1111001111110111",
45095 => "1111001111111000",
45096 => "1111001111111001",
45097 => "1111001111111001",
45098 => "1111001111111010",
45099 => "1111001111111011",
45100 => "1111001111111100",
45101 => "1111001111111100",
45102 => "1111001111111101",
45103 => "1111001111111110",
45104 => "1111001111111110",
45105 => "1111001111111111",
45106 => "1111010000000000",
45107 => "1111010000000001",
45108 => "1111010000000001",
45109 => "1111010000000010",
45110 => "1111010000000011",
45111 => "1111010000000011",
45112 => "1111010000000100",
45113 => "1111010000000101",
45114 => "1111010000000110",
45115 => "1111010000000110",
45116 => "1111010000000111",
45117 => "1111010000001000",
45118 => "1111010000001000",
45119 => "1111010000001001",
45120 => "1111010000001010",
45121 => "1111010000001011",
45122 => "1111010000001011",
45123 => "1111010000001100",
45124 => "1111010000001101",
45125 => "1111010000001101",
45126 => "1111010000001110",
45127 => "1111010000001111",
45128 => "1111010000010000",
45129 => "1111010000010000",
45130 => "1111010000010001",
45131 => "1111010000010010",
45132 => "1111010000010010",
45133 => "1111010000010011",
45134 => "1111010000010100",
45135 => "1111010000010100",
45136 => "1111010000010101",
45137 => "1111010000010110",
45138 => "1111010000010111",
45139 => "1111010000010111",
45140 => "1111010000011000",
45141 => "1111010000011001",
45142 => "1111010000011001",
45143 => "1111010000011010",
45144 => "1111010000011011",
45145 => "1111010000011100",
45146 => "1111010000011100",
45147 => "1111010000011101",
45148 => "1111010000011110",
45149 => "1111010000011110",
45150 => "1111010000011111",
45151 => "1111010000100000",
45152 => "1111010000100001",
45153 => "1111010000100001",
45154 => "1111010000100010",
45155 => "1111010000100011",
45156 => "1111010000100011",
45157 => "1111010000100100",
45158 => "1111010000100101",
45159 => "1111010000100101",
45160 => "1111010000100110",
45161 => "1111010000100111",
45162 => "1111010000101000",
45163 => "1111010000101000",
45164 => "1111010000101001",
45165 => "1111010000101010",
45166 => "1111010000101010",
45167 => "1111010000101011",
45168 => "1111010000101100",
45169 => "1111010000101101",
45170 => "1111010000101101",
45171 => "1111010000101110",
45172 => "1111010000101111",
45173 => "1111010000101111",
45174 => "1111010000110000",
45175 => "1111010000110001",
45176 => "1111010000110001",
45177 => "1111010000110010",
45178 => "1111010000110011",
45179 => "1111010000110100",
45180 => "1111010000110100",
45181 => "1111010000110101",
45182 => "1111010000110110",
45183 => "1111010000110110",
45184 => "1111010000110111",
45185 => "1111010000111000",
45186 => "1111010000111001",
45187 => "1111010000111001",
45188 => "1111010000111010",
45189 => "1111010000111011",
45190 => "1111010000111011",
45191 => "1111010000111100",
45192 => "1111010000111101",
45193 => "1111010000111101",
45194 => "1111010000111110",
45195 => "1111010000111111",
45196 => "1111010001000000",
45197 => "1111010001000000",
45198 => "1111010001000001",
45199 => "1111010001000010",
45200 => "1111010001000010",
45201 => "1111010001000011",
45202 => "1111010001000100",
45203 => "1111010001000100",
45204 => "1111010001000101",
45205 => "1111010001000110",
45206 => "1111010001000111",
45207 => "1111010001000111",
45208 => "1111010001001000",
45209 => "1111010001001001",
45210 => "1111010001001001",
45211 => "1111010001001010",
45212 => "1111010001001011",
45213 => "1111010001001011",
45214 => "1111010001001100",
45215 => "1111010001001101",
45216 => "1111010001001110",
45217 => "1111010001001110",
45218 => "1111010001001111",
45219 => "1111010001010000",
45220 => "1111010001010000",
45221 => "1111010001010001",
45222 => "1111010001010010",
45223 => "1111010001010010",
45224 => "1111010001010011",
45225 => "1111010001010100",
45226 => "1111010001010100",
45227 => "1111010001010101",
45228 => "1111010001010110",
45229 => "1111010001010111",
45230 => "1111010001010111",
45231 => "1111010001011000",
45232 => "1111010001011001",
45233 => "1111010001011001",
45234 => "1111010001011010",
45235 => "1111010001011011",
45236 => "1111010001011011",
45237 => "1111010001011100",
45238 => "1111010001011101",
45239 => "1111010001011110",
45240 => "1111010001011110",
45241 => "1111010001011111",
45242 => "1111010001100000",
45243 => "1111010001100000",
45244 => "1111010001100001",
45245 => "1111010001100010",
45246 => "1111010001100010",
45247 => "1111010001100011",
45248 => "1111010001100100",
45249 => "1111010001100100",
45250 => "1111010001100101",
45251 => "1111010001100110",
45252 => "1111010001100111",
45253 => "1111010001100111",
45254 => "1111010001101000",
45255 => "1111010001101001",
45256 => "1111010001101001",
45257 => "1111010001101010",
45258 => "1111010001101011",
45259 => "1111010001101011",
45260 => "1111010001101100",
45261 => "1111010001101101",
45262 => "1111010001101101",
45263 => "1111010001101110",
45264 => "1111010001101111",
45265 => "1111010001110000",
45266 => "1111010001110000",
45267 => "1111010001110001",
45268 => "1111010001110010",
45269 => "1111010001110010",
45270 => "1111010001110011",
45271 => "1111010001110100",
45272 => "1111010001110100",
45273 => "1111010001110101",
45274 => "1111010001110110",
45275 => "1111010001110110",
45276 => "1111010001110111",
45277 => "1111010001111000",
45278 => "1111010001111000",
45279 => "1111010001111001",
45280 => "1111010001111010",
45281 => "1111010001111011",
45282 => "1111010001111011",
45283 => "1111010001111100",
45284 => "1111010001111101",
45285 => "1111010001111101",
45286 => "1111010001111110",
45287 => "1111010001111111",
45288 => "1111010001111111",
45289 => "1111010010000000",
45290 => "1111010010000001",
45291 => "1111010010000001",
45292 => "1111010010000010",
45293 => "1111010010000011",
45294 => "1111010010000011",
45295 => "1111010010000100",
45296 => "1111010010000101",
45297 => "1111010010000110",
45298 => "1111010010000110",
45299 => "1111010010000111",
45300 => "1111010010001000",
45301 => "1111010010001000",
45302 => "1111010010001001",
45303 => "1111010010001010",
45304 => "1111010010001010",
45305 => "1111010010001011",
45306 => "1111010010001100",
45307 => "1111010010001100",
45308 => "1111010010001101",
45309 => "1111010010001110",
45310 => "1111010010001110",
45311 => "1111010010001111",
45312 => "1111010010010000",
45313 => "1111010010010000",
45314 => "1111010010010001",
45315 => "1111010010010010",
45316 => "1111010010010010",
45317 => "1111010010010011",
45318 => "1111010010010100",
45319 => "1111010010010101",
45320 => "1111010010010101",
45321 => "1111010010010110",
45322 => "1111010010010111",
45323 => "1111010010010111",
45324 => "1111010010011000",
45325 => "1111010010011001",
45326 => "1111010010011001",
45327 => "1111010010011010",
45328 => "1111010010011011",
45329 => "1111010010011011",
45330 => "1111010010011100",
45331 => "1111010010011101",
45332 => "1111010010011101",
45333 => "1111010010011110",
45334 => "1111010010011111",
45335 => "1111010010011111",
45336 => "1111010010100000",
45337 => "1111010010100001",
45338 => "1111010010100001",
45339 => "1111010010100010",
45340 => "1111010010100011",
45341 => "1111010010100100",
45342 => "1111010010100100",
45343 => "1111010010100101",
45344 => "1111010010100110",
45345 => "1111010010100110",
45346 => "1111010010100111",
45347 => "1111010010101000",
45348 => "1111010010101000",
45349 => "1111010010101001",
45350 => "1111010010101010",
45351 => "1111010010101010",
45352 => "1111010010101011",
45353 => "1111010010101100",
45354 => "1111010010101100",
45355 => "1111010010101101",
45356 => "1111010010101110",
45357 => "1111010010101110",
45358 => "1111010010101111",
45359 => "1111010010110000",
45360 => "1111010010110000",
45361 => "1111010010110001",
45362 => "1111010010110010",
45363 => "1111010010110010",
45364 => "1111010010110011",
45365 => "1111010010110100",
45366 => "1111010010110100",
45367 => "1111010010110101",
45368 => "1111010010110110",
45369 => "1111010010110110",
45370 => "1111010010110111",
45371 => "1111010010111000",
45372 => "1111010010111000",
45373 => "1111010010111001",
45374 => "1111010010111010",
45375 => "1111010010111010",
45376 => "1111010010111011",
45377 => "1111010010111100",
45378 => "1111010010111101",
45379 => "1111010010111101",
45380 => "1111010010111110",
45381 => "1111010010111111",
45382 => "1111010010111111",
45383 => "1111010011000000",
45384 => "1111010011000001",
45385 => "1111010011000001",
45386 => "1111010011000010",
45387 => "1111010011000011",
45388 => "1111010011000011",
45389 => "1111010011000100",
45390 => "1111010011000101",
45391 => "1111010011000101",
45392 => "1111010011000110",
45393 => "1111010011000111",
45394 => "1111010011000111",
45395 => "1111010011001000",
45396 => "1111010011001001",
45397 => "1111010011001001",
45398 => "1111010011001010",
45399 => "1111010011001011",
45400 => "1111010011001011",
45401 => "1111010011001100",
45402 => "1111010011001101",
45403 => "1111010011001101",
45404 => "1111010011001110",
45405 => "1111010011001111",
45406 => "1111010011001111",
45407 => "1111010011010000",
45408 => "1111010011010001",
45409 => "1111010011010001",
45410 => "1111010011010010",
45411 => "1111010011010011",
45412 => "1111010011010011",
45413 => "1111010011010100",
45414 => "1111010011010101",
45415 => "1111010011010101",
45416 => "1111010011010110",
45417 => "1111010011010111",
45418 => "1111010011010111",
45419 => "1111010011011000",
45420 => "1111010011011001",
45421 => "1111010011011001",
45422 => "1111010011011010",
45423 => "1111010011011011",
45424 => "1111010011011011",
45425 => "1111010011011100",
45426 => "1111010011011101",
45427 => "1111010011011101",
45428 => "1111010011011110",
45429 => "1111010011011111",
45430 => "1111010011011111",
45431 => "1111010011100000",
45432 => "1111010011100001",
45433 => "1111010011100001",
45434 => "1111010011100010",
45435 => "1111010011100011",
45436 => "1111010011100011",
45437 => "1111010011100100",
45438 => "1111010011100101",
45439 => "1111010011100101",
45440 => "1111010011100110",
45441 => "1111010011100111",
45442 => "1111010011100111",
45443 => "1111010011101000",
45444 => "1111010011101001",
45445 => "1111010011101001",
45446 => "1111010011101010",
45447 => "1111010011101011",
45448 => "1111010011101011",
45449 => "1111010011101100",
45450 => "1111010011101101",
45451 => "1111010011101101",
45452 => "1111010011101110",
45453 => "1111010011101111",
45454 => "1111010011101111",
45455 => "1111010011110000",
45456 => "1111010011110001",
45457 => "1111010011110001",
45458 => "1111010011110010",
45459 => "1111010011110011",
45460 => "1111010011110011",
45461 => "1111010011110100",
45462 => "1111010011110101",
45463 => "1111010011110101",
45464 => "1111010011110110",
45465 => "1111010011110110",
45466 => "1111010011110111",
45467 => "1111010011111000",
45468 => "1111010011111000",
45469 => "1111010011111001",
45470 => "1111010011111010",
45471 => "1111010011111010",
45472 => "1111010011111011",
45473 => "1111010011111100",
45474 => "1111010011111100",
45475 => "1111010011111101",
45476 => "1111010011111110",
45477 => "1111010011111110",
45478 => "1111010011111111",
45479 => "1111010100000000",
45480 => "1111010100000000",
45481 => "1111010100000001",
45482 => "1111010100000010",
45483 => "1111010100000010",
45484 => "1111010100000011",
45485 => "1111010100000100",
45486 => "1111010100000100",
45487 => "1111010100000101",
45488 => "1111010100000110",
45489 => "1111010100000110",
45490 => "1111010100000111",
45491 => "1111010100001000",
45492 => "1111010100001000",
45493 => "1111010100001001",
45494 => "1111010100001010",
45495 => "1111010100001010",
45496 => "1111010100001011",
45497 => "1111010100001100",
45498 => "1111010100001100",
45499 => "1111010100001101",
45500 => "1111010100001101",
45501 => "1111010100001110",
45502 => "1111010100001111",
45503 => "1111010100001111",
45504 => "1111010100010000",
45505 => "1111010100010001",
45506 => "1111010100010001",
45507 => "1111010100010010",
45508 => "1111010100010011",
45509 => "1111010100010011",
45510 => "1111010100010100",
45511 => "1111010100010101",
45512 => "1111010100010101",
45513 => "1111010100010110",
45514 => "1111010100010111",
45515 => "1111010100010111",
45516 => "1111010100011000",
45517 => "1111010100011001",
45518 => "1111010100011001",
45519 => "1111010100011010",
45520 => "1111010100011011",
45521 => "1111010100011011",
45522 => "1111010100011100",
45523 => "1111010100011101",
45524 => "1111010100011101",
45525 => "1111010100011110",
45526 => "1111010100011110",
45527 => "1111010100011111",
45528 => "1111010100100000",
45529 => "1111010100100000",
45530 => "1111010100100001",
45531 => "1111010100100010",
45532 => "1111010100100010",
45533 => "1111010100100011",
45534 => "1111010100100100",
45535 => "1111010100100100",
45536 => "1111010100100101",
45537 => "1111010100100110",
45538 => "1111010100100110",
45539 => "1111010100100111",
45540 => "1111010100101000",
45541 => "1111010100101000",
45542 => "1111010100101001",
45543 => "1111010100101010",
45544 => "1111010100101010",
45545 => "1111010100101011",
45546 => "1111010100101011",
45547 => "1111010100101100",
45548 => "1111010100101101",
45549 => "1111010100101101",
45550 => "1111010100101110",
45551 => "1111010100101111",
45552 => "1111010100101111",
45553 => "1111010100110000",
45554 => "1111010100110001",
45555 => "1111010100110001",
45556 => "1111010100110010",
45557 => "1111010100110011",
45558 => "1111010100110011",
45559 => "1111010100110100",
45560 => "1111010100110101",
45561 => "1111010100110101",
45562 => "1111010100110110",
45563 => "1111010100110110",
45564 => "1111010100110111",
45565 => "1111010100111000",
45566 => "1111010100111000",
45567 => "1111010100111001",
45568 => "1111010100111010",
45569 => "1111010100111010",
45570 => "1111010100111011",
45571 => "1111010100111100",
45572 => "1111010100111100",
45573 => "1111010100111101",
45574 => "1111010100111110",
45575 => "1111010100111110",
45576 => "1111010100111111",
45577 => "1111010100111111",
45578 => "1111010101000000",
45579 => "1111010101000001",
45580 => "1111010101000001",
45581 => "1111010101000010",
45582 => "1111010101000011",
45583 => "1111010101000011",
45584 => "1111010101000100",
45585 => "1111010101000101",
45586 => "1111010101000101",
45587 => "1111010101000110",
45588 => "1111010101000111",
45589 => "1111010101000111",
45590 => "1111010101001000",
45591 => "1111010101001000",
45592 => "1111010101001001",
45593 => "1111010101001010",
45594 => "1111010101001010",
45595 => "1111010101001011",
45596 => "1111010101001100",
45597 => "1111010101001100",
45598 => "1111010101001101",
45599 => "1111010101001110",
45600 => "1111010101001110",
45601 => "1111010101001111",
45602 => "1111010101010000",
45603 => "1111010101010000",
45604 => "1111010101010001",
45605 => "1111010101010001",
45606 => "1111010101010010",
45607 => "1111010101010011",
45608 => "1111010101010011",
45609 => "1111010101010100",
45610 => "1111010101010101",
45611 => "1111010101010101",
45612 => "1111010101010110",
45613 => "1111010101010111",
45614 => "1111010101010111",
45615 => "1111010101011000",
45616 => "1111010101011000",
45617 => "1111010101011001",
45618 => "1111010101011010",
45619 => "1111010101011010",
45620 => "1111010101011011",
45621 => "1111010101011100",
45622 => "1111010101011100",
45623 => "1111010101011101",
45624 => "1111010101011110",
45625 => "1111010101011110",
45626 => "1111010101011111",
45627 => "1111010101011111",
45628 => "1111010101100000",
45629 => "1111010101100001",
45630 => "1111010101100001",
45631 => "1111010101100010",
45632 => "1111010101100011",
45633 => "1111010101100011",
45634 => "1111010101100100",
45635 => "1111010101100101",
45636 => "1111010101100101",
45637 => "1111010101100110",
45638 => "1111010101100110",
45639 => "1111010101100111",
45640 => "1111010101101000",
45641 => "1111010101101000",
45642 => "1111010101101001",
45643 => "1111010101101010",
45644 => "1111010101101010",
45645 => "1111010101101011",
45646 => "1111010101101100",
45647 => "1111010101101100",
45648 => "1111010101101101",
45649 => "1111010101101101",
45650 => "1111010101101110",
45651 => "1111010101101111",
45652 => "1111010101101111",
45653 => "1111010101110000",
45654 => "1111010101110001",
45655 => "1111010101110001",
45656 => "1111010101110010",
45657 => "1111010101110011",
45658 => "1111010101110011",
45659 => "1111010101110100",
45660 => "1111010101110100",
45661 => "1111010101110101",
45662 => "1111010101110110",
45663 => "1111010101110110",
45664 => "1111010101110111",
45665 => "1111010101111000",
45666 => "1111010101111000",
45667 => "1111010101111001",
45668 => "1111010101111001",
45669 => "1111010101111010",
45670 => "1111010101111011",
45671 => "1111010101111011",
45672 => "1111010101111100",
45673 => "1111010101111101",
45674 => "1111010101111101",
45675 => "1111010101111110",
45676 => "1111010101111111",
45677 => "1111010101111111",
45678 => "1111010110000000",
45679 => "1111010110000000",
45680 => "1111010110000001",
45681 => "1111010110000010",
45682 => "1111010110000010",
45683 => "1111010110000011",
45684 => "1111010110000100",
45685 => "1111010110000100",
45686 => "1111010110000101",
45687 => "1111010110000101",
45688 => "1111010110000110",
45689 => "1111010110000111",
45690 => "1111010110000111",
45691 => "1111010110001000",
45692 => "1111010110001001",
45693 => "1111010110001001",
45694 => "1111010110001010",
45695 => "1111010110001010",
45696 => "1111010110001011",
45697 => "1111010110001100",
45698 => "1111010110001100",
45699 => "1111010110001101",
45700 => "1111010110001110",
45701 => "1111010110001110",
45702 => "1111010110001111",
45703 => "1111010110001111",
45704 => "1111010110010000",
45705 => "1111010110010001",
45706 => "1111010110010001",
45707 => "1111010110010010",
45708 => "1111010110010011",
45709 => "1111010110010011",
45710 => "1111010110010100",
45711 => "1111010110010100",
45712 => "1111010110010101",
45713 => "1111010110010110",
45714 => "1111010110010110",
45715 => "1111010110010111",
45716 => "1111010110011000",
45717 => "1111010110011000",
45718 => "1111010110011001",
45719 => "1111010110011001",
45720 => "1111010110011010",
45721 => "1111010110011011",
45722 => "1111010110011011",
45723 => "1111010110011100",
45724 => "1111010110011101",
45725 => "1111010110011101",
45726 => "1111010110011110",
45727 => "1111010110011110",
45728 => "1111010110011111",
45729 => "1111010110100000",
45730 => "1111010110100000",
45731 => "1111010110100001",
45732 => "1111010110100010",
45733 => "1111010110100010",
45734 => "1111010110100011",
45735 => "1111010110100011",
45736 => "1111010110100100",
45737 => "1111010110100101",
45738 => "1111010110100101",
45739 => "1111010110100110",
45740 => "1111010110100111",
45741 => "1111010110100111",
45742 => "1111010110101000",
45743 => "1111010110101000",
45744 => "1111010110101001",
45745 => "1111010110101010",
45746 => "1111010110101010",
45747 => "1111010110101011",
45748 => "1111010110101011",
45749 => "1111010110101100",
45750 => "1111010110101101",
45751 => "1111010110101101",
45752 => "1111010110101110",
45753 => "1111010110101111",
45754 => "1111010110101111",
45755 => "1111010110110000",
45756 => "1111010110110000",
45757 => "1111010110110001",
45758 => "1111010110110010",
45759 => "1111010110110010",
45760 => "1111010110110011",
45761 => "1111010110110100",
45762 => "1111010110110100",
45763 => "1111010110110101",
45764 => "1111010110110101",
45765 => "1111010110110110",
45766 => "1111010110110111",
45767 => "1111010110110111",
45768 => "1111010110111000",
45769 => "1111010110111000",
45770 => "1111010110111001",
45771 => "1111010110111010",
45772 => "1111010110111010",
45773 => "1111010110111011",
45774 => "1111010110111100",
45775 => "1111010110111100",
45776 => "1111010110111101",
45777 => "1111010110111101",
45778 => "1111010110111110",
45779 => "1111010110111111",
45780 => "1111010110111111",
45781 => "1111010111000000",
45782 => "1111010111000000",
45783 => "1111010111000001",
45784 => "1111010111000010",
45785 => "1111010111000010",
45786 => "1111010111000011",
45787 => "1111010111000100",
45788 => "1111010111000100",
45789 => "1111010111000101",
45790 => "1111010111000101",
45791 => "1111010111000110",
45792 => "1111010111000111",
45793 => "1111010111000111",
45794 => "1111010111001000",
45795 => "1111010111001000",
45796 => "1111010111001001",
45797 => "1111010111001010",
45798 => "1111010111001010",
45799 => "1111010111001011",
45800 => "1111010111001011",
45801 => "1111010111001100",
45802 => "1111010111001101",
45803 => "1111010111001101",
45804 => "1111010111001110",
45805 => "1111010111001111",
45806 => "1111010111001111",
45807 => "1111010111010000",
45808 => "1111010111010000",
45809 => "1111010111010001",
45810 => "1111010111010010",
45811 => "1111010111010010",
45812 => "1111010111010011",
45813 => "1111010111010011",
45814 => "1111010111010100",
45815 => "1111010111010101",
45816 => "1111010111010101",
45817 => "1111010111010110",
45818 => "1111010111010110",
45819 => "1111010111010111",
45820 => "1111010111011000",
45821 => "1111010111011000",
45822 => "1111010111011001",
45823 => "1111010111011010",
45824 => "1111010111011010",
45825 => "1111010111011011",
45826 => "1111010111011011",
45827 => "1111010111011100",
45828 => "1111010111011101",
45829 => "1111010111011101",
45830 => "1111010111011110",
45831 => "1111010111011110",
45832 => "1111010111011111",
45833 => "1111010111100000",
45834 => "1111010111100000",
45835 => "1111010111100001",
45836 => "1111010111100001",
45837 => "1111010111100010",
45838 => "1111010111100011",
45839 => "1111010111100011",
45840 => "1111010111100100",
45841 => "1111010111100100",
45842 => "1111010111100101",
45843 => "1111010111100110",
45844 => "1111010111100110",
45845 => "1111010111100111",
45846 => "1111010111101000",
45847 => "1111010111101000",
45848 => "1111010111101001",
45849 => "1111010111101001",
45850 => "1111010111101010",
45851 => "1111010111101011",
45852 => "1111010111101011",
45853 => "1111010111101100",
45854 => "1111010111101100",
45855 => "1111010111101101",
45856 => "1111010111101110",
45857 => "1111010111101110",
45858 => "1111010111101111",
45859 => "1111010111101111",
45860 => "1111010111110000",
45861 => "1111010111110001",
45862 => "1111010111110001",
45863 => "1111010111110010",
45864 => "1111010111110010",
45865 => "1111010111110011",
45866 => "1111010111110100",
45867 => "1111010111110100",
45868 => "1111010111110101",
45869 => "1111010111110101",
45870 => "1111010111110110",
45871 => "1111010111110111",
45872 => "1111010111110111",
45873 => "1111010111111000",
45874 => "1111010111111000",
45875 => "1111010111111001",
45876 => "1111010111111010",
45877 => "1111010111111010",
45878 => "1111010111111011",
45879 => "1111010111111011",
45880 => "1111010111111100",
45881 => "1111010111111101",
45882 => "1111010111111101",
45883 => "1111010111111110",
45884 => "1111010111111110",
45885 => "1111010111111111",
45886 => "1111011000000000",
45887 => "1111011000000000",
45888 => "1111011000000001",
45889 => "1111011000000001",
45890 => "1111011000000010",
45891 => "1111011000000011",
45892 => "1111011000000011",
45893 => "1111011000000100",
45894 => "1111011000000100",
45895 => "1111011000000101",
45896 => "1111011000000110",
45897 => "1111011000000110",
45898 => "1111011000000111",
45899 => "1111011000000111",
45900 => "1111011000001000",
45901 => "1111011000001001",
45902 => "1111011000001001",
45903 => "1111011000001010",
45904 => "1111011000001010",
45905 => "1111011000001011",
45906 => "1111011000001100",
45907 => "1111011000001100",
45908 => "1111011000001101",
45909 => "1111011000001101",
45910 => "1111011000001110",
45911 => "1111011000001111",
45912 => "1111011000001111",
45913 => "1111011000010000",
45914 => "1111011000010000",
45915 => "1111011000010001",
45916 => "1111011000010010",
45917 => "1111011000010010",
45918 => "1111011000010011",
45919 => "1111011000010011",
45920 => "1111011000010100",
45921 => "1111011000010101",
45922 => "1111011000010101",
45923 => "1111011000010110",
45924 => "1111011000010110",
45925 => "1111011000010111",
45926 => "1111011000011000",
45927 => "1111011000011000",
45928 => "1111011000011001",
45929 => "1111011000011001",
45930 => "1111011000011010",
45931 => "1111011000011011",
45932 => "1111011000011011",
45933 => "1111011000011100",
45934 => "1111011000011100",
45935 => "1111011000011101",
45936 => "1111011000011110",
45937 => "1111011000011110",
45938 => "1111011000011111",
45939 => "1111011000011111",
45940 => "1111011000100000",
45941 => "1111011000100000",
45942 => "1111011000100001",
45943 => "1111011000100010",
45944 => "1111011000100010",
45945 => "1111011000100011",
45946 => "1111011000100011",
45947 => "1111011000100100",
45948 => "1111011000100101",
45949 => "1111011000100101",
45950 => "1111011000100110",
45951 => "1111011000100110",
45952 => "1111011000100111",
45953 => "1111011000101000",
45954 => "1111011000101000",
45955 => "1111011000101001",
45956 => "1111011000101001",
45957 => "1111011000101010",
45958 => "1111011000101011",
45959 => "1111011000101011",
45960 => "1111011000101100",
45961 => "1111011000101100",
45962 => "1111011000101101",
45963 => "1111011000101101",
45964 => "1111011000101110",
45965 => "1111011000101111",
45966 => "1111011000101111",
45967 => "1111011000110000",
45968 => "1111011000110000",
45969 => "1111011000110001",
45970 => "1111011000110010",
45971 => "1111011000110010",
45972 => "1111011000110011",
45973 => "1111011000110011",
45974 => "1111011000110100",
45975 => "1111011000110101",
45976 => "1111011000110101",
45977 => "1111011000110110",
45978 => "1111011000110110",
45979 => "1111011000110111",
45980 => "1111011000111000",
45981 => "1111011000111000",
45982 => "1111011000111001",
45983 => "1111011000111001",
45984 => "1111011000111010",
45985 => "1111011000111010",
45986 => "1111011000111011",
45987 => "1111011000111100",
45988 => "1111011000111100",
45989 => "1111011000111101",
45990 => "1111011000111101",
45991 => "1111011000111110",
45992 => "1111011000111111",
45993 => "1111011000111111",
45994 => "1111011001000000",
45995 => "1111011001000000",
45996 => "1111011001000001",
45997 => "1111011001000001",
45998 => "1111011001000010",
45999 => "1111011001000011",
46000 => "1111011001000011",
46001 => "1111011001000100",
46002 => "1111011001000100",
46003 => "1111011001000101",
46004 => "1111011001000110",
46005 => "1111011001000110",
46006 => "1111011001000111",
46007 => "1111011001000111",
46008 => "1111011001001000",
46009 => "1111011001001001",
46010 => "1111011001001001",
46011 => "1111011001001010",
46012 => "1111011001001010",
46013 => "1111011001001011",
46014 => "1111011001001011",
46015 => "1111011001001100",
46016 => "1111011001001101",
46017 => "1111011001001101",
46018 => "1111011001001110",
46019 => "1111011001001110",
46020 => "1111011001001111",
46021 => "1111011001010000",
46022 => "1111011001010000",
46023 => "1111011001010001",
46024 => "1111011001010001",
46025 => "1111011001010010",
46026 => "1111011001010010",
46027 => "1111011001010011",
46028 => "1111011001010100",
46029 => "1111011001010100",
46030 => "1111011001010101",
46031 => "1111011001010101",
46032 => "1111011001010110",
46033 => "1111011001010110",
46034 => "1111011001010111",
46035 => "1111011001011000",
46036 => "1111011001011000",
46037 => "1111011001011001",
46038 => "1111011001011001",
46039 => "1111011001011010",
46040 => "1111011001011011",
46041 => "1111011001011011",
46042 => "1111011001011100",
46043 => "1111011001011100",
46044 => "1111011001011101",
46045 => "1111011001011101",
46046 => "1111011001011110",
46047 => "1111011001011111",
46048 => "1111011001011111",
46049 => "1111011001100000",
46050 => "1111011001100000",
46051 => "1111011001100001",
46052 => "1111011001100010",
46053 => "1111011001100010",
46054 => "1111011001100011",
46055 => "1111011001100011",
46056 => "1111011001100100",
46057 => "1111011001100100",
46058 => "1111011001100101",
46059 => "1111011001100110",
46060 => "1111011001100110",
46061 => "1111011001100111",
46062 => "1111011001100111",
46063 => "1111011001101000",
46064 => "1111011001101000",
46065 => "1111011001101001",
46066 => "1111011001101010",
46067 => "1111011001101010",
46068 => "1111011001101011",
46069 => "1111011001101011",
46070 => "1111011001101100",
46071 => "1111011001101100",
46072 => "1111011001101101",
46073 => "1111011001101110",
46074 => "1111011001101110",
46075 => "1111011001101111",
46076 => "1111011001101111",
46077 => "1111011001110000",
46078 => "1111011001110000",
46079 => "1111011001110001",
46080 => "1111011001110010",
46081 => "1111011001110010",
46082 => "1111011001110011",
46083 => "1111011001110011",
46084 => "1111011001110100",
46085 => "1111011001110101",
46086 => "1111011001110101",
46087 => "1111011001110110",
46088 => "1111011001110110",
46089 => "1111011001110111",
46090 => "1111011001110111",
46091 => "1111011001111000",
46092 => "1111011001111001",
46093 => "1111011001111001",
46094 => "1111011001111010",
46095 => "1111011001111010",
46096 => "1111011001111011",
46097 => "1111011001111011",
46098 => "1111011001111100",
46099 => "1111011001111101",
46100 => "1111011001111101",
46101 => "1111011001111110",
46102 => "1111011001111110",
46103 => "1111011001111111",
46104 => "1111011001111111",
46105 => "1111011010000000",
46106 => "1111011010000001",
46107 => "1111011010000001",
46108 => "1111011010000010",
46109 => "1111011010000010",
46110 => "1111011010000011",
46111 => "1111011010000011",
46112 => "1111011010000100",
46113 => "1111011010000101",
46114 => "1111011010000101",
46115 => "1111011010000110",
46116 => "1111011010000110",
46117 => "1111011010000111",
46118 => "1111011010000111",
46119 => "1111011010001000",
46120 => "1111011010001001",
46121 => "1111011010001001",
46122 => "1111011010001010",
46123 => "1111011010001010",
46124 => "1111011010001011",
46125 => "1111011010001011",
46126 => "1111011010001100",
46127 => "1111011010001101",
46128 => "1111011010001101",
46129 => "1111011010001110",
46130 => "1111011010001110",
46131 => "1111011010001111",
46132 => "1111011010001111",
46133 => "1111011010010000",
46134 => "1111011010010001",
46135 => "1111011010010001",
46136 => "1111011010010010",
46137 => "1111011010010010",
46138 => "1111011010010011",
46139 => "1111011010010011",
46140 => "1111011010010100",
46141 => "1111011010010100",
46142 => "1111011010010101",
46143 => "1111011010010110",
46144 => "1111011010010110",
46145 => "1111011010010111",
46146 => "1111011010010111",
46147 => "1111011010011000",
46148 => "1111011010011000",
46149 => "1111011010011001",
46150 => "1111011010011010",
46151 => "1111011010011010",
46152 => "1111011010011011",
46153 => "1111011010011011",
46154 => "1111011010011100",
46155 => "1111011010011100",
46156 => "1111011010011101",
46157 => "1111011010011110",
46158 => "1111011010011110",
46159 => "1111011010011111",
46160 => "1111011010011111",
46161 => "1111011010100000",
46162 => "1111011010100000",
46163 => "1111011010100001",
46164 => "1111011010100001",
46165 => "1111011010100010",
46166 => "1111011010100011",
46167 => "1111011010100011",
46168 => "1111011010100100",
46169 => "1111011010100100",
46170 => "1111011010100101",
46171 => "1111011010100101",
46172 => "1111011010100110",
46173 => "1111011010100111",
46174 => "1111011010100111",
46175 => "1111011010101000",
46176 => "1111011010101000",
46177 => "1111011010101001",
46178 => "1111011010101001",
46179 => "1111011010101010",
46180 => "1111011010101010",
46181 => "1111011010101011",
46182 => "1111011010101100",
46183 => "1111011010101100",
46184 => "1111011010101101",
46185 => "1111011010101101",
46186 => "1111011010101110",
46187 => "1111011010101110",
46188 => "1111011010101111",
46189 => "1111011010110000",
46190 => "1111011010110000",
46191 => "1111011010110001",
46192 => "1111011010110001",
46193 => "1111011010110010",
46194 => "1111011010110010",
46195 => "1111011010110011",
46196 => "1111011010110011",
46197 => "1111011010110100",
46198 => "1111011010110101",
46199 => "1111011010110101",
46200 => "1111011010110110",
46201 => "1111011010110110",
46202 => "1111011010110111",
46203 => "1111011010110111",
46204 => "1111011010111000",
46205 => "1111011010111001",
46206 => "1111011010111001",
46207 => "1111011010111010",
46208 => "1111011010111010",
46209 => "1111011010111011",
46210 => "1111011010111011",
46211 => "1111011010111100",
46212 => "1111011010111100",
46213 => "1111011010111101",
46214 => "1111011010111110",
46215 => "1111011010111110",
46216 => "1111011010111111",
46217 => "1111011010111111",
46218 => "1111011011000000",
46219 => "1111011011000000",
46220 => "1111011011000001",
46221 => "1111011011000001",
46222 => "1111011011000010",
46223 => "1111011011000011",
46224 => "1111011011000011",
46225 => "1111011011000100",
46226 => "1111011011000100",
46227 => "1111011011000101",
46228 => "1111011011000101",
46229 => "1111011011000110",
46230 => "1111011011000110",
46231 => "1111011011000111",
46232 => "1111011011001000",
46233 => "1111011011001000",
46234 => "1111011011001001",
46235 => "1111011011001001",
46236 => "1111011011001010",
46237 => "1111011011001010",
46238 => "1111011011001011",
46239 => "1111011011001011",
46240 => "1111011011001100",
46241 => "1111011011001101",
46242 => "1111011011001101",
46243 => "1111011011001110",
46244 => "1111011011001110",
46245 => "1111011011001111",
46246 => "1111011011001111",
46247 => "1111011011010000",
46248 => "1111011011010000",
46249 => "1111011011010001",
46250 => "1111011011010010",
46251 => "1111011011010010",
46252 => "1111011011010011",
46253 => "1111011011010011",
46254 => "1111011011010100",
46255 => "1111011011010100",
46256 => "1111011011010101",
46257 => "1111011011010101",
46258 => "1111011011010110",
46259 => "1111011011010110",
46260 => "1111011011010111",
46261 => "1111011011011000",
46262 => "1111011011011000",
46263 => "1111011011011001",
46264 => "1111011011011001",
46265 => "1111011011011010",
46266 => "1111011011011010",
46267 => "1111011011011011",
46268 => "1111011011011011",
46269 => "1111011011011100",
46270 => "1111011011011101",
46271 => "1111011011011101",
46272 => "1111011011011110",
46273 => "1111011011011110",
46274 => "1111011011011111",
46275 => "1111011011011111",
46276 => "1111011011100000",
46277 => "1111011011100000",
46278 => "1111011011100001",
46279 => "1111011011100010",
46280 => "1111011011100010",
46281 => "1111011011100011",
46282 => "1111011011100011",
46283 => "1111011011100100",
46284 => "1111011011100100",
46285 => "1111011011100101",
46286 => "1111011011100101",
46287 => "1111011011100110",
46288 => "1111011011100110",
46289 => "1111011011100111",
46290 => "1111011011101000",
46291 => "1111011011101000",
46292 => "1111011011101001",
46293 => "1111011011101001",
46294 => "1111011011101010",
46295 => "1111011011101010",
46296 => "1111011011101011",
46297 => "1111011011101011",
46298 => "1111011011101100",
46299 => "1111011011101100",
46300 => "1111011011101101",
46301 => "1111011011101110",
46302 => "1111011011101110",
46303 => "1111011011101111",
46304 => "1111011011101111",
46305 => "1111011011110000",
46306 => "1111011011110000",
46307 => "1111011011110001",
46308 => "1111011011110001",
46309 => "1111011011110010",
46310 => "1111011011110010",
46311 => "1111011011110011",
46312 => "1111011011110100",
46313 => "1111011011110100",
46314 => "1111011011110101",
46315 => "1111011011110101",
46316 => "1111011011110110",
46317 => "1111011011110110",
46318 => "1111011011110111",
46319 => "1111011011110111",
46320 => "1111011011111000",
46321 => "1111011011111000",
46322 => "1111011011111001",
46323 => "1111011011111010",
46324 => "1111011011111010",
46325 => "1111011011111011",
46326 => "1111011011111011",
46327 => "1111011011111100",
46328 => "1111011011111100",
46329 => "1111011011111101",
46330 => "1111011011111101",
46331 => "1111011011111110",
46332 => "1111011011111110",
46333 => "1111011011111111",
46334 => "1111011100000000",
46335 => "1111011100000000",
46336 => "1111011100000001",
46337 => "1111011100000001",
46338 => "1111011100000010",
46339 => "1111011100000010",
46340 => "1111011100000011",
46341 => "1111011100000011",
46342 => "1111011100000100",
46343 => "1111011100000100",
46344 => "1111011100000101",
46345 => "1111011100000110",
46346 => "1111011100000110",
46347 => "1111011100000111",
46348 => "1111011100000111",
46349 => "1111011100001000",
46350 => "1111011100001000",
46351 => "1111011100001001",
46352 => "1111011100001001",
46353 => "1111011100001010",
46354 => "1111011100001010",
46355 => "1111011100001011",
46356 => "1111011100001011",
46357 => "1111011100001100",
46358 => "1111011100001101",
46359 => "1111011100001101",
46360 => "1111011100001110",
46361 => "1111011100001110",
46362 => "1111011100001111",
46363 => "1111011100001111",
46364 => "1111011100010000",
46365 => "1111011100010000",
46366 => "1111011100010001",
46367 => "1111011100010001",
46368 => "1111011100010010",
46369 => "1111011100010010",
46370 => "1111011100010011",
46371 => "1111011100010100",
46372 => "1111011100010100",
46373 => "1111011100010101",
46374 => "1111011100010101",
46375 => "1111011100010110",
46376 => "1111011100010110",
46377 => "1111011100010111",
46378 => "1111011100010111",
46379 => "1111011100011000",
46380 => "1111011100011000",
46381 => "1111011100011001",
46382 => "1111011100011001",
46383 => "1111011100011010",
46384 => "1111011100011011",
46385 => "1111011100011011",
46386 => "1111011100011100",
46387 => "1111011100011100",
46388 => "1111011100011101",
46389 => "1111011100011101",
46390 => "1111011100011110",
46391 => "1111011100011110",
46392 => "1111011100011111",
46393 => "1111011100011111",
46394 => "1111011100100000",
46395 => "1111011100100000",
46396 => "1111011100100001",
46397 => "1111011100100001",
46398 => "1111011100100010",
46399 => "1111011100100011",
46400 => "1111011100100011",
46401 => "1111011100100100",
46402 => "1111011100100100",
46403 => "1111011100100101",
46404 => "1111011100100101",
46405 => "1111011100100110",
46406 => "1111011100100110",
46407 => "1111011100100111",
46408 => "1111011100100111",
46409 => "1111011100101000",
46410 => "1111011100101000",
46411 => "1111011100101001",
46412 => "1111011100101010",
46413 => "1111011100101010",
46414 => "1111011100101011",
46415 => "1111011100101011",
46416 => "1111011100101100",
46417 => "1111011100101100",
46418 => "1111011100101101",
46419 => "1111011100101101",
46420 => "1111011100101110",
46421 => "1111011100101110",
46422 => "1111011100101111",
46423 => "1111011100101111",
46424 => "1111011100110000",
46425 => "1111011100110000",
46426 => "1111011100110001",
46427 => "1111011100110001",
46428 => "1111011100110010",
46429 => "1111011100110011",
46430 => "1111011100110011",
46431 => "1111011100110100",
46432 => "1111011100110100",
46433 => "1111011100110101",
46434 => "1111011100110101",
46435 => "1111011100110110",
46436 => "1111011100110110",
46437 => "1111011100110111",
46438 => "1111011100110111",
46439 => "1111011100111000",
46440 => "1111011100111000",
46441 => "1111011100111001",
46442 => "1111011100111001",
46443 => "1111011100111010",
46444 => "1111011100111011",
46445 => "1111011100111011",
46446 => "1111011100111100",
46447 => "1111011100111100",
46448 => "1111011100111101",
46449 => "1111011100111101",
46450 => "1111011100111110",
46451 => "1111011100111110",
46452 => "1111011100111111",
46453 => "1111011100111111",
46454 => "1111011101000000",
46455 => "1111011101000000",
46456 => "1111011101000001",
46457 => "1111011101000001",
46458 => "1111011101000010",
46459 => "1111011101000010",
46460 => "1111011101000011",
46461 => "1111011101000011",
46462 => "1111011101000100",
46463 => "1111011101000101",
46464 => "1111011101000101",
46465 => "1111011101000110",
46466 => "1111011101000110",
46467 => "1111011101000111",
46468 => "1111011101000111",
46469 => "1111011101001000",
46470 => "1111011101001000",
46471 => "1111011101001001",
46472 => "1111011101001001",
46473 => "1111011101001010",
46474 => "1111011101001010",
46475 => "1111011101001011",
46476 => "1111011101001011",
46477 => "1111011101001100",
46478 => "1111011101001100",
46479 => "1111011101001101",
46480 => "1111011101001101",
46481 => "1111011101001110",
46482 => "1111011101001111",
46483 => "1111011101001111",
46484 => "1111011101010000",
46485 => "1111011101010000",
46486 => "1111011101010001",
46487 => "1111011101010001",
46488 => "1111011101010010",
46489 => "1111011101010010",
46490 => "1111011101010011",
46491 => "1111011101010011",
46492 => "1111011101010100",
46493 => "1111011101010100",
46494 => "1111011101010101",
46495 => "1111011101010101",
46496 => "1111011101010110",
46497 => "1111011101010110",
46498 => "1111011101010111",
46499 => "1111011101010111",
46500 => "1111011101011000",
46501 => "1111011101011000",
46502 => "1111011101011001",
46503 => "1111011101011010",
46504 => "1111011101011010",
46505 => "1111011101011011",
46506 => "1111011101011011",
46507 => "1111011101011100",
46508 => "1111011101011100",
46509 => "1111011101011101",
46510 => "1111011101011101",
46511 => "1111011101011110",
46512 => "1111011101011110",
46513 => "1111011101011111",
46514 => "1111011101011111",
46515 => "1111011101100000",
46516 => "1111011101100000",
46517 => "1111011101100001",
46518 => "1111011101100001",
46519 => "1111011101100010",
46520 => "1111011101100010",
46521 => "1111011101100011",
46522 => "1111011101100011",
46523 => "1111011101100100",
46524 => "1111011101100100",
46525 => "1111011101100101",
46526 => "1111011101100110",
46527 => "1111011101100110",
46528 => "1111011101100111",
46529 => "1111011101100111",
46530 => "1111011101101000",
46531 => "1111011101101000",
46532 => "1111011101101001",
46533 => "1111011101101001",
46534 => "1111011101101010",
46535 => "1111011101101010",
46536 => "1111011101101011",
46537 => "1111011101101011",
46538 => "1111011101101100",
46539 => "1111011101101100",
46540 => "1111011101101101",
46541 => "1111011101101101",
46542 => "1111011101101110",
46543 => "1111011101101110",
46544 => "1111011101101111",
46545 => "1111011101101111",
46546 => "1111011101110000",
46547 => "1111011101110000",
46548 => "1111011101110001",
46549 => "1111011101110001",
46550 => "1111011101110010",
46551 => "1111011101110010",
46552 => "1111011101110011",
46553 => "1111011101110011",
46554 => "1111011101110100",
46555 => "1111011101110101",
46556 => "1111011101110101",
46557 => "1111011101110110",
46558 => "1111011101110110",
46559 => "1111011101110111",
46560 => "1111011101110111",
46561 => "1111011101111000",
46562 => "1111011101111000",
46563 => "1111011101111001",
46564 => "1111011101111001",
46565 => "1111011101111010",
46566 => "1111011101111010",
46567 => "1111011101111011",
46568 => "1111011101111011",
46569 => "1111011101111100",
46570 => "1111011101111100",
46571 => "1111011101111101",
46572 => "1111011101111101",
46573 => "1111011101111110",
46574 => "1111011101111110",
46575 => "1111011101111111",
46576 => "1111011101111111",
46577 => "1111011110000000",
46578 => "1111011110000000",
46579 => "1111011110000001",
46580 => "1111011110000001",
46581 => "1111011110000010",
46582 => "1111011110000010",
46583 => "1111011110000011",
46584 => "1111011110000011",
46585 => "1111011110000100",
46586 => "1111011110000100",
46587 => "1111011110000101",
46588 => "1111011110000101",
46589 => "1111011110000110",
46590 => "1111011110000111",
46591 => "1111011110000111",
46592 => "1111011110001000",
46593 => "1111011110001000",
46594 => "1111011110001001",
46595 => "1111011110001001",
46596 => "1111011110001010",
46597 => "1111011110001010",
46598 => "1111011110001011",
46599 => "1111011110001011",
46600 => "1111011110001100",
46601 => "1111011110001100",
46602 => "1111011110001101",
46603 => "1111011110001101",
46604 => "1111011110001110",
46605 => "1111011110001110",
46606 => "1111011110001111",
46607 => "1111011110001111",
46608 => "1111011110010000",
46609 => "1111011110010000",
46610 => "1111011110010001",
46611 => "1111011110010001",
46612 => "1111011110010010",
46613 => "1111011110010010",
46614 => "1111011110010011",
46615 => "1111011110010011",
46616 => "1111011110010100",
46617 => "1111011110010100",
46618 => "1111011110010101",
46619 => "1111011110010101",
46620 => "1111011110010110",
46621 => "1111011110010110",
46622 => "1111011110010111",
46623 => "1111011110010111",
46624 => "1111011110011000",
46625 => "1111011110011000",
46626 => "1111011110011001",
46627 => "1111011110011001",
46628 => "1111011110011010",
46629 => "1111011110011010",
46630 => "1111011110011011",
46631 => "1111011110011011",
46632 => "1111011110011100",
46633 => "1111011110011100",
46634 => "1111011110011101",
46635 => "1111011110011101",
46636 => "1111011110011110",
46637 => "1111011110011110",
46638 => "1111011110011111",
46639 => "1111011110011111",
46640 => "1111011110100000",
46641 => "1111011110100000",
46642 => "1111011110100001",
46643 => "1111011110100001",
46644 => "1111011110100010",
46645 => "1111011110100011",
46646 => "1111011110100011",
46647 => "1111011110100100",
46648 => "1111011110100100",
46649 => "1111011110100101",
46650 => "1111011110100101",
46651 => "1111011110100110",
46652 => "1111011110100110",
46653 => "1111011110100111",
46654 => "1111011110100111",
46655 => "1111011110101000",
46656 => "1111011110101000",
46657 => "1111011110101001",
46658 => "1111011110101001",
46659 => "1111011110101010",
46660 => "1111011110101010",
46661 => "1111011110101011",
46662 => "1111011110101011",
46663 => "1111011110101100",
46664 => "1111011110101100",
46665 => "1111011110101101",
46666 => "1111011110101101",
46667 => "1111011110101110",
46668 => "1111011110101110",
46669 => "1111011110101111",
46670 => "1111011110101111",
46671 => "1111011110110000",
46672 => "1111011110110000",
46673 => "1111011110110001",
46674 => "1111011110110001",
46675 => "1111011110110010",
46676 => "1111011110110010",
46677 => "1111011110110011",
46678 => "1111011110110011",
46679 => "1111011110110100",
46680 => "1111011110110100",
46681 => "1111011110110101",
46682 => "1111011110110101",
46683 => "1111011110110110",
46684 => "1111011110110110",
46685 => "1111011110110111",
46686 => "1111011110110111",
46687 => "1111011110111000",
46688 => "1111011110111000",
46689 => "1111011110111001",
46690 => "1111011110111001",
46691 => "1111011110111010",
46692 => "1111011110111010",
46693 => "1111011110111011",
46694 => "1111011110111011",
46695 => "1111011110111100",
46696 => "1111011110111100",
46697 => "1111011110111101",
46698 => "1111011110111101",
46699 => "1111011110111110",
46700 => "1111011110111110",
46701 => "1111011110111111",
46702 => "1111011110111111",
46703 => "1111011111000000",
46704 => "1111011111000000",
46705 => "1111011111000001",
46706 => "1111011111000001",
46707 => "1111011111000010",
46708 => "1111011111000010",
46709 => "1111011111000011",
46710 => "1111011111000011",
46711 => "1111011111000100",
46712 => "1111011111000100",
46713 => "1111011111000101",
46714 => "1111011111000101",
46715 => "1111011111000110",
46716 => "1111011111000110",
46717 => "1111011111000111",
46718 => "1111011111000111",
46719 => "1111011111001000",
46720 => "1111011111001000",
46721 => "1111011111001001",
46722 => "1111011111001001",
46723 => "1111011111001010",
46724 => "1111011111001010",
46725 => "1111011111001011",
46726 => "1111011111001011",
46727 => "1111011111001100",
46728 => "1111011111001100",
46729 => "1111011111001101",
46730 => "1111011111001101",
46731 => "1111011111001110",
46732 => "1111011111001110",
46733 => "1111011111001111",
46734 => "1111011111001111",
46735 => "1111011111010000",
46736 => "1111011111010000",
46737 => "1111011111010001",
46738 => "1111011111010001",
46739 => "1111011111010010",
46740 => "1111011111010010",
46741 => "1111011111010011",
46742 => "1111011111010011",
46743 => "1111011111010100",
46744 => "1111011111010100",
46745 => "1111011111010100",
46746 => "1111011111010101",
46747 => "1111011111010101",
46748 => "1111011111010110",
46749 => "1111011111010110",
46750 => "1111011111010111",
46751 => "1111011111010111",
46752 => "1111011111011000",
46753 => "1111011111011000",
46754 => "1111011111011001",
46755 => "1111011111011001",
46756 => "1111011111011010",
46757 => "1111011111011010",
46758 => "1111011111011011",
46759 => "1111011111011011",
46760 => "1111011111011100",
46761 => "1111011111011100",
46762 => "1111011111011101",
46763 => "1111011111011101",
46764 => "1111011111011110",
46765 => "1111011111011110",
46766 => "1111011111011111",
46767 => "1111011111011111",
46768 => "1111011111100000",
46769 => "1111011111100000",
46770 => "1111011111100001",
46771 => "1111011111100001",
46772 => "1111011111100010",
46773 => "1111011111100010",
46774 => "1111011111100011",
46775 => "1111011111100011",
46776 => "1111011111100100",
46777 => "1111011111100100",
46778 => "1111011111100101",
46779 => "1111011111100101",
46780 => "1111011111100110",
46781 => "1111011111100110",
46782 => "1111011111100111",
46783 => "1111011111100111",
46784 => "1111011111101000",
46785 => "1111011111101000",
46786 => "1111011111101001",
46787 => "1111011111101001",
46788 => "1111011111101010",
46789 => "1111011111101010",
46790 => "1111011111101011",
46791 => "1111011111101011",
46792 => "1111011111101100",
46793 => "1111011111101100",
46794 => "1111011111101101",
46795 => "1111011111101101",
46796 => "1111011111101110",
46797 => "1111011111101110",
46798 => "1111011111101111",
46799 => "1111011111101111",
46800 => "1111011111110000",
46801 => "1111011111110000",
46802 => "1111011111110000",
46803 => "1111011111110001",
46804 => "1111011111110001",
46805 => "1111011111110010",
46806 => "1111011111110010",
46807 => "1111011111110011",
46808 => "1111011111110011",
46809 => "1111011111110100",
46810 => "1111011111110100",
46811 => "1111011111110101",
46812 => "1111011111110101",
46813 => "1111011111110110",
46814 => "1111011111110110",
46815 => "1111011111110111",
46816 => "1111011111110111",
46817 => "1111011111111000",
46818 => "1111011111111000",
46819 => "1111011111111001",
46820 => "1111011111111001",
46821 => "1111011111111010",
46822 => "1111011111111010",
46823 => "1111011111111011",
46824 => "1111011111111011",
46825 => "1111011111111100",
46826 => "1111011111111100",
46827 => "1111011111111101",
46828 => "1111011111111101",
46829 => "1111011111111110",
46830 => "1111011111111110",
46831 => "1111011111111111",
46832 => "1111011111111111",
46833 => "1111100000000000",
46834 => "1111100000000000",
46835 => "1111100000000001",
46836 => "1111100000000001",
46837 => "1111100000000001",
46838 => "1111100000000010",
46839 => "1111100000000010",
46840 => "1111100000000011",
46841 => "1111100000000011",
46842 => "1111100000000100",
46843 => "1111100000000100",
46844 => "1111100000000101",
46845 => "1111100000000101",
46846 => "1111100000000110",
46847 => "1111100000000110",
46848 => "1111100000000111",
46849 => "1111100000000111",
46850 => "1111100000001000",
46851 => "1111100000001000",
46852 => "1111100000001001",
46853 => "1111100000001001",
46854 => "1111100000001010",
46855 => "1111100000001010",
46856 => "1111100000001011",
46857 => "1111100000001011",
46858 => "1111100000001100",
46859 => "1111100000001100",
46860 => "1111100000001101",
46861 => "1111100000001101",
46862 => "1111100000001110",
46863 => "1111100000001110",
46864 => "1111100000001111",
46865 => "1111100000001111",
46866 => "1111100000001111",
46867 => "1111100000010000",
46868 => "1111100000010000",
46869 => "1111100000010001",
46870 => "1111100000010001",
46871 => "1111100000010010",
46872 => "1111100000010010",
46873 => "1111100000010011",
46874 => "1111100000010011",
46875 => "1111100000010100",
46876 => "1111100000010100",
46877 => "1111100000010101",
46878 => "1111100000010101",
46879 => "1111100000010110",
46880 => "1111100000010110",
46881 => "1111100000010111",
46882 => "1111100000010111",
46883 => "1111100000011000",
46884 => "1111100000011000",
46885 => "1111100000011001",
46886 => "1111100000011001",
46887 => "1111100000011010",
46888 => "1111100000011010",
46889 => "1111100000011011",
46890 => "1111100000011011",
46891 => "1111100000011011",
46892 => "1111100000011100",
46893 => "1111100000011100",
46894 => "1111100000011101",
46895 => "1111100000011101",
46896 => "1111100000011110",
46897 => "1111100000011110",
46898 => "1111100000011111",
46899 => "1111100000011111",
46900 => "1111100000100000",
46901 => "1111100000100000",
46902 => "1111100000100001",
46903 => "1111100000100001",
46904 => "1111100000100010",
46905 => "1111100000100010",
46906 => "1111100000100011",
46907 => "1111100000100011",
46908 => "1111100000100100",
46909 => "1111100000100100",
46910 => "1111100000100101",
46911 => "1111100000100101",
46912 => "1111100000100101",
46913 => "1111100000100110",
46914 => "1111100000100110",
46915 => "1111100000100111",
46916 => "1111100000100111",
46917 => "1111100000101000",
46918 => "1111100000101000",
46919 => "1111100000101001",
46920 => "1111100000101001",
46921 => "1111100000101010",
46922 => "1111100000101010",
46923 => "1111100000101011",
46924 => "1111100000101011",
46925 => "1111100000101100",
46926 => "1111100000101100",
46927 => "1111100000101101",
46928 => "1111100000101101",
46929 => "1111100000101110",
46930 => "1111100000101110",
46931 => "1111100000101110",
46932 => "1111100000101111",
46933 => "1111100000101111",
46934 => "1111100000110000",
46935 => "1111100000110000",
46936 => "1111100000110001",
46937 => "1111100000110001",
46938 => "1111100000110010",
46939 => "1111100000110010",
46940 => "1111100000110011",
46941 => "1111100000110011",
46942 => "1111100000110100",
46943 => "1111100000110100",
46944 => "1111100000110101",
46945 => "1111100000110101",
46946 => "1111100000110110",
46947 => "1111100000110110",
46948 => "1111100000110111",
46949 => "1111100000110111",
46950 => "1111100000110111",
46951 => "1111100000111000",
46952 => "1111100000111000",
46953 => "1111100000111001",
46954 => "1111100000111001",
46955 => "1111100000111010",
46956 => "1111100000111010",
46957 => "1111100000111011",
46958 => "1111100000111011",
46959 => "1111100000111100",
46960 => "1111100000111100",
46961 => "1111100000111101",
46962 => "1111100000111101",
46963 => "1111100000111110",
46964 => "1111100000111110",
46965 => "1111100000111111",
46966 => "1111100000111111",
46967 => "1111100000111111",
46968 => "1111100001000000",
46969 => "1111100001000000",
46970 => "1111100001000001",
46971 => "1111100001000001",
46972 => "1111100001000010",
46973 => "1111100001000010",
46974 => "1111100001000011",
46975 => "1111100001000011",
46976 => "1111100001000100",
46977 => "1111100001000100",
46978 => "1111100001000101",
46979 => "1111100001000101",
46980 => "1111100001000110",
46981 => "1111100001000110",
46982 => "1111100001000111",
46983 => "1111100001000111",
46984 => "1111100001000111",
46985 => "1111100001001000",
46986 => "1111100001001000",
46987 => "1111100001001001",
46988 => "1111100001001001",
46989 => "1111100001001010",
46990 => "1111100001001010",
46991 => "1111100001001011",
46992 => "1111100001001011",
46993 => "1111100001001100",
46994 => "1111100001001100",
46995 => "1111100001001101",
46996 => "1111100001001101",
46997 => "1111100001001110",
46998 => "1111100001001110",
46999 => "1111100001001110",
47000 => "1111100001001111",
47001 => "1111100001001111",
47002 => "1111100001010000",
47003 => "1111100001010000",
47004 => "1111100001010001",
47005 => "1111100001010001",
47006 => "1111100001010010",
47007 => "1111100001010010",
47008 => "1111100001010011",
47009 => "1111100001010011",
47010 => "1111100001010100",
47011 => "1111100001010100",
47012 => "1111100001010100",
47013 => "1111100001010101",
47014 => "1111100001010101",
47015 => "1111100001010110",
47016 => "1111100001010110",
47017 => "1111100001010111",
47018 => "1111100001010111",
47019 => "1111100001011000",
47020 => "1111100001011000",
47021 => "1111100001011001",
47022 => "1111100001011001",
47023 => "1111100001011010",
47024 => "1111100001011010",
47025 => "1111100001011011",
47026 => "1111100001011011",
47027 => "1111100001011011",
47028 => "1111100001011100",
47029 => "1111100001011100",
47030 => "1111100001011101",
47031 => "1111100001011101",
47032 => "1111100001011110",
47033 => "1111100001011110",
47034 => "1111100001011111",
47035 => "1111100001011111",
47036 => "1111100001100000",
47037 => "1111100001100000",
47038 => "1111100001100001",
47039 => "1111100001100001",
47040 => "1111100001100001",
47041 => "1111100001100010",
47042 => "1111100001100010",
47043 => "1111100001100011",
47044 => "1111100001100011",
47045 => "1111100001100100",
47046 => "1111100001100100",
47047 => "1111100001100101",
47048 => "1111100001100101",
47049 => "1111100001100110",
47050 => "1111100001100110",
47051 => "1111100001100111",
47052 => "1111100001100111",
47053 => "1111100001100111",
47054 => "1111100001101000",
47055 => "1111100001101000",
47056 => "1111100001101001",
47057 => "1111100001101001",
47058 => "1111100001101010",
47059 => "1111100001101010",
47060 => "1111100001101011",
47061 => "1111100001101011",
47062 => "1111100001101100",
47063 => "1111100001101100",
47064 => "1111100001101101",
47065 => "1111100001101101",
47066 => "1111100001101101",
47067 => "1111100001101110",
47068 => "1111100001101110",
47069 => "1111100001101111",
47070 => "1111100001101111",
47071 => "1111100001110000",
47072 => "1111100001110000",
47073 => "1111100001110001",
47074 => "1111100001110001",
47075 => "1111100001110010",
47076 => "1111100001110010",
47077 => "1111100001110010",
47078 => "1111100001110011",
47079 => "1111100001110011",
47080 => "1111100001110100",
47081 => "1111100001110100",
47082 => "1111100001110101",
47083 => "1111100001110101",
47084 => "1111100001110110",
47085 => "1111100001110110",
47086 => "1111100001110111",
47087 => "1111100001110111",
47088 => "1111100001111000",
47089 => "1111100001111000",
47090 => "1111100001111000",
47091 => "1111100001111001",
47092 => "1111100001111001",
47093 => "1111100001111010",
47094 => "1111100001111010",
47095 => "1111100001111011",
47096 => "1111100001111011",
47097 => "1111100001111100",
47098 => "1111100001111100",
47099 => "1111100001111101",
47100 => "1111100001111101",
47101 => "1111100001111101",
47102 => "1111100001111110",
47103 => "1111100001111110",
47104 => "1111100001111111",
47105 => "1111100001111111",
47106 => "1111100010000000",
47107 => "1111100010000000",
47108 => "1111100010000001",
47109 => "1111100010000001",
47110 => "1111100010000010",
47111 => "1111100010000010",
47112 => "1111100010000010",
47113 => "1111100010000011",
47114 => "1111100010000011",
47115 => "1111100010000100",
47116 => "1111100010000100",
47117 => "1111100010000101",
47118 => "1111100010000101",
47119 => "1111100010000110",
47120 => "1111100010000110",
47121 => "1111100010000111",
47122 => "1111100010000111",
47123 => "1111100010000111",
47124 => "1111100010001000",
47125 => "1111100010001000",
47126 => "1111100010001001",
47127 => "1111100010001001",
47128 => "1111100010001010",
47129 => "1111100010001010",
47130 => "1111100010001011",
47131 => "1111100010001011",
47132 => "1111100010001100",
47133 => "1111100010001100",
47134 => "1111100010001100",
47135 => "1111100010001101",
47136 => "1111100010001101",
47137 => "1111100010001110",
47138 => "1111100010001110",
47139 => "1111100010001111",
47140 => "1111100010001111",
47141 => "1111100010010000",
47142 => "1111100010010000",
47143 => "1111100010010000",
47144 => "1111100010010001",
47145 => "1111100010010001",
47146 => "1111100010010010",
47147 => "1111100010010010",
47148 => "1111100010010011",
47149 => "1111100010010011",
47150 => "1111100010010100",
47151 => "1111100010010100",
47152 => "1111100010010101",
47153 => "1111100010010101",
47154 => "1111100010010101",
47155 => "1111100010010110",
47156 => "1111100010010110",
47157 => "1111100010010111",
47158 => "1111100010010111",
47159 => "1111100010011000",
47160 => "1111100010011000",
47161 => "1111100010011001",
47162 => "1111100010011001",
47163 => "1111100010011001",
47164 => "1111100010011010",
47165 => "1111100010011010",
47166 => "1111100010011011",
47167 => "1111100010011011",
47168 => "1111100010011100",
47169 => "1111100010011100",
47170 => "1111100010011101",
47171 => "1111100010011101",
47172 => "1111100010011110",
47173 => "1111100010011110",
47174 => "1111100010011110",
47175 => "1111100010011111",
47176 => "1111100010011111",
47177 => "1111100010100000",
47178 => "1111100010100000",
47179 => "1111100010100001",
47180 => "1111100010100001",
47181 => "1111100010100010",
47182 => "1111100010100010",
47183 => "1111100010100010",
47184 => "1111100010100011",
47185 => "1111100010100011",
47186 => "1111100010100100",
47187 => "1111100010100100",
47188 => "1111100010100101",
47189 => "1111100010100101",
47190 => "1111100010100110",
47191 => "1111100010100110",
47192 => "1111100010100110",
47193 => "1111100010100111",
47194 => "1111100010100111",
47195 => "1111100010101000",
47196 => "1111100010101000",
47197 => "1111100010101001",
47198 => "1111100010101001",
47199 => "1111100010101010",
47200 => "1111100010101010",
47201 => "1111100010101010",
47202 => "1111100010101011",
47203 => "1111100010101011",
47204 => "1111100010101100",
47205 => "1111100010101100",
47206 => "1111100010101101",
47207 => "1111100010101101",
47208 => "1111100010101110",
47209 => "1111100010101110",
47210 => "1111100010101110",
47211 => "1111100010101111",
47212 => "1111100010101111",
47213 => "1111100010110000",
47214 => "1111100010110000",
47215 => "1111100010110001",
47216 => "1111100010110001",
47217 => "1111100010110010",
47218 => "1111100010110010",
47219 => "1111100010110010",
47220 => "1111100010110011",
47221 => "1111100010110011",
47222 => "1111100010110100",
47223 => "1111100010110100",
47224 => "1111100010110101",
47225 => "1111100010110101",
47226 => "1111100010110110",
47227 => "1111100010110110",
47228 => "1111100010110110",
47229 => "1111100010110111",
47230 => "1111100010110111",
47231 => "1111100010111000",
47232 => "1111100010111000",
47233 => "1111100010111001",
47234 => "1111100010111001",
47235 => "1111100010111010",
47236 => "1111100010111010",
47237 => "1111100010111010",
47238 => "1111100010111011",
47239 => "1111100010111011",
47240 => "1111100010111100",
47241 => "1111100010111100",
47242 => "1111100010111101",
47243 => "1111100010111101",
47244 => "1111100010111110",
47245 => "1111100010111110",
47246 => "1111100010111110",
47247 => "1111100010111111",
47248 => "1111100010111111",
47249 => "1111100011000000",
47250 => "1111100011000000",
47251 => "1111100011000001",
47252 => "1111100011000001",
47253 => "1111100011000001",
47254 => "1111100011000010",
47255 => "1111100011000010",
47256 => "1111100011000011",
47257 => "1111100011000011",
47258 => "1111100011000100",
47259 => "1111100011000100",
47260 => "1111100011000101",
47261 => "1111100011000101",
47262 => "1111100011000101",
47263 => "1111100011000110",
47264 => "1111100011000110",
47265 => "1111100011000111",
47266 => "1111100011000111",
47267 => "1111100011001000",
47268 => "1111100011001000",
47269 => "1111100011001001",
47270 => "1111100011001001",
47271 => "1111100011001001",
47272 => "1111100011001010",
47273 => "1111100011001010",
47274 => "1111100011001011",
47275 => "1111100011001011",
47276 => "1111100011001100",
47277 => "1111100011001100",
47278 => "1111100011001100",
47279 => "1111100011001101",
47280 => "1111100011001101",
47281 => "1111100011001110",
47282 => "1111100011001110",
47283 => "1111100011001111",
47284 => "1111100011001111",
47285 => "1111100011010000",
47286 => "1111100011010000",
47287 => "1111100011010000",
47288 => "1111100011010001",
47289 => "1111100011010001",
47290 => "1111100011010010",
47291 => "1111100011010010",
47292 => "1111100011010011",
47293 => "1111100011010011",
47294 => "1111100011010011",
47295 => "1111100011010100",
47296 => "1111100011010100",
47297 => "1111100011010101",
47298 => "1111100011010101",
47299 => "1111100011010110",
47300 => "1111100011010110",
47301 => "1111100011010110",
47302 => "1111100011010111",
47303 => "1111100011010111",
47304 => "1111100011011000",
47305 => "1111100011011000",
47306 => "1111100011011001",
47307 => "1111100011011001",
47308 => "1111100011011010",
47309 => "1111100011011010",
47310 => "1111100011011010",
47311 => "1111100011011011",
47312 => "1111100011011011",
47313 => "1111100011011100",
47314 => "1111100011011100",
47315 => "1111100011011101",
47316 => "1111100011011101",
47317 => "1111100011011101",
47318 => "1111100011011110",
47319 => "1111100011011110",
47320 => "1111100011011111",
47321 => "1111100011011111",
47322 => "1111100011100000",
47323 => "1111100011100000",
47324 => "1111100011100000",
47325 => "1111100011100001",
47326 => "1111100011100001",
47327 => "1111100011100010",
47328 => "1111100011100010",
47329 => "1111100011100011",
47330 => "1111100011100011",
47331 => "1111100011100011",
47332 => "1111100011100100",
47333 => "1111100011100100",
47334 => "1111100011100101",
47335 => "1111100011100101",
47336 => "1111100011100110",
47337 => "1111100011100110",
47338 => "1111100011100111",
47339 => "1111100011100111",
47340 => "1111100011100111",
47341 => "1111100011101000",
47342 => "1111100011101000",
47343 => "1111100011101001",
47344 => "1111100011101001",
47345 => "1111100011101010",
47346 => "1111100011101010",
47347 => "1111100011101010",
47348 => "1111100011101011",
47349 => "1111100011101011",
47350 => "1111100011101100",
47351 => "1111100011101100",
47352 => "1111100011101101",
47353 => "1111100011101101",
47354 => "1111100011101101",
47355 => "1111100011101110",
47356 => "1111100011101110",
47357 => "1111100011101111",
47358 => "1111100011101111",
47359 => "1111100011110000",
47360 => "1111100011110000",
47361 => "1111100011110000",
47362 => "1111100011110001",
47363 => "1111100011110001",
47364 => "1111100011110010",
47365 => "1111100011110010",
47366 => "1111100011110011",
47367 => "1111100011110011",
47368 => "1111100011110011",
47369 => "1111100011110100",
47370 => "1111100011110100",
47371 => "1111100011110101",
47372 => "1111100011110101",
47373 => "1111100011110110",
47374 => "1111100011110110",
47375 => "1111100011110110",
47376 => "1111100011110111",
47377 => "1111100011110111",
47378 => "1111100011111000",
47379 => "1111100011111000",
47380 => "1111100011111001",
47381 => "1111100011111001",
47382 => "1111100011111001",
47383 => "1111100011111010",
47384 => "1111100011111010",
47385 => "1111100011111011",
47386 => "1111100011111011",
47387 => "1111100011111100",
47388 => "1111100011111100",
47389 => "1111100011111100",
47390 => "1111100011111101",
47391 => "1111100011111101",
47392 => "1111100011111110",
47393 => "1111100011111110",
47394 => "1111100011111111",
47395 => "1111100011111111",
47396 => "1111100011111111",
47397 => "1111100100000000",
47398 => "1111100100000000",
47399 => "1111100100000001",
47400 => "1111100100000001",
47401 => "1111100100000001",
47402 => "1111100100000010",
47403 => "1111100100000010",
47404 => "1111100100000011",
47405 => "1111100100000011",
47406 => "1111100100000100",
47407 => "1111100100000100",
47408 => "1111100100000100",
47409 => "1111100100000101",
47410 => "1111100100000101",
47411 => "1111100100000110",
47412 => "1111100100000110",
47413 => "1111100100000111",
47414 => "1111100100000111",
47415 => "1111100100000111",
47416 => "1111100100001000",
47417 => "1111100100001000",
47418 => "1111100100001001",
47419 => "1111100100001001",
47420 => "1111100100001010",
47421 => "1111100100001010",
47422 => "1111100100001010",
47423 => "1111100100001011",
47424 => "1111100100001011",
47425 => "1111100100001100",
47426 => "1111100100001100",
47427 => "1111100100001101",
47428 => "1111100100001101",
47429 => "1111100100001101",
47430 => "1111100100001110",
47431 => "1111100100001110",
47432 => "1111100100001111",
47433 => "1111100100001111",
47434 => "1111100100001111",
47435 => "1111100100010000",
47436 => "1111100100010000",
47437 => "1111100100010001",
47438 => "1111100100010001",
47439 => "1111100100010010",
47440 => "1111100100010010",
47441 => "1111100100010010",
47442 => "1111100100010011",
47443 => "1111100100010011",
47444 => "1111100100010100",
47445 => "1111100100010100",
47446 => "1111100100010101",
47447 => "1111100100010101",
47448 => "1111100100010101",
47449 => "1111100100010110",
47450 => "1111100100010110",
47451 => "1111100100010111",
47452 => "1111100100010111",
47453 => "1111100100010111",
47454 => "1111100100011000",
47455 => "1111100100011000",
47456 => "1111100100011001",
47457 => "1111100100011001",
47458 => "1111100100011010",
47459 => "1111100100011010",
47460 => "1111100100011010",
47461 => "1111100100011011",
47462 => "1111100100011011",
47463 => "1111100100011100",
47464 => "1111100100011100",
47465 => "1111100100011100",
47466 => "1111100100011101",
47467 => "1111100100011101",
47468 => "1111100100011110",
47469 => "1111100100011110",
47470 => "1111100100011111",
47471 => "1111100100011111",
47472 => "1111100100011111",
47473 => "1111100100100000",
47474 => "1111100100100000",
47475 => "1111100100100001",
47476 => "1111100100100001",
47477 => "1111100100100010",
47478 => "1111100100100010",
47479 => "1111100100100010",
47480 => "1111100100100011",
47481 => "1111100100100011",
47482 => "1111100100100100",
47483 => "1111100100100100",
47484 => "1111100100100100",
47485 => "1111100100100101",
47486 => "1111100100100101",
47487 => "1111100100100110",
47488 => "1111100100100110",
47489 => "1111100100100111",
47490 => "1111100100100111",
47491 => "1111100100100111",
47492 => "1111100100101000",
47493 => "1111100100101000",
47494 => "1111100100101001",
47495 => "1111100100101001",
47496 => "1111100100101001",
47497 => "1111100100101010",
47498 => "1111100100101010",
47499 => "1111100100101011",
47500 => "1111100100101011",
47501 => "1111100100101100",
47502 => "1111100100101100",
47503 => "1111100100101100",
47504 => "1111100100101101",
47505 => "1111100100101101",
47506 => "1111100100101110",
47507 => "1111100100101110",
47508 => "1111100100101110",
47509 => "1111100100101111",
47510 => "1111100100101111",
47511 => "1111100100110000",
47512 => "1111100100110000",
47513 => "1111100100110000",
47514 => "1111100100110001",
47515 => "1111100100110001",
47516 => "1111100100110010",
47517 => "1111100100110010",
47518 => "1111100100110011",
47519 => "1111100100110011",
47520 => "1111100100110011",
47521 => "1111100100110100",
47522 => "1111100100110100",
47523 => "1111100100110101",
47524 => "1111100100110101",
47525 => "1111100100110101",
47526 => "1111100100110110",
47527 => "1111100100110110",
47528 => "1111100100110111",
47529 => "1111100100110111",
47530 => "1111100100111000",
47531 => "1111100100111000",
47532 => "1111100100111000",
47533 => "1111100100111001",
47534 => "1111100100111001",
47535 => "1111100100111010",
47536 => "1111100100111010",
47537 => "1111100100111010",
47538 => "1111100100111011",
47539 => "1111100100111011",
47540 => "1111100100111100",
47541 => "1111100100111100",
47542 => "1111100100111100",
47543 => "1111100100111101",
47544 => "1111100100111101",
47545 => "1111100100111110",
47546 => "1111100100111110",
47547 => "1111100100111111",
47548 => "1111100100111111",
47549 => "1111100100111111",
47550 => "1111100101000000",
47551 => "1111100101000000",
47552 => "1111100101000001",
47553 => "1111100101000001",
47554 => "1111100101000001",
47555 => "1111100101000010",
47556 => "1111100101000010",
47557 => "1111100101000011",
47558 => "1111100101000011",
47559 => "1111100101000011",
47560 => "1111100101000100",
47561 => "1111100101000100",
47562 => "1111100101000101",
47563 => "1111100101000101",
47564 => "1111100101000101",
47565 => "1111100101000110",
47566 => "1111100101000110",
47567 => "1111100101000111",
47568 => "1111100101000111",
47569 => "1111100101001000",
47570 => "1111100101001000",
47571 => "1111100101001000",
47572 => "1111100101001001",
47573 => "1111100101001001",
47574 => "1111100101001010",
47575 => "1111100101001010",
47576 => "1111100101001010",
47577 => "1111100101001011",
47578 => "1111100101001011",
47579 => "1111100101001100",
47580 => "1111100101001100",
47581 => "1111100101001100",
47582 => "1111100101001101",
47583 => "1111100101001101",
47584 => "1111100101001110",
47585 => "1111100101001110",
47586 => "1111100101001110",
47587 => "1111100101001111",
47588 => "1111100101001111",
47589 => "1111100101010000",
47590 => "1111100101010000",
47591 => "1111100101010001",
47592 => "1111100101010001",
47593 => "1111100101010001",
47594 => "1111100101010010",
47595 => "1111100101010010",
47596 => "1111100101010011",
47597 => "1111100101010011",
47598 => "1111100101010011",
47599 => "1111100101010100",
47600 => "1111100101010100",
47601 => "1111100101010101",
47602 => "1111100101010101",
47603 => "1111100101010101",
47604 => "1111100101010110",
47605 => "1111100101010110",
47606 => "1111100101010111",
47607 => "1111100101010111",
47608 => "1111100101010111",
47609 => "1111100101011000",
47610 => "1111100101011000",
47611 => "1111100101011001",
47612 => "1111100101011001",
47613 => "1111100101011001",
47614 => "1111100101011010",
47615 => "1111100101011010",
47616 => "1111100101011011",
47617 => "1111100101011011",
47618 => "1111100101011011",
47619 => "1111100101011100",
47620 => "1111100101011100",
47621 => "1111100101011101",
47622 => "1111100101011101",
47623 => "1111100101011101",
47624 => "1111100101011110",
47625 => "1111100101011110",
47626 => "1111100101011111",
47627 => "1111100101011111",
47628 => "1111100101011111",
47629 => "1111100101100000",
47630 => "1111100101100000",
47631 => "1111100101100001",
47632 => "1111100101100001",
47633 => "1111100101100010",
47634 => "1111100101100010",
47635 => "1111100101100010",
47636 => "1111100101100011",
47637 => "1111100101100011",
47638 => "1111100101100100",
47639 => "1111100101100100",
47640 => "1111100101100100",
47641 => "1111100101100101",
47642 => "1111100101100101",
47643 => "1111100101100110",
47644 => "1111100101100110",
47645 => "1111100101100110",
47646 => "1111100101100111",
47647 => "1111100101100111",
47648 => "1111100101101000",
47649 => "1111100101101000",
47650 => "1111100101101000",
47651 => "1111100101101001",
47652 => "1111100101101001",
47653 => "1111100101101010",
47654 => "1111100101101010",
47655 => "1111100101101010",
47656 => "1111100101101011",
47657 => "1111100101101011",
47658 => "1111100101101100",
47659 => "1111100101101100",
47660 => "1111100101101100",
47661 => "1111100101101101",
47662 => "1111100101101101",
47663 => "1111100101101110",
47664 => "1111100101101110",
47665 => "1111100101101110",
47666 => "1111100101101111",
47667 => "1111100101101111",
47668 => "1111100101110000",
47669 => "1111100101110000",
47670 => "1111100101110000",
47671 => "1111100101110001",
47672 => "1111100101110001",
47673 => "1111100101110010",
47674 => "1111100101110010",
47675 => "1111100101110010",
47676 => "1111100101110011",
47677 => "1111100101110011",
47678 => "1111100101110100",
47679 => "1111100101110100",
47680 => "1111100101110100",
47681 => "1111100101110101",
47682 => "1111100101110101",
47683 => "1111100101110110",
47684 => "1111100101110110",
47685 => "1111100101110110",
47686 => "1111100101110111",
47687 => "1111100101110111",
47688 => "1111100101111000",
47689 => "1111100101111000",
47690 => "1111100101111000",
47691 => "1111100101111001",
47692 => "1111100101111001",
47693 => "1111100101111010",
47694 => "1111100101111010",
47695 => "1111100101111010",
47696 => "1111100101111011",
47697 => "1111100101111011",
47698 => "1111100101111100",
47699 => "1111100101111100",
47700 => "1111100101111100",
47701 => "1111100101111101",
47702 => "1111100101111101",
47703 => "1111100101111101",
47704 => "1111100101111110",
47705 => "1111100101111110",
47706 => "1111100101111111",
47707 => "1111100101111111",
47708 => "1111100101111111",
47709 => "1111100110000000",
47710 => "1111100110000000",
47711 => "1111100110000001",
47712 => "1111100110000001",
47713 => "1111100110000001",
47714 => "1111100110000010",
47715 => "1111100110000010",
47716 => "1111100110000011",
47717 => "1111100110000011",
47718 => "1111100110000011",
47719 => "1111100110000100",
47720 => "1111100110000100",
47721 => "1111100110000101",
47722 => "1111100110000101",
47723 => "1111100110000101",
47724 => "1111100110000110",
47725 => "1111100110000110",
47726 => "1111100110000111",
47727 => "1111100110000111",
47728 => "1111100110000111",
47729 => "1111100110001000",
47730 => "1111100110001000",
47731 => "1111100110001001",
47732 => "1111100110001001",
47733 => "1111100110001001",
47734 => "1111100110001010",
47735 => "1111100110001010",
47736 => "1111100110001011",
47737 => "1111100110001011",
47738 => "1111100110001011",
47739 => "1111100110001100",
47740 => "1111100110001100",
47741 => "1111100110001100",
47742 => "1111100110001101",
47743 => "1111100110001101",
47744 => "1111100110001110",
47745 => "1111100110001110",
47746 => "1111100110001110",
47747 => "1111100110001111",
47748 => "1111100110001111",
47749 => "1111100110010000",
47750 => "1111100110010000",
47751 => "1111100110010000",
47752 => "1111100110010001",
47753 => "1111100110010001",
47754 => "1111100110010010",
47755 => "1111100110010010",
47756 => "1111100110010010",
47757 => "1111100110010011",
47758 => "1111100110010011",
47759 => "1111100110010100",
47760 => "1111100110010100",
47761 => "1111100110010100",
47762 => "1111100110010101",
47763 => "1111100110010101",
47764 => "1111100110010110",
47765 => "1111100110010110",
47766 => "1111100110010110",
47767 => "1111100110010111",
47768 => "1111100110010111",
47769 => "1111100110010111",
47770 => "1111100110011000",
47771 => "1111100110011000",
47772 => "1111100110011001",
47773 => "1111100110011001",
47774 => "1111100110011001",
47775 => "1111100110011010",
47776 => "1111100110011010",
47777 => "1111100110011011",
47778 => "1111100110011011",
47779 => "1111100110011011",
47780 => "1111100110011100",
47781 => "1111100110011100",
47782 => "1111100110011101",
47783 => "1111100110011101",
47784 => "1111100110011101",
47785 => "1111100110011110",
47786 => "1111100110011110",
47787 => "1111100110011110",
47788 => "1111100110011111",
47789 => "1111100110011111",
47790 => "1111100110100000",
47791 => "1111100110100000",
47792 => "1111100110100000",
47793 => "1111100110100001",
47794 => "1111100110100001",
47795 => "1111100110100010",
47796 => "1111100110100010",
47797 => "1111100110100010",
47798 => "1111100110100011",
47799 => "1111100110100011",
47800 => "1111100110100100",
47801 => "1111100110100100",
47802 => "1111100110100100",
47803 => "1111100110100101",
47804 => "1111100110100101",
47805 => "1111100110100101",
47806 => "1111100110100110",
47807 => "1111100110100110",
47808 => "1111100110100111",
47809 => "1111100110100111",
47810 => "1111100110100111",
47811 => "1111100110101000",
47812 => "1111100110101000",
47813 => "1111100110101001",
47814 => "1111100110101001",
47815 => "1111100110101001",
47816 => "1111100110101010",
47817 => "1111100110101010",
47818 => "1111100110101010",
47819 => "1111100110101011",
47820 => "1111100110101011",
47821 => "1111100110101100",
47822 => "1111100110101100",
47823 => "1111100110101100",
47824 => "1111100110101101",
47825 => "1111100110101101",
47826 => "1111100110101110",
47827 => "1111100110101110",
47828 => "1111100110101110",
47829 => "1111100110101111",
47830 => "1111100110101111",
47831 => "1111100110101111",
47832 => "1111100110110000",
47833 => "1111100110110000",
47834 => "1111100110110001",
47835 => "1111100110110001",
47836 => "1111100110110001",
47837 => "1111100110110010",
47838 => "1111100110110010",
47839 => "1111100110110011",
47840 => "1111100110110011",
47841 => "1111100110110011",
47842 => "1111100110110100",
47843 => "1111100110110100",
47844 => "1111100110110100",
47845 => "1111100110110101",
47846 => "1111100110110101",
47847 => "1111100110110110",
47848 => "1111100110110110",
47849 => "1111100110110110",
47850 => "1111100110110111",
47851 => "1111100110110111",
47852 => "1111100110111000",
47853 => "1111100110111000",
47854 => "1111100110111000",
47855 => "1111100110111001",
47856 => "1111100110111001",
47857 => "1111100110111001",
47858 => "1111100110111010",
47859 => "1111100110111010",
47860 => "1111100110111011",
47861 => "1111100110111011",
47862 => "1111100110111011",
47863 => "1111100110111100",
47864 => "1111100110111100",
47865 => "1111100110111101",
47866 => "1111100110111101",
47867 => "1111100110111101",
47868 => "1111100110111110",
47869 => "1111100110111110",
47870 => "1111100110111110",
47871 => "1111100110111111",
47872 => "1111100110111111",
47873 => "1111100111000000",
47874 => "1111100111000000",
47875 => "1111100111000000",
47876 => "1111100111000001",
47877 => "1111100111000001",
47878 => "1111100111000001",
47879 => "1111100111000010",
47880 => "1111100111000010",
47881 => "1111100111000011",
47882 => "1111100111000011",
47883 => "1111100111000011",
47884 => "1111100111000100",
47885 => "1111100111000100",
47886 => "1111100111000101",
47887 => "1111100111000101",
47888 => "1111100111000101",
47889 => "1111100111000110",
47890 => "1111100111000110",
47891 => "1111100111000110",
47892 => "1111100111000111",
47893 => "1111100111000111",
47894 => "1111100111001000",
47895 => "1111100111001000",
47896 => "1111100111001000",
47897 => "1111100111001001",
47898 => "1111100111001001",
47899 => "1111100111001001",
47900 => "1111100111001010",
47901 => "1111100111001010",
47902 => "1111100111001011",
47903 => "1111100111001011",
47904 => "1111100111001011",
47905 => "1111100111001100",
47906 => "1111100111001100",
47907 => "1111100111001100",
47908 => "1111100111001101",
47909 => "1111100111001101",
47910 => "1111100111001110",
47911 => "1111100111001110",
47912 => "1111100111001110",
47913 => "1111100111001111",
47914 => "1111100111001111",
47915 => "1111100111001111",
47916 => "1111100111010000",
47917 => "1111100111010000",
47918 => "1111100111010001",
47919 => "1111100111010001",
47920 => "1111100111010001",
47921 => "1111100111010010",
47922 => "1111100111010010",
47923 => "1111100111010011",
47924 => "1111100111010011",
47925 => "1111100111010011",
47926 => "1111100111010100",
47927 => "1111100111010100",
47928 => "1111100111010100",
47929 => "1111100111010101",
47930 => "1111100111010101",
47931 => "1111100111010110",
47932 => "1111100111010110",
47933 => "1111100111010110",
47934 => "1111100111010111",
47935 => "1111100111010111",
47936 => "1111100111010111",
47937 => "1111100111011000",
47938 => "1111100111011000",
47939 => "1111100111011001",
47940 => "1111100111011001",
47941 => "1111100111011001",
47942 => "1111100111011010",
47943 => "1111100111011010",
47944 => "1111100111011010",
47945 => "1111100111011011",
47946 => "1111100111011011",
47947 => "1111100111011100",
47948 => "1111100111011100",
47949 => "1111100111011100",
47950 => "1111100111011101",
47951 => "1111100111011101",
47952 => "1111100111011101",
47953 => "1111100111011110",
47954 => "1111100111011110",
47955 => "1111100111011111",
47956 => "1111100111011111",
47957 => "1111100111011111",
47958 => "1111100111100000",
47959 => "1111100111100000",
47960 => "1111100111100000",
47961 => "1111100111100001",
47962 => "1111100111100001",
47963 => "1111100111100010",
47964 => "1111100111100010",
47965 => "1111100111100010",
47966 => "1111100111100011",
47967 => "1111100111100011",
47968 => "1111100111100011",
47969 => "1111100111100100",
47970 => "1111100111100100",
47971 => "1111100111100100",
47972 => "1111100111100101",
47973 => "1111100111100101",
47974 => "1111100111100110",
47975 => "1111100111100110",
47976 => "1111100111100110",
47977 => "1111100111100111",
47978 => "1111100111100111",
47979 => "1111100111100111",
47980 => "1111100111101000",
47981 => "1111100111101000",
47982 => "1111100111101001",
47983 => "1111100111101001",
47984 => "1111100111101001",
47985 => "1111100111101010",
47986 => "1111100111101010",
47987 => "1111100111101010",
47988 => "1111100111101011",
47989 => "1111100111101011",
47990 => "1111100111101100",
47991 => "1111100111101100",
47992 => "1111100111101100",
47993 => "1111100111101101",
47994 => "1111100111101101",
47995 => "1111100111101101",
47996 => "1111100111101110",
47997 => "1111100111101110",
47998 => "1111100111101111",
47999 => "1111100111101111",
48000 => "1111100111101111",
48001 => "1111100111110000",
48002 => "1111100111110000",
48003 => "1111100111110000",
48004 => "1111100111110001",
48005 => "1111100111110001",
48006 => "1111100111110001",
48007 => "1111100111110010",
48008 => "1111100111110010",
48009 => "1111100111110011",
48010 => "1111100111110011",
48011 => "1111100111110011",
48012 => "1111100111110100",
48013 => "1111100111110100",
48014 => "1111100111110100",
48015 => "1111100111110101",
48016 => "1111100111110101",
48017 => "1111100111110110",
48018 => "1111100111110110",
48019 => "1111100111110110",
48020 => "1111100111110111",
48021 => "1111100111110111",
48022 => "1111100111110111",
48023 => "1111100111111000",
48024 => "1111100111111000",
48025 => "1111100111111000",
48026 => "1111100111111001",
48027 => "1111100111111001",
48028 => "1111100111111010",
48029 => "1111100111111010",
48030 => "1111100111111010",
48031 => "1111100111111011",
48032 => "1111100111111011",
48033 => "1111100111111011",
48034 => "1111100111111100",
48035 => "1111100111111100",
48036 => "1111100111111101",
48037 => "1111100111111101",
48038 => "1111100111111101",
48039 => "1111100111111110",
48040 => "1111100111111110",
48041 => "1111100111111110",
48042 => "1111100111111111",
48043 => "1111100111111111",
48044 => "1111100111111111",
48045 => "1111101000000000",
48046 => "1111101000000000",
48047 => "1111101000000001",
48048 => "1111101000000001",
48049 => "1111101000000001",
48050 => "1111101000000010",
48051 => "1111101000000010",
48052 => "1111101000000010",
48053 => "1111101000000011",
48054 => "1111101000000011",
48055 => "1111101000000011",
48056 => "1111101000000100",
48057 => "1111101000000100",
48058 => "1111101000000101",
48059 => "1111101000000101",
48060 => "1111101000000101",
48061 => "1111101000000110",
48062 => "1111101000000110",
48063 => "1111101000000110",
48064 => "1111101000000111",
48065 => "1111101000000111",
48066 => "1111101000000111",
48067 => "1111101000001000",
48068 => "1111101000001000",
48069 => "1111101000001001",
48070 => "1111101000001001",
48071 => "1111101000001001",
48072 => "1111101000001010",
48073 => "1111101000001010",
48074 => "1111101000001010",
48075 => "1111101000001011",
48076 => "1111101000001011",
48077 => "1111101000001011",
48078 => "1111101000001100",
48079 => "1111101000001100",
48080 => "1111101000001101",
48081 => "1111101000001101",
48082 => "1111101000001101",
48083 => "1111101000001110",
48084 => "1111101000001110",
48085 => "1111101000001110",
48086 => "1111101000001111",
48087 => "1111101000001111",
48088 => "1111101000001111",
48089 => "1111101000010000",
48090 => "1111101000010000",
48091 => "1111101000010001",
48092 => "1111101000010001",
48093 => "1111101000010001",
48094 => "1111101000010010",
48095 => "1111101000010010",
48096 => "1111101000010010",
48097 => "1111101000010011",
48098 => "1111101000010011",
48099 => "1111101000010011",
48100 => "1111101000010100",
48101 => "1111101000010100",
48102 => "1111101000010101",
48103 => "1111101000010101",
48104 => "1111101000010101",
48105 => "1111101000010110",
48106 => "1111101000010110",
48107 => "1111101000010110",
48108 => "1111101000010111",
48109 => "1111101000010111",
48110 => "1111101000010111",
48111 => "1111101000011000",
48112 => "1111101000011000",
48113 => "1111101000011001",
48114 => "1111101000011001",
48115 => "1111101000011001",
48116 => "1111101000011010",
48117 => "1111101000011010",
48118 => "1111101000011010",
48119 => "1111101000011011",
48120 => "1111101000011011",
48121 => "1111101000011011",
48122 => "1111101000011100",
48123 => "1111101000011100",
48124 => "1111101000011100",
48125 => "1111101000011101",
48126 => "1111101000011101",
48127 => "1111101000011110",
48128 => "1111101000011110",
48129 => "1111101000011110",
48130 => "1111101000011111",
48131 => "1111101000011111",
48132 => "1111101000011111",
48133 => "1111101000100000",
48134 => "1111101000100000",
48135 => "1111101000100000",
48136 => "1111101000100001",
48137 => "1111101000100001",
48138 => "1111101000100010",
48139 => "1111101000100010",
48140 => "1111101000100010",
48141 => "1111101000100011",
48142 => "1111101000100011",
48143 => "1111101000100011",
48144 => "1111101000100100",
48145 => "1111101000100100",
48146 => "1111101000100100",
48147 => "1111101000100101",
48148 => "1111101000100101",
48149 => "1111101000100101",
48150 => "1111101000100110",
48151 => "1111101000100110",
48152 => "1111101000100111",
48153 => "1111101000100111",
48154 => "1111101000100111",
48155 => "1111101000101000",
48156 => "1111101000101000",
48157 => "1111101000101000",
48158 => "1111101000101001",
48159 => "1111101000101001",
48160 => "1111101000101001",
48161 => "1111101000101010",
48162 => "1111101000101010",
48163 => "1111101000101010",
48164 => "1111101000101011",
48165 => "1111101000101011",
48166 => "1111101000101100",
48167 => "1111101000101100",
48168 => "1111101000101100",
48169 => "1111101000101101",
48170 => "1111101000101101",
48171 => "1111101000101101",
48172 => "1111101000101110",
48173 => "1111101000101110",
48174 => "1111101000101110",
48175 => "1111101000101111",
48176 => "1111101000101111",
48177 => "1111101000101111",
48178 => "1111101000110000",
48179 => "1111101000110000",
48180 => "1111101000110000",
48181 => "1111101000110001",
48182 => "1111101000110001",
48183 => "1111101000110010",
48184 => "1111101000110010",
48185 => "1111101000110010",
48186 => "1111101000110011",
48187 => "1111101000110011",
48188 => "1111101000110011",
48189 => "1111101000110100",
48190 => "1111101000110100",
48191 => "1111101000110100",
48192 => "1111101000110101",
48193 => "1111101000110101",
48194 => "1111101000110101",
48195 => "1111101000110110",
48196 => "1111101000110110",
48197 => "1111101000110111",
48198 => "1111101000110111",
48199 => "1111101000110111",
48200 => "1111101000111000",
48201 => "1111101000111000",
48202 => "1111101000111000",
48203 => "1111101000111001",
48204 => "1111101000111001",
48205 => "1111101000111001",
48206 => "1111101000111010",
48207 => "1111101000111010",
48208 => "1111101000111010",
48209 => "1111101000111011",
48210 => "1111101000111011",
48211 => "1111101000111011",
48212 => "1111101000111100",
48213 => "1111101000111100",
48214 => "1111101000111100",
48215 => "1111101000111101",
48216 => "1111101000111101",
48217 => "1111101000111110",
48218 => "1111101000111110",
48219 => "1111101000111110",
48220 => "1111101000111111",
48221 => "1111101000111111",
48222 => "1111101000111111",
48223 => "1111101001000000",
48224 => "1111101001000000",
48225 => "1111101001000000",
48226 => "1111101001000001",
48227 => "1111101001000001",
48228 => "1111101001000001",
48229 => "1111101001000010",
48230 => "1111101001000010",
48231 => "1111101001000010",
48232 => "1111101001000011",
48233 => "1111101001000011",
48234 => "1111101001000100",
48235 => "1111101001000100",
48236 => "1111101001000100",
48237 => "1111101001000101",
48238 => "1111101001000101",
48239 => "1111101001000101",
48240 => "1111101001000110",
48241 => "1111101001000110",
48242 => "1111101001000110",
48243 => "1111101001000111",
48244 => "1111101001000111",
48245 => "1111101001000111",
48246 => "1111101001001000",
48247 => "1111101001001000",
48248 => "1111101001001000",
48249 => "1111101001001001",
48250 => "1111101001001001",
48251 => "1111101001001001",
48252 => "1111101001001010",
48253 => "1111101001001010",
48254 => "1111101001001011",
48255 => "1111101001001011",
48256 => "1111101001001011",
48257 => "1111101001001100",
48258 => "1111101001001100",
48259 => "1111101001001100",
48260 => "1111101001001101",
48261 => "1111101001001101",
48262 => "1111101001001101",
48263 => "1111101001001110",
48264 => "1111101001001110",
48265 => "1111101001001110",
48266 => "1111101001001111",
48267 => "1111101001001111",
48268 => "1111101001001111",
48269 => "1111101001010000",
48270 => "1111101001010000",
48271 => "1111101001010000",
48272 => "1111101001010001",
48273 => "1111101001010001",
48274 => "1111101001010001",
48275 => "1111101001010010",
48276 => "1111101001010010",
48277 => "1111101001010011",
48278 => "1111101001010011",
48279 => "1111101001010011",
48280 => "1111101001010100",
48281 => "1111101001010100",
48282 => "1111101001010100",
48283 => "1111101001010101",
48284 => "1111101001010101",
48285 => "1111101001010101",
48286 => "1111101001010110",
48287 => "1111101001010110",
48288 => "1111101001010110",
48289 => "1111101001010111",
48290 => "1111101001010111",
48291 => "1111101001010111",
48292 => "1111101001011000",
48293 => "1111101001011000",
48294 => "1111101001011000",
48295 => "1111101001011001",
48296 => "1111101001011001",
48297 => "1111101001011001",
48298 => "1111101001011010",
48299 => "1111101001011010",
48300 => "1111101001011010",
48301 => "1111101001011011",
48302 => "1111101001011011",
48303 => "1111101001011100",
48304 => "1111101001011100",
48305 => "1111101001011100",
48306 => "1111101001011101",
48307 => "1111101001011101",
48308 => "1111101001011101",
48309 => "1111101001011110",
48310 => "1111101001011110",
48311 => "1111101001011110",
48312 => "1111101001011111",
48313 => "1111101001011111",
48314 => "1111101001011111",
48315 => "1111101001100000",
48316 => "1111101001100000",
48317 => "1111101001100000",
48318 => "1111101001100001",
48319 => "1111101001100001",
48320 => "1111101001100001",
48321 => "1111101001100010",
48322 => "1111101001100010",
48323 => "1111101001100010",
48324 => "1111101001100011",
48325 => "1111101001100011",
48326 => "1111101001100011",
48327 => "1111101001100100",
48328 => "1111101001100100",
48329 => "1111101001100100",
48330 => "1111101001100101",
48331 => "1111101001100101",
48332 => "1111101001100101",
48333 => "1111101001100110",
48334 => "1111101001100110",
48335 => "1111101001100110",
48336 => "1111101001100111",
48337 => "1111101001100111",
48338 => "1111101001101000",
48339 => "1111101001101000",
48340 => "1111101001101000",
48341 => "1111101001101001",
48342 => "1111101001101001",
48343 => "1111101001101001",
48344 => "1111101001101010",
48345 => "1111101001101010",
48346 => "1111101001101010",
48347 => "1111101001101011",
48348 => "1111101001101011",
48349 => "1111101001101011",
48350 => "1111101001101100",
48351 => "1111101001101100",
48352 => "1111101001101100",
48353 => "1111101001101101",
48354 => "1111101001101101",
48355 => "1111101001101101",
48356 => "1111101001101110",
48357 => "1111101001101110",
48358 => "1111101001101110",
48359 => "1111101001101111",
48360 => "1111101001101111",
48361 => "1111101001101111",
48362 => "1111101001110000",
48363 => "1111101001110000",
48364 => "1111101001110000",
48365 => "1111101001110001",
48366 => "1111101001110001",
48367 => "1111101001110001",
48368 => "1111101001110010",
48369 => "1111101001110010",
48370 => "1111101001110010",
48371 => "1111101001110011",
48372 => "1111101001110011",
48373 => "1111101001110011",
48374 => "1111101001110100",
48375 => "1111101001110100",
48376 => "1111101001110100",
48377 => "1111101001110101",
48378 => "1111101001110101",
48379 => "1111101001110101",
48380 => "1111101001110110",
48381 => "1111101001110110",
48382 => "1111101001110110",
48383 => "1111101001110111",
48384 => "1111101001110111",
48385 => "1111101001111000",
48386 => "1111101001111000",
48387 => "1111101001111000",
48388 => "1111101001111001",
48389 => "1111101001111001",
48390 => "1111101001111001",
48391 => "1111101001111010",
48392 => "1111101001111010",
48393 => "1111101001111010",
48394 => "1111101001111011",
48395 => "1111101001111011",
48396 => "1111101001111011",
48397 => "1111101001111100",
48398 => "1111101001111100",
48399 => "1111101001111100",
48400 => "1111101001111101",
48401 => "1111101001111101",
48402 => "1111101001111101",
48403 => "1111101001111110",
48404 => "1111101001111110",
48405 => "1111101001111110",
48406 => "1111101001111111",
48407 => "1111101001111111",
48408 => "1111101001111111",
48409 => "1111101010000000",
48410 => "1111101010000000",
48411 => "1111101010000000",
48412 => "1111101010000001",
48413 => "1111101010000001",
48414 => "1111101010000001",
48415 => "1111101010000010",
48416 => "1111101010000010",
48417 => "1111101010000010",
48418 => "1111101010000011",
48419 => "1111101010000011",
48420 => "1111101010000011",
48421 => "1111101010000100",
48422 => "1111101010000100",
48423 => "1111101010000100",
48424 => "1111101010000101",
48425 => "1111101010000101",
48426 => "1111101010000101",
48427 => "1111101010000110",
48428 => "1111101010000110",
48429 => "1111101010000110",
48430 => "1111101010000111",
48431 => "1111101010000111",
48432 => "1111101010000111",
48433 => "1111101010001000",
48434 => "1111101010001000",
48435 => "1111101010001000",
48436 => "1111101010001001",
48437 => "1111101010001001",
48438 => "1111101010001001",
48439 => "1111101010001010",
48440 => "1111101010001010",
48441 => "1111101010001010",
48442 => "1111101010001011",
48443 => "1111101010001011",
48444 => "1111101010001011",
48445 => "1111101010001100",
48446 => "1111101010001100",
48447 => "1111101010001100",
48448 => "1111101010001101",
48449 => "1111101010001101",
48450 => "1111101010001101",
48451 => "1111101010001110",
48452 => "1111101010001110",
48453 => "1111101010001110",
48454 => "1111101010001111",
48455 => "1111101010001111",
48456 => "1111101010001111",
48457 => "1111101010010000",
48458 => "1111101010010000",
48459 => "1111101010010000",
48460 => "1111101010010001",
48461 => "1111101010010001",
48462 => "1111101010010001",
48463 => "1111101010010010",
48464 => "1111101010010010",
48465 => "1111101010010010",
48466 => "1111101010010011",
48467 => "1111101010010011",
48468 => "1111101010010011",
48469 => "1111101010010100",
48470 => "1111101010010100",
48471 => "1111101010010100",
48472 => "1111101010010101",
48473 => "1111101010010101",
48474 => "1111101010010101",
48475 => "1111101010010110",
48476 => "1111101010010110",
48477 => "1111101010010110",
48478 => "1111101010010111",
48479 => "1111101010010111",
48480 => "1111101010010111",
48481 => "1111101010011000",
48482 => "1111101010011000",
48483 => "1111101010011000",
48484 => "1111101010011001",
48485 => "1111101010011001",
48486 => "1111101010011001",
48487 => "1111101010011010",
48488 => "1111101010011010",
48489 => "1111101010011010",
48490 => "1111101010011011",
48491 => "1111101010011011",
48492 => "1111101010011011",
48493 => "1111101010011100",
48494 => "1111101010011100",
48495 => "1111101010011100",
48496 => "1111101010011101",
48497 => "1111101010011101",
48498 => "1111101010011101",
48499 => "1111101010011110",
48500 => "1111101010011110",
48501 => "1111101010011110",
48502 => "1111101010011111",
48503 => "1111101010011111",
48504 => "1111101010011111",
48505 => "1111101010100000",
48506 => "1111101010100000",
48507 => "1111101010100000",
48508 => "1111101010100001",
48509 => "1111101010100001",
48510 => "1111101010100001",
48511 => "1111101010100010",
48512 => "1111101010100010",
48513 => "1111101010100010",
48514 => "1111101010100010",
48515 => "1111101010100011",
48516 => "1111101010100011",
48517 => "1111101010100011",
48518 => "1111101010100100",
48519 => "1111101010100100",
48520 => "1111101010100100",
48521 => "1111101010100101",
48522 => "1111101010100101",
48523 => "1111101010100101",
48524 => "1111101010100110",
48525 => "1111101010100110",
48526 => "1111101010100110",
48527 => "1111101010100111",
48528 => "1111101010100111",
48529 => "1111101010100111",
48530 => "1111101010101000",
48531 => "1111101010101000",
48532 => "1111101010101000",
48533 => "1111101010101001",
48534 => "1111101010101001",
48535 => "1111101010101001",
48536 => "1111101010101010",
48537 => "1111101010101010",
48538 => "1111101010101010",
48539 => "1111101010101011",
48540 => "1111101010101011",
48541 => "1111101010101011",
48542 => "1111101010101100",
48543 => "1111101010101100",
48544 => "1111101010101100",
48545 => "1111101010101101",
48546 => "1111101010101101",
48547 => "1111101010101101",
48548 => "1111101010101110",
48549 => "1111101010101110",
48550 => "1111101010101110",
48551 => "1111101010101111",
48552 => "1111101010101111",
48553 => "1111101010101111",
48554 => "1111101010110000",
48555 => "1111101010110000",
48556 => "1111101010110000",
48557 => "1111101010110001",
48558 => "1111101010110001",
48559 => "1111101010110001",
48560 => "1111101010110010",
48561 => "1111101010110010",
48562 => "1111101010110010",
48563 => "1111101010110010",
48564 => "1111101010110011",
48565 => "1111101010110011",
48566 => "1111101010110011",
48567 => "1111101010110100",
48568 => "1111101010110100",
48569 => "1111101010110100",
48570 => "1111101010110101",
48571 => "1111101010110101",
48572 => "1111101010110101",
48573 => "1111101010110110",
48574 => "1111101010110110",
48575 => "1111101010110110",
48576 => "1111101010110111",
48577 => "1111101010110111",
48578 => "1111101010110111",
48579 => "1111101010111000",
48580 => "1111101010111000",
48581 => "1111101010111000",
48582 => "1111101010111001",
48583 => "1111101010111001",
48584 => "1111101010111001",
48585 => "1111101010111010",
48586 => "1111101010111010",
48587 => "1111101010111010",
48588 => "1111101010111011",
48589 => "1111101010111011",
48590 => "1111101010111011",
48591 => "1111101010111100",
48592 => "1111101010111100",
48593 => "1111101010111100",
48594 => "1111101010111100",
48595 => "1111101010111101",
48596 => "1111101010111101",
48597 => "1111101010111101",
48598 => "1111101010111110",
48599 => "1111101010111110",
48600 => "1111101010111110",
48601 => "1111101010111111",
48602 => "1111101010111111",
48603 => "1111101010111111",
48604 => "1111101011000000",
48605 => "1111101011000000",
48606 => "1111101011000000",
48607 => "1111101011000001",
48608 => "1111101011000001",
48609 => "1111101011000001",
48610 => "1111101011000010",
48611 => "1111101011000010",
48612 => "1111101011000010",
48613 => "1111101011000011",
48614 => "1111101011000011",
48615 => "1111101011000011",
48616 => "1111101011000100",
48617 => "1111101011000100",
48618 => "1111101011000100",
48619 => "1111101011000101",
48620 => "1111101011000101",
48621 => "1111101011000101",
48622 => "1111101011000101",
48623 => "1111101011000110",
48624 => "1111101011000110",
48625 => "1111101011000110",
48626 => "1111101011000111",
48627 => "1111101011000111",
48628 => "1111101011000111",
48629 => "1111101011001000",
48630 => "1111101011001000",
48631 => "1111101011001000",
48632 => "1111101011001001",
48633 => "1111101011001001",
48634 => "1111101011001001",
48635 => "1111101011001010",
48636 => "1111101011001010",
48637 => "1111101011001010",
48638 => "1111101011001011",
48639 => "1111101011001011",
48640 => "1111101011001011",
48641 => "1111101011001100",
48642 => "1111101011001100",
48643 => "1111101011001100",
48644 => "1111101011001101",
48645 => "1111101011001101",
48646 => "1111101011001101",
48647 => "1111101011001101",
48648 => "1111101011001110",
48649 => "1111101011001110",
48650 => "1111101011001110",
48651 => "1111101011001111",
48652 => "1111101011001111",
48653 => "1111101011001111",
48654 => "1111101011010000",
48655 => "1111101011010000",
48656 => "1111101011010000",
48657 => "1111101011010001",
48658 => "1111101011010001",
48659 => "1111101011010001",
48660 => "1111101011010010",
48661 => "1111101011010010",
48662 => "1111101011010010",
48663 => "1111101011010011",
48664 => "1111101011010011",
48665 => "1111101011010011",
48666 => "1111101011010011",
48667 => "1111101011010100",
48668 => "1111101011010100",
48669 => "1111101011010100",
48670 => "1111101011010101",
48671 => "1111101011010101",
48672 => "1111101011010101",
48673 => "1111101011010110",
48674 => "1111101011010110",
48675 => "1111101011010110",
48676 => "1111101011010111",
48677 => "1111101011010111",
48678 => "1111101011010111",
48679 => "1111101011011000",
48680 => "1111101011011000",
48681 => "1111101011011000",
48682 => "1111101011011001",
48683 => "1111101011011001",
48684 => "1111101011011001",
48685 => "1111101011011001",
48686 => "1111101011011010",
48687 => "1111101011011010",
48688 => "1111101011011010",
48689 => "1111101011011011",
48690 => "1111101011011011",
48691 => "1111101011011011",
48692 => "1111101011011100",
48693 => "1111101011011100",
48694 => "1111101011011100",
48695 => "1111101011011101",
48696 => "1111101011011101",
48697 => "1111101011011101",
48698 => "1111101011011110",
48699 => "1111101011011110",
48700 => "1111101011011110",
48701 => "1111101011011111",
48702 => "1111101011011111",
48703 => "1111101011011111",
48704 => "1111101011011111",
48705 => "1111101011100000",
48706 => "1111101011100000",
48707 => "1111101011100000",
48708 => "1111101011100001",
48709 => "1111101011100001",
48710 => "1111101011100001",
48711 => "1111101011100010",
48712 => "1111101011100010",
48713 => "1111101011100010",
48714 => "1111101011100011",
48715 => "1111101011100011",
48716 => "1111101011100011",
48717 => "1111101011100100",
48718 => "1111101011100100",
48719 => "1111101011100100",
48720 => "1111101011100100",
48721 => "1111101011100101",
48722 => "1111101011100101",
48723 => "1111101011100101",
48724 => "1111101011100110",
48725 => "1111101011100110",
48726 => "1111101011100110",
48727 => "1111101011100111",
48728 => "1111101011100111",
48729 => "1111101011100111",
48730 => "1111101011101000",
48731 => "1111101011101000",
48732 => "1111101011101000",
48733 => "1111101011101001",
48734 => "1111101011101001",
48735 => "1111101011101001",
48736 => "1111101011101001",
48737 => "1111101011101010",
48738 => "1111101011101010",
48739 => "1111101011101010",
48740 => "1111101011101011",
48741 => "1111101011101011",
48742 => "1111101011101011",
48743 => "1111101011101100",
48744 => "1111101011101100",
48745 => "1111101011101100",
48746 => "1111101011101101",
48747 => "1111101011101101",
48748 => "1111101011101101",
48749 => "1111101011101110",
48750 => "1111101011101110",
48751 => "1111101011101110",
48752 => "1111101011101110",
48753 => "1111101011101111",
48754 => "1111101011101111",
48755 => "1111101011101111",
48756 => "1111101011110000",
48757 => "1111101011110000",
48758 => "1111101011110000",
48759 => "1111101011110001",
48760 => "1111101011110001",
48761 => "1111101011110001",
48762 => "1111101011110010",
48763 => "1111101011110010",
48764 => "1111101011110010",
48765 => "1111101011110010",
48766 => "1111101011110011",
48767 => "1111101011110011",
48768 => "1111101011110011",
48769 => "1111101011110100",
48770 => "1111101011110100",
48771 => "1111101011110100",
48772 => "1111101011110101",
48773 => "1111101011110101",
48774 => "1111101011110101",
48775 => "1111101011110110",
48776 => "1111101011110110",
48777 => "1111101011110110",
48778 => "1111101011110111",
48779 => "1111101011110111",
48780 => "1111101011110111",
48781 => "1111101011110111",
48782 => "1111101011111000",
48783 => "1111101011111000",
48784 => "1111101011111000",
48785 => "1111101011111001",
48786 => "1111101011111001",
48787 => "1111101011111001",
48788 => "1111101011111010",
48789 => "1111101011111010",
48790 => "1111101011111010",
48791 => "1111101011111011",
48792 => "1111101011111011",
48793 => "1111101011111011",
48794 => "1111101011111011",
48795 => "1111101011111100",
48796 => "1111101011111100",
48797 => "1111101011111100",
48798 => "1111101011111101",
48799 => "1111101011111101",
48800 => "1111101011111101",
48801 => "1111101011111110",
48802 => "1111101011111110",
48803 => "1111101011111110",
48804 => "1111101011111111",
48805 => "1111101011111111",
48806 => "1111101011111111",
48807 => "1111101011111111",
48808 => "1111101100000000",
48809 => "1111101100000000",
48810 => "1111101100000000",
48811 => "1111101100000001",
48812 => "1111101100000001",
48813 => "1111101100000001",
48814 => "1111101100000010",
48815 => "1111101100000010",
48816 => "1111101100000010",
48817 => "1111101100000010",
48818 => "1111101100000011",
48819 => "1111101100000011",
48820 => "1111101100000011",
48821 => "1111101100000100",
48822 => "1111101100000100",
48823 => "1111101100000100",
48824 => "1111101100000101",
48825 => "1111101100000101",
48826 => "1111101100000101",
48827 => "1111101100000110",
48828 => "1111101100000110",
48829 => "1111101100000110",
48830 => "1111101100000110",
48831 => "1111101100000111",
48832 => "1111101100000111",
48833 => "1111101100000111",
48834 => "1111101100001000",
48835 => "1111101100001000",
48836 => "1111101100001000",
48837 => "1111101100001001",
48838 => "1111101100001001",
48839 => "1111101100001001",
48840 => "1111101100001001",
48841 => "1111101100001010",
48842 => "1111101100001010",
48843 => "1111101100001010",
48844 => "1111101100001011",
48845 => "1111101100001011",
48846 => "1111101100001011",
48847 => "1111101100001100",
48848 => "1111101100001100",
48849 => "1111101100001100",
48850 => "1111101100001101",
48851 => "1111101100001101",
48852 => "1111101100001101",
48853 => "1111101100001101",
48854 => "1111101100001110",
48855 => "1111101100001110",
48856 => "1111101100001110",
48857 => "1111101100001111",
48858 => "1111101100001111",
48859 => "1111101100001111",
48860 => "1111101100010000",
48861 => "1111101100010000",
48862 => "1111101100010000",
48863 => "1111101100010000",
48864 => "1111101100010001",
48865 => "1111101100010001",
48866 => "1111101100010001",
48867 => "1111101100010010",
48868 => "1111101100010010",
48869 => "1111101100010010",
48870 => "1111101100010011",
48871 => "1111101100010011",
48872 => "1111101100010011",
48873 => "1111101100010011",
48874 => "1111101100010100",
48875 => "1111101100010100",
48876 => "1111101100010100",
48877 => "1111101100010101",
48878 => "1111101100010101",
48879 => "1111101100010101",
48880 => "1111101100010110",
48881 => "1111101100010110",
48882 => "1111101100010110",
48883 => "1111101100010111",
48884 => "1111101100010111",
48885 => "1111101100010111",
48886 => "1111101100010111",
48887 => "1111101100011000",
48888 => "1111101100011000",
48889 => "1111101100011000",
48890 => "1111101100011001",
48891 => "1111101100011001",
48892 => "1111101100011001",
48893 => "1111101100011010",
48894 => "1111101100011010",
48895 => "1111101100011010",
48896 => "1111101100011010",
48897 => "1111101100011011",
48898 => "1111101100011011",
48899 => "1111101100011011",
48900 => "1111101100011100",
48901 => "1111101100011100",
48902 => "1111101100011100",
48903 => "1111101100011101",
48904 => "1111101100011101",
48905 => "1111101100011101",
48906 => "1111101100011101",
48907 => "1111101100011110",
48908 => "1111101100011110",
48909 => "1111101100011110",
48910 => "1111101100011111",
48911 => "1111101100011111",
48912 => "1111101100011111",
48913 => "1111101100100000",
48914 => "1111101100100000",
48915 => "1111101100100000",
48916 => "1111101100100000",
48917 => "1111101100100001",
48918 => "1111101100100001",
48919 => "1111101100100001",
48920 => "1111101100100010",
48921 => "1111101100100010",
48922 => "1111101100100010",
48923 => "1111101100100010",
48924 => "1111101100100011",
48925 => "1111101100100011",
48926 => "1111101100100011",
48927 => "1111101100100100",
48928 => "1111101100100100",
48929 => "1111101100100100",
48930 => "1111101100100101",
48931 => "1111101100100101",
48932 => "1111101100100101",
48933 => "1111101100100101",
48934 => "1111101100100110",
48935 => "1111101100100110",
48936 => "1111101100100110",
48937 => "1111101100100111",
48938 => "1111101100100111",
48939 => "1111101100100111",
48940 => "1111101100101000",
48941 => "1111101100101000",
48942 => "1111101100101000",
48943 => "1111101100101000",
48944 => "1111101100101001",
48945 => "1111101100101001",
48946 => "1111101100101001",
48947 => "1111101100101010",
48948 => "1111101100101010",
48949 => "1111101100101010",
48950 => "1111101100101011",
48951 => "1111101100101011",
48952 => "1111101100101011",
48953 => "1111101100101011",
48954 => "1111101100101100",
48955 => "1111101100101100",
48956 => "1111101100101100",
48957 => "1111101100101101",
48958 => "1111101100101101",
48959 => "1111101100101101",
48960 => "1111101100101101",
48961 => "1111101100101110",
48962 => "1111101100101110",
48963 => "1111101100101110",
48964 => "1111101100101111",
48965 => "1111101100101111",
48966 => "1111101100101111",
48967 => "1111101100110000",
48968 => "1111101100110000",
48969 => "1111101100110000",
48970 => "1111101100110000",
48971 => "1111101100110001",
48972 => "1111101100110001",
48973 => "1111101100110001",
48974 => "1111101100110010",
48975 => "1111101100110010",
48976 => "1111101100110010",
48977 => "1111101100110010",
48978 => "1111101100110011",
48979 => "1111101100110011",
48980 => "1111101100110011",
48981 => "1111101100110100",
48982 => "1111101100110100",
48983 => "1111101100110100",
48984 => "1111101100110101",
48985 => "1111101100110101",
48986 => "1111101100110101",
48987 => "1111101100110101",
48988 => "1111101100110110",
48989 => "1111101100110110",
48990 => "1111101100110110",
48991 => "1111101100110111",
48992 => "1111101100110111",
48993 => "1111101100110111",
48994 => "1111101100110111",
48995 => "1111101100111000",
48996 => "1111101100111000",
48997 => "1111101100111000",
48998 => "1111101100111001",
48999 => "1111101100111001",
49000 => "1111101100111001",
49001 => "1111101100111010",
49002 => "1111101100111010",
49003 => "1111101100111010",
49004 => "1111101100111010",
49005 => "1111101100111011",
49006 => "1111101100111011",
49007 => "1111101100111011",
49008 => "1111101100111100",
49009 => "1111101100111100",
49010 => "1111101100111100",
49011 => "1111101100111100",
49012 => "1111101100111101",
49013 => "1111101100111101",
49014 => "1111101100111101",
49015 => "1111101100111110",
49016 => "1111101100111110",
49017 => "1111101100111110",
49018 => "1111101100111111",
49019 => "1111101100111111",
49020 => "1111101100111111",
49021 => "1111101100111111",
49022 => "1111101101000000",
49023 => "1111101101000000",
49024 => "1111101101000000",
49025 => "1111101101000001",
49026 => "1111101101000001",
49027 => "1111101101000001",
49028 => "1111101101000001",
49029 => "1111101101000010",
49030 => "1111101101000010",
49031 => "1111101101000010",
49032 => "1111101101000011",
49033 => "1111101101000011",
49034 => "1111101101000011",
49035 => "1111101101000011",
49036 => "1111101101000100",
49037 => "1111101101000100",
49038 => "1111101101000100",
49039 => "1111101101000101",
49040 => "1111101101000101",
49041 => "1111101101000101",
49042 => "1111101101000101",
49043 => "1111101101000110",
49044 => "1111101101000110",
49045 => "1111101101000110",
49046 => "1111101101000111",
49047 => "1111101101000111",
49048 => "1111101101000111",
49049 => "1111101101001000",
49050 => "1111101101001000",
49051 => "1111101101001000",
49052 => "1111101101001000",
49053 => "1111101101001001",
49054 => "1111101101001001",
49055 => "1111101101001001",
49056 => "1111101101001010",
49057 => "1111101101001010",
49058 => "1111101101001010",
49059 => "1111101101001010",
49060 => "1111101101001011",
49061 => "1111101101001011",
49062 => "1111101101001011",
49063 => "1111101101001100",
49064 => "1111101101001100",
49065 => "1111101101001100",
49066 => "1111101101001100",
49067 => "1111101101001101",
49068 => "1111101101001101",
49069 => "1111101101001101",
49070 => "1111101101001110",
49071 => "1111101101001110",
49072 => "1111101101001110",
49073 => "1111101101001110",
49074 => "1111101101001111",
49075 => "1111101101001111",
49076 => "1111101101001111",
49077 => "1111101101010000",
49078 => "1111101101010000",
49079 => "1111101101010000",
49080 => "1111101101010000",
49081 => "1111101101010001",
49082 => "1111101101010001",
49083 => "1111101101010001",
49084 => "1111101101010010",
49085 => "1111101101010010",
49086 => "1111101101010010",
49087 => "1111101101010010",
49088 => "1111101101010011",
49089 => "1111101101010011",
49090 => "1111101101010011",
49091 => "1111101101010100",
49092 => "1111101101010100",
49093 => "1111101101010100",
49094 => "1111101101010100",
49095 => "1111101101010101",
49096 => "1111101101010101",
49097 => "1111101101010101",
49098 => "1111101101010110",
49099 => "1111101101010110",
49100 => "1111101101010110",
49101 => "1111101101010110",
49102 => "1111101101010111",
49103 => "1111101101010111",
49104 => "1111101101010111",
49105 => "1111101101011000",
49106 => "1111101101011000",
49107 => "1111101101011000",
49108 => "1111101101011000",
49109 => "1111101101011001",
49110 => "1111101101011001",
49111 => "1111101101011001",
49112 => "1111101101011010",
49113 => "1111101101011010",
49114 => "1111101101011010",
49115 => "1111101101011010",
49116 => "1111101101011011",
49117 => "1111101101011011",
49118 => "1111101101011011",
49119 => "1111101101011100",
49120 => "1111101101011100",
49121 => "1111101101011100",
49122 => "1111101101011100",
49123 => "1111101101011101",
49124 => "1111101101011101",
49125 => "1111101101011101",
49126 => "1111101101011110",
49127 => "1111101101011110",
49128 => "1111101101011110",
49129 => "1111101101011110",
49130 => "1111101101011111",
49131 => "1111101101011111",
49132 => "1111101101011111",
49133 => "1111101101100000",
49134 => "1111101101100000",
49135 => "1111101101100000",
49136 => "1111101101100000",
49137 => "1111101101100001",
49138 => "1111101101100001",
49139 => "1111101101100001",
49140 => "1111101101100010",
49141 => "1111101101100010",
49142 => "1111101101100010",
49143 => "1111101101100010",
49144 => "1111101101100011",
49145 => "1111101101100011",
49146 => "1111101101100011",
49147 => "1111101101100100",
49148 => "1111101101100100",
49149 => "1111101101100100",
49150 => "1111101101100100",
49151 => "1111101101100101",
49152 => "1111101101100101",
49153 => "1111101101100101",
49154 => "1111101101100110",
49155 => "1111101101100110",
49156 => "1111101101100110",
49157 => "1111101101100110",
49158 => "1111101101100111",
49159 => "1111101101100111",
49160 => "1111101101100111",
49161 => "1111101101101000",
49162 => "1111101101101000",
49163 => "1111101101101000",
49164 => "1111101101101000",
49165 => "1111101101101001",
49166 => "1111101101101001",
49167 => "1111101101101001",
49168 => "1111101101101001",
49169 => "1111101101101010",
49170 => "1111101101101010",
49171 => "1111101101101010",
49172 => "1111101101101011",
49173 => "1111101101101011",
49174 => "1111101101101011",
49175 => "1111101101101011",
49176 => "1111101101101100",
49177 => "1111101101101100",
49178 => "1111101101101100",
49179 => "1111101101101101",
49180 => "1111101101101101",
49181 => "1111101101101101",
49182 => "1111101101101101",
49183 => "1111101101101110",
49184 => "1111101101101110",
49185 => "1111101101101110",
49186 => "1111101101101111",
49187 => "1111101101101111",
49188 => "1111101101101111",
49189 => "1111101101101111",
49190 => "1111101101110000",
49191 => "1111101101110000",
49192 => "1111101101110000",
49193 => "1111101101110000",
49194 => "1111101101110001",
49195 => "1111101101110001",
49196 => "1111101101110001",
49197 => "1111101101110010",
49198 => "1111101101110010",
49199 => "1111101101110010",
49200 => "1111101101110010",
49201 => "1111101101110011",
49202 => "1111101101110011",
49203 => "1111101101110011",
49204 => "1111101101110100",
49205 => "1111101101110100",
49206 => "1111101101110100",
49207 => "1111101101110100",
49208 => "1111101101110101",
49209 => "1111101101110101",
49210 => "1111101101110101",
49211 => "1111101101110110",
49212 => "1111101101110110",
49213 => "1111101101110110",
49214 => "1111101101110110",
49215 => "1111101101110111",
49216 => "1111101101110111",
49217 => "1111101101110111",
49218 => "1111101101110111",
49219 => "1111101101111000",
49220 => "1111101101111000",
49221 => "1111101101111000",
49222 => "1111101101111001",
49223 => "1111101101111001",
49224 => "1111101101111001",
49225 => "1111101101111001",
49226 => "1111101101111010",
49227 => "1111101101111010",
49228 => "1111101101111010",
49229 => "1111101101111011",
49230 => "1111101101111011",
49231 => "1111101101111011",
49232 => "1111101101111011",
49233 => "1111101101111100",
49234 => "1111101101111100",
49235 => "1111101101111100",
49236 => "1111101101111100",
49237 => "1111101101111101",
49238 => "1111101101111101",
49239 => "1111101101111101",
49240 => "1111101101111110",
49241 => "1111101101111110",
49242 => "1111101101111110",
49243 => "1111101101111110",
49244 => "1111101101111111",
49245 => "1111101101111111",
49246 => "1111101101111111",
49247 => "1111101110000000",
49248 => "1111101110000000",
49249 => "1111101110000000",
49250 => "1111101110000000",
49251 => "1111101110000001",
49252 => "1111101110000001",
49253 => "1111101110000001",
49254 => "1111101110000001",
49255 => "1111101110000010",
49256 => "1111101110000010",
49257 => "1111101110000010",
49258 => "1111101110000011",
49259 => "1111101110000011",
49260 => "1111101110000011",
49261 => "1111101110000011",
49262 => "1111101110000100",
49263 => "1111101110000100",
49264 => "1111101110000100",
49265 => "1111101110000100",
49266 => "1111101110000101",
49267 => "1111101110000101",
49268 => "1111101110000101",
49269 => "1111101110000110",
49270 => "1111101110000110",
49271 => "1111101110000110",
49272 => "1111101110000110",
49273 => "1111101110000111",
49274 => "1111101110000111",
49275 => "1111101110000111",
49276 => "1111101110000111",
49277 => "1111101110001000",
49278 => "1111101110001000",
49279 => "1111101110001000",
49280 => "1111101110001001",
49281 => "1111101110001001",
49282 => "1111101110001001",
49283 => "1111101110001001",
49284 => "1111101110001010",
49285 => "1111101110001010",
49286 => "1111101110001010",
49287 => "1111101110001011",
49288 => "1111101110001011",
49289 => "1111101110001011",
49290 => "1111101110001011",
49291 => "1111101110001100",
49292 => "1111101110001100",
49293 => "1111101110001100",
49294 => "1111101110001100",
49295 => "1111101110001101",
49296 => "1111101110001101",
49297 => "1111101110001101",
49298 => "1111101110001110",
49299 => "1111101110001110",
49300 => "1111101110001110",
49301 => "1111101110001110",
49302 => "1111101110001111",
49303 => "1111101110001111",
49304 => "1111101110001111",
49305 => "1111101110001111",
49306 => "1111101110010000",
49307 => "1111101110010000",
49308 => "1111101110010000",
49309 => "1111101110010001",
49310 => "1111101110010001",
49311 => "1111101110010001",
49312 => "1111101110010001",
49313 => "1111101110010010",
49314 => "1111101110010010",
49315 => "1111101110010010",
49316 => "1111101110010010",
49317 => "1111101110010011",
49318 => "1111101110010011",
49319 => "1111101110010011",
49320 => "1111101110010100",
49321 => "1111101110010100",
49322 => "1111101110010100",
49323 => "1111101110010100",
49324 => "1111101110010101",
49325 => "1111101110010101",
49326 => "1111101110010101",
49327 => "1111101110010101",
49328 => "1111101110010110",
49329 => "1111101110010110",
49330 => "1111101110010110",
49331 => "1111101110010110",
49332 => "1111101110010111",
49333 => "1111101110010111",
49334 => "1111101110010111",
49335 => "1111101110011000",
49336 => "1111101110011000",
49337 => "1111101110011000",
49338 => "1111101110011000",
49339 => "1111101110011001",
49340 => "1111101110011001",
49341 => "1111101110011001",
49342 => "1111101110011001",
49343 => "1111101110011010",
49344 => "1111101110011010",
49345 => "1111101110011010",
49346 => "1111101110011011",
49347 => "1111101110011011",
49348 => "1111101110011011",
49349 => "1111101110011011",
49350 => "1111101110011100",
49351 => "1111101110011100",
49352 => "1111101110011100",
49353 => "1111101110011100",
49354 => "1111101110011101",
49355 => "1111101110011101",
49356 => "1111101110011101",
49357 => "1111101110011110",
49358 => "1111101110011110",
49359 => "1111101110011110",
49360 => "1111101110011110",
49361 => "1111101110011111",
49362 => "1111101110011111",
49363 => "1111101110011111",
49364 => "1111101110011111",
49365 => "1111101110100000",
49366 => "1111101110100000",
49367 => "1111101110100000",
49368 => "1111101110100000",
49369 => "1111101110100001",
49370 => "1111101110100001",
49371 => "1111101110100001",
49372 => "1111101110100010",
49373 => "1111101110100010",
49374 => "1111101110100010",
49375 => "1111101110100010",
49376 => "1111101110100011",
49377 => "1111101110100011",
49378 => "1111101110100011",
49379 => "1111101110100011",
49380 => "1111101110100100",
49381 => "1111101110100100",
49382 => "1111101110100100",
49383 => "1111101110100100",
49384 => "1111101110100101",
49385 => "1111101110100101",
49386 => "1111101110100101",
49387 => "1111101110100110",
49388 => "1111101110100110",
49389 => "1111101110100110",
49390 => "1111101110100110",
49391 => "1111101110100111",
49392 => "1111101110100111",
49393 => "1111101110100111",
49394 => "1111101110100111",
49395 => "1111101110101000",
49396 => "1111101110101000",
49397 => "1111101110101000",
49398 => "1111101110101001",
49399 => "1111101110101001",
49400 => "1111101110101001",
49401 => "1111101110101001",
49402 => "1111101110101010",
49403 => "1111101110101010",
49404 => "1111101110101010",
49405 => "1111101110101010",
49406 => "1111101110101011",
49407 => "1111101110101011",
49408 => "1111101110101011",
49409 => "1111101110101011",
49410 => "1111101110101100",
49411 => "1111101110101100",
49412 => "1111101110101100",
49413 => "1111101110101100",
49414 => "1111101110101101",
49415 => "1111101110101101",
49416 => "1111101110101101",
49417 => "1111101110101110",
49418 => "1111101110101110",
49419 => "1111101110101110",
49420 => "1111101110101110",
49421 => "1111101110101111",
49422 => "1111101110101111",
49423 => "1111101110101111",
49424 => "1111101110101111",
49425 => "1111101110110000",
49426 => "1111101110110000",
49427 => "1111101110110000",
49428 => "1111101110110000",
49429 => "1111101110110001",
49430 => "1111101110110001",
49431 => "1111101110110001",
49432 => "1111101110110010",
49433 => "1111101110110010",
49434 => "1111101110110010",
49435 => "1111101110110010",
49436 => "1111101110110011",
49437 => "1111101110110011",
49438 => "1111101110110011",
49439 => "1111101110110011",
49440 => "1111101110110100",
49441 => "1111101110110100",
49442 => "1111101110110100",
49443 => "1111101110110100",
49444 => "1111101110110101",
49445 => "1111101110110101",
49446 => "1111101110110101",
49447 => "1111101110110101",
49448 => "1111101110110110",
49449 => "1111101110110110",
49450 => "1111101110110110",
49451 => "1111101110110111",
49452 => "1111101110110111",
49453 => "1111101110110111",
49454 => "1111101110110111",
49455 => "1111101110111000",
49456 => "1111101110111000",
49457 => "1111101110111000",
49458 => "1111101110111000",
49459 => "1111101110111001",
49460 => "1111101110111001",
49461 => "1111101110111001",
49462 => "1111101110111001",
49463 => "1111101110111010",
49464 => "1111101110111010",
49465 => "1111101110111010",
49466 => "1111101110111010",
49467 => "1111101110111011",
49468 => "1111101110111011",
49469 => "1111101110111011",
49470 => "1111101110111100",
49471 => "1111101110111100",
49472 => "1111101110111100",
49473 => "1111101110111100",
49474 => "1111101110111101",
49475 => "1111101110111101",
49476 => "1111101110111101",
49477 => "1111101110111101",
49478 => "1111101110111110",
49479 => "1111101110111110",
49480 => "1111101110111110",
49481 => "1111101110111110",
49482 => "1111101110111111",
49483 => "1111101110111111",
49484 => "1111101110111111",
49485 => "1111101110111111",
49486 => "1111101111000000",
49487 => "1111101111000000",
49488 => "1111101111000000",
49489 => "1111101111000001",
49490 => "1111101111000001",
49491 => "1111101111000001",
49492 => "1111101111000001",
49493 => "1111101111000010",
49494 => "1111101111000010",
49495 => "1111101111000010",
49496 => "1111101111000010",
49497 => "1111101111000011",
49498 => "1111101111000011",
49499 => "1111101111000011",
49500 => "1111101111000011",
49501 => "1111101111000100",
49502 => "1111101111000100",
49503 => "1111101111000100",
49504 => "1111101111000100",
49505 => "1111101111000101",
49506 => "1111101111000101",
49507 => "1111101111000101",
49508 => "1111101111000101",
49509 => "1111101111000110",
49510 => "1111101111000110",
49511 => "1111101111000110",
49512 => "1111101111000110",
49513 => "1111101111000111",
49514 => "1111101111000111",
49515 => "1111101111000111",
49516 => "1111101111001000",
49517 => "1111101111001000",
49518 => "1111101111001000",
49519 => "1111101111001000",
49520 => "1111101111001001",
49521 => "1111101111001001",
49522 => "1111101111001001",
49523 => "1111101111001001",
49524 => "1111101111001010",
49525 => "1111101111001010",
49526 => "1111101111001010",
49527 => "1111101111001010",
49528 => "1111101111001011",
49529 => "1111101111001011",
49530 => "1111101111001011",
49531 => "1111101111001011",
49532 => "1111101111001100",
49533 => "1111101111001100",
49534 => "1111101111001100",
49535 => "1111101111001100",
49536 => "1111101111001101",
49537 => "1111101111001101",
49538 => "1111101111001101",
49539 => "1111101111001101",
49540 => "1111101111001110",
49541 => "1111101111001110",
49542 => "1111101111001110",
49543 => "1111101111001111",
49544 => "1111101111001111",
49545 => "1111101111001111",
49546 => "1111101111001111",
49547 => "1111101111010000",
49548 => "1111101111010000",
49549 => "1111101111010000",
49550 => "1111101111010000",
49551 => "1111101111010001",
49552 => "1111101111010001",
49553 => "1111101111010001",
49554 => "1111101111010001",
49555 => "1111101111010010",
49556 => "1111101111010010",
49557 => "1111101111010010",
49558 => "1111101111010010",
49559 => "1111101111010011",
49560 => "1111101111010011",
49561 => "1111101111010011",
49562 => "1111101111010011",
49563 => "1111101111010100",
49564 => "1111101111010100",
49565 => "1111101111010100",
49566 => "1111101111010100",
49567 => "1111101111010101",
49568 => "1111101111010101",
49569 => "1111101111010101",
49570 => "1111101111010101",
49571 => "1111101111010110",
49572 => "1111101111010110",
49573 => "1111101111010110",
49574 => "1111101111010110",
49575 => "1111101111010111",
49576 => "1111101111010111",
49577 => "1111101111010111",
49578 => "1111101111010111",
49579 => "1111101111011000",
49580 => "1111101111011000",
49581 => "1111101111011000",
49582 => "1111101111011001",
49583 => "1111101111011001",
49584 => "1111101111011001",
49585 => "1111101111011001",
49586 => "1111101111011010",
49587 => "1111101111011010",
49588 => "1111101111011010",
49589 => "1111101111011010",
49590 => "1111101111011011",
49591 => "1111101111011011",
49592 => "1111101111011011",
49593 => "1111101111011011",
49594 => "1111101111011100",
49595 => "1111101111011100",
49596 => "1111101111011100",
49597 => "1111101111011100",
49598 => "1111101111011101",
49599 => "1111101111011101",
49600 => "1111101111011101",
49601 => "1111101111011101",
49602 => "1111101111011110",
49603 => "1111101111011110",
49604 => "1111101111011110",
49605 => "1111101111011110",
49606 => "1111101111011111",
49607 => "1111101111011111",
49608 => "1111101111011111",
49609 => "1111101111011111",
49610 => "1111101111100000",
49611 => "1111101111100000",
49612 => "1111101111100000",
49613 => "1111101111100000",
49614 => "1111101111100001",
49615 => "1111101111100001",
49616 => "1111101111100001",
49617 => "1111101111100001",
49618 => "1111101111100010",
49619 => "1111101111100010",
49620 => "1111101111100010",
49621 => "1111101111100010",
49622 => "1111101111100011",
49623 => "1111101111100011",
49624 => "1111101111100011",
49625 => "1111101111100011",
49626 => "1111101111100100",
49627 => "1111101111100100",
49628 => "1111101111100100",
49629 => "1111101111100100",
49630 => "1111101111100101",
49631 => "1111101111100101",
49632 => "1111101111100101",
49633 => "1111101111100101",
49634 => "1111101111100110",
49635 => "1111101111100110",
49636 => "1111101111100110",
49637 => "1111101111100110",
49638 => "1111101111100111",
49639 => "1111101111100111",
49640 => "1111101111100111",
49641 => "1111101111100111",
49642 => "1111101111101000",
49643 => "1111101111101000",
49644 => "1111101111101000",
49645 => "1111101111101000",
49646 => "1111101111101001",
49647 => "1111101111101001",
49648 => "1111101111101001",
49649 => "1111101111101001",
49650 => "1111101111101010",
49651 => "1111101111101010",
49652 => "1111101111101010",
49653 => "1111101111101010",
49654 => "1111101111101011",
49655 => "1111101111101011",
49656 => "1111101111101011",
49657 => "1111101111101011",
49658 => "1111101111101100",
49659 => "1111101111101100",
49660 => "1111101111101100",
49661 => "1111101111101100",
49662 => "1111101111101101",
49663 => "1111101111101101",
49664 => "1111101111101101",
49665 => "1111101111101101",
49666 => "1111101111101110",
49667 => "1111101111101110",
49668 => "1111101111101110",
49669 => "1111101111101110",
49670 => "1111101111101111",
49671 => "1111101111101111",
49672 => "1111101111101111",
49673 => "1111101111101111",
49674 => "1111101111110000",
49675 => "1111101111110000",
49676 => "1111101111110000",
49677 => "1111101111110000",
49678 => "1111101111110001",
49679 => "1111101111110001",
49680 => "1111101111110001",
49681 => "1111101111110001",
49682 => "1111101111110010",
49683 => "1111101111110010",
49684 => "1111101111110010",
49685 => "1111101111110010",
49686 => "1111101111110011",
49687 => "1111101111110011",
49688 => "1111101111110011",
49689 => "1111101111110011",
49690 => "1111101111110100",
49691 => "1111101111110100",
49692 => "1111101111110100",
49693 => "1111101111110100",
49694 => "1111101111110101",
49695 => "1111101111110101",
49696 => "1111101111110101",
49697 => "1111101111110101",
49698 => "1111101111110110",
49699 => "1111101111110110",
49700 => "1111101111110110",
49701 => "1111101111110110",
49702 => "1111101111110111",
49703 => "1111101111110111",
49704 => "1111101111110111",
49705 => "1111101111110111",
49706 => "1111101111111000",
49707 => "1111101111111000",
49708 => "1111101111111000",
49709 => "1111101111111000",
49710 => "1111101111111001",
49711 => "1111101111111001",
49712 => "1111101111111001",
49713 => "1111101111111001",
49714 => "1111101111111010",
49715 => "1111101111111010",
49716 => "1111101111111010",
49717 => "1111101111111010",
49718 => "1111101111111011",
49719 => "1111101111111011",
49720 => "1111101111111011",
49721 => "1111101111111011",
49722 => "1111101111111100",
49723 => "1111101111111100",
49724 => "1111101111111100",
49725 => "1111101111111100",
49726 => "1111101111111101",
49727 => "1111101111111101",
49728 => "1111101111111101",
49729 => "1111101111111101",
49730 => "1111101111111110",
49731 => "1111101111111110",
49732 => "1111101111111110",
49733 => "1111101111111110",
49734 => "1111101111111111",
49735 => "1111101111111111",
49736 => "1111101111111111",
49737 => "1111101111111111",
49738 => "1111110000000000",
49739 => "1111110000000000",
49740 => "1111110000000000",
49741 => "1111110000000000",
49742 => "1111110000000001",
49743 => "1111110000000001",
49744 => "1111110000000001",
49745 => "1111110000000001",
49746 => "1111110000000010",
49747 => "1111110000000010",
49748 => "1111110000000010",
49749 => "1111110000000010",
49750 => "1111110000000011",
49751 => "1111110000000011",
49752 => "1111110000000011",
49753 => "1111110000000011",
49754 => "1111110000000100",
49755 => "1111110000000100",
49756 => "1111110000000100",
49757 => "1111110000000100",
49758 => "1111110000000101",
49759 => "1111110000000101",
49760 => "1111110000000101",
49761 => "1111110000000101",
49762 => "1111110000000110",
49763 => "1111110000000110",
49764 => "1111110000000110",
49765 => "1111110000000110",
49766 => "1111110000000110",
49767 => "1111110000000111",
49768 => "1111110000000111",
49769 => "1111110000000111",
49770 => "1111110000000111",
49771 => "1111110000001000",
49772 => "1111110000001000",
49773 => "1111110000001000",
49774 => "1111110000001000",
49775 => "1111110000001001",
49776 => "1111110000001001",
49777 => "1111110000001001",
49778 => "1111110000001001",
49779 => "1111110000001010",
49780 => "1111110000001010",
49781 => "1111110000001010",
49782 => "1111110000001010",
49783 => "1111110000001011",
49784 => "1111110000001011",
49785 => "1111110000001011",
49786 => "1111110000001011",
49787 => "1111110000001100",
49788 => "1111110000001100",
49789 => "1111110000001100",
49790 => "1111110000001100",
49791 => "1111110000001101",
49792 => "1111110000001101",
49793 => "1111110000001101",
49794 => "1111110000001101",
49795 => "1111110000001110",
49796 => "1111110000001110",
49797 => "1111110000001110",
49798 => "1111110000001110",
49799 => "1111110000001111",
49800 => "1111110000001111",
49801 => "1111110000001111",
49802 => "1111110000001111",
49803 => "1111110000001111",
49804 => "1111110000010000",
49805 => "1111110000010000",
49806 => "1111110000010000",
49807 => "1111110000010000",
49808 => "1111110000010001",
49809 => "1111110000010001",
49810 => "1111110000010001",
49811 => "1111110000010001",
49812 => "1111110000010010",
49813 => "1111110000010010",
49814 => "1111110000010010",
49815 => "1111110000010010",
49816 => "1111110000010011",
49817 => "1111110000010011",
49818 => "1111110000010011",
49819 => "1111110000010011",
49820 => "1111110000010100",
49821 => "1111110000010100",
49822 => "1111110000010100",
49823 => "1111110000010100",
49824 => "1111110000010101",
49825 => "1111110000010101",
49826 => "1111110000010101",
49827 => "1111110000010101",
49828 => "1111110000010110",
49829 => "1111110000010110",
49830 => "1111110000010110",
49831 => "1111110000010110",
49832 => "1111110000010110",
49833 => "1111110000010111",
49834 => "1111110000010111",
49835 => "1111110000010111",
49836 => "1111110000010111",
49837 => "1111110000011000",
49838 => "1111110000011000",
49839 => "1111110000011000",
49840 => "1111110000011000",
49841 => "1111110000011001",
49842 => "1111110000011001",
49843 => "1111110000011001",
49844 => "1111110000011001",
49845 => "1111110000011010",
49846 => "1111110000011010",
49847 => "1111110000011010",
49848 => "1111110000011010",
49849 => "1111110000011011",
49850 => "1111110000011011",
49851 => "1111110000011011",
49852 => "1111110000011011",
49853 => "1111110000011100",
49854 => "1111110000011100",
49855 => "1111110000011100",
49856 => "1111110000011100",
49857 => "1111110000011100",
49858 => "1111110000011101",
49859 => "1111110000011101",
49860 => "1111110000011101",
49861 => "1111110000011101",
49862 => "1111110000011110",
49863 => "1111110000011110",
49864 => "1111110000011110",
49865 => "1111110000011110",
49866 => "1111110000011111",
49867 => "1111110000011111",
49868 => "1111110000011111",
49869 => "1111110000011111",
49870 => "1111110000100000",
49871 => "1111110000100000",
49872 => "1111110000100000",
49873 => "1111110000100000",
49874 => "1111110000100001",
49875 => "1111110000100001",
49876 => "1111110000100001",
49877 => "1111110000100001",
49878 => "1111110000100010",
49879 => "1111110000100010",
49880 => "1111110000100010",
49881 => "1111110000100010",
49882 => "1111110000100010",
49883 => "1111110000100011",
49884 => "1111110000100011",
49885 => "1111110000100011",
49886 => "1111110000100011",
49887 => "1111110000100100",
49888 => "1111110000100100",
49889 => "1111110000100100",
49890 => "1111110000100100",
49891 => "1111110000100101",
49892 => "1111110000100101",
49893 => "1111110000100101",
49894 => "1111110000100101",
49895 => "1111110000100110",
49896 => "1111110000100110",
49897 => "1111110000100110",
49898 => "1111110000100110",
49899 => "1111110000100110",
49900 => "1111110000100111",
49901 => "1111110000100111",
49902 => "1111110000100111",
49903 => "1111110000100111",
49904 => "1111110000101000",
49905 => "1111110000101000",
49906 => "1111110000101000",
49907 => "1111110000101000",
49908 => "1111110000101001",
49909 => "1111110000101001",
49910 => "1111110000101001",
49911 => "1111110000101001",
49912 => "1111110000101010",
49913 => "1111110000101010",
49914 => "1111110000101010",
49915 => "1111110000101010",
49916 => "1111110000101011",
49917 => "1111110000101011",
49918 => "1111110000101011",
49919 => "1111110000101011",
49920 => "1111110000101011",
49921 => "1111110000101100",
49922 => "1111110000101100",
49923 => "1111110000101100",
49924 => "1111110000101100",
49925 => "1111110000101101",
49926 => "1111110000101101",
49927 => "1111110000101101",
49928 => "1111110000101101",
49929 => "1111110000101110",
49930 => "1111110000101110",
49931 => "1111110000101110",
49932 => "1111110000101110",
49933 => "1111110000101111",
49934 => "1111110000101111",
49935 => "1111110000101111",
49936 => "1111110000101111",
49937 => "1111110000101111",
49938 => "1111110000110000",
49939 => "1111110000110000",
49940 => "1111110000110000",
49941 => "1111110000110000",
49942 => "1111110000110001",
49943 => "1111110000110001",
49944 => "1111110000110001",
49945 => "1111110000110001",
49946 => "1111110000110010",
49947 => "1111110000110010",
49948 => "1111110000110010",
49949 => "1111110000110010",
49950 => "1111110000110010",
49951 => "1111110000110011",
49952 => "1111110000110011",
49953 => "1111110000110011",
49954 => "1111110000110011",
49955 => "1111110000110100",
49956 => "1111110000110100",
49957 => "1111110000110100",
49958 => "1111110000110100",
49959 => "1111110000110101",
49960 => "1111110000110101",
49961 => "1111110000110101",
49962 => "1111110000110101",
49963 => "1111110000110110",
49964 => "1111110000110110",
49965 => "1111110000110110",
49966 => "1111110000110110",
49967 => "1111110000110110",
49968 => "1111110000110111",
49969 => "1111110000110111",
49970 => "1111110000110111",
49971 => "1111110000110111",
49972 => "1111110000111000",
49973 => "1111110000111000",
49974 => "1111110000111000",
49975 => "1111110000111000",
49976 => "1111110000111001",
49977 => "1111110000111001",
49978 => "1111110000111001",
49979 => "1111110000111001",
49980 => "1111110000111001",
49981 => "1111110000111010",
49982 => "1111110000111010",
49983 => "1111110000111010",
49984 => "1111110000111010",
49985 => "1111110000111011",
49986 => "1111110000111011",
49987 => "1111110000111011",
49988 => "1111110000111011",
49989 => "1111110000111100",
49990 => "1111110000111100",
49991 => "1111110000111100",
49992 => "1111110000111100",
49993 => "1111110000111101",
49994 => "1111110000111101",
49995 => "1111110000111101",
49996 => "1111110000111101",
49997 => "1111110000111101",
49998 => "1111110000111110",
49999 => "1111110000111110",
50000 => "1111110000111110",
50001 => "1111110000111110",
50002 => "1111110000111111",
50003 => "1111110000111111",
50004 => "1111110000111111",
50005 => "1111110000111111",
50006 => "1111110001000000",
50007 => "1111110001000000",
50008 => "1111110001000000",
50009 => "1111110001000000",
50010 => "1111110001000000",
50011 => "1111110001000001",
50012 => "1111110001000001",
50013 => "1111110001000001",
50014 => "1111110001000001",
50015 => "1111110001000010",
50016 => "1111110001000010",
50017 => "1111110001000010",
50018 => "1111110001000010",
50019 => "1111110001000011",
50020 => "1111110001000011",
50021 => "1111110001000011",
50022 => "1111110001000011",
50023 => "1111110001000011",
50024 => "1111110001000100",
50025 => "1111110001000100",
50026 => "1111110001000100",
50027 => "1111110001000100",
50028 => "1111110001000101",
50029 => "1111110001000101",
50030 => "1111110001000101",
50031 => "1111110001000101",
50032 => "1111110001000110",
50033 => "1111110001000110",
50034 => "1111110001000110",
50035 => "1111110001000110",
50036 => "1111110001000110",
50037 => "1111110001000111",
50038 => "1111110001000111",
50039 => "1111110001000111",
50040 => "1111110001000111",
50041 => "1111110001001000",
50042 => "1111110001001000",
50043 => "1111110001001000",
50044 => "1111110001001000",
50045 => "1111110001001000",
50046 => "1111110001001001",
50047 => "1111110001001001",
50048 => "1111110001001001",
50049 => "1111110001001001",
50050 => "1111110001001010",
50051 => "1111110001001010",
50052 => "1111110001001010",
50053 => "1111110001001010",
50054 => "1111110001001011",
50055 => "1111110001001011",
50056 => "1111110001001011",
50057 => "1111110001001011",
50058 => "1111110001001011",
50059 => "1111110001001100",
50060 => "1111110001001100",
50061 => "1111110001001100",
50062 => "1111110001001100",
50063 => "1111110001001101",
50064 => "1111110001001101",
50065 => "1111110001001101",
50066 => "1111110001001101",
50067 => "1111110001001110",
50068 => "1111110001001110",
50069 => "1111110001001110",
50070 => "1111110001001110",
50071 => "1111110001001110",
50072 => "1111110001001111",
50073 => "1111110001001111",
50074 => "1111110001001111",
50075 => "1111110001001111",
50076 => "1111110001010000",
50077 => "1111110001010000",
50078 => "1111110001010000",
50079 => "1111110001010000",
50080 => "1111110001010000",
50081 => "1111110001010001",
50082 => "1111110001010001",
50083 => "1111110001010001",
50084 => "1111110001010001",
50085 => "1111110001010010",
50086 => "1111110001010010",
50087 => "1111110001010010",
50088 => "1111110001010010",
50089 => "1111110001010010",
50090 => "1111110001010011",
50091 => "1111110001010011",
50092 => "1111110001010011",
50093 => "1111110001010011",
50094 => "1111110001010100",
50095 => "1111110001010100",
50096 => "1111110001010100",
50097 => "1111110001010100",
50098 => "1111110001010101",
50099 => "1111110001010101",
50100 => "1111110001010101",
50101 => "1111110001010101",
50102 => "1111110001010101",
50103 => "1111110001010110",
50104 => "1111110001010110",
50105 => "1111110001010110",
50106 => "1111110001010110",
50107 => "1111110001010111",
50108 => "1111110001010111",
50109 => "1111110001010111",
50110 => "1111110001010111",
50111 => "1111110001010111",
50112 => "1111110001011000",
50113 => "1111110001011000",
50114 => "1111110001011000",
50115 => "1111110001011000",
50116 => "1111110001011001",
50117 => "1111110001011001",
50118 => "1111110001011001",
50119 => "1111110001011001",
50120 => "1111110001011001",
50121 => "1111110001011010",
50122 => "1111110001011010",
50123 => "1111110001011010",
50124 => "1111110001011010",
50125 => "1111110001011011",
50126 => "1111110001011011",
50127 => "1111110001011011",
50128 => "1111110001011011",
50129 => "1111110001011100",
50130 => "1111110001011100",
50131 => "1111110001011100",
50132 => "1111110001011100",
50133 => "1111110001011100",
50134 => "1111110001011101",
50135 => "1111110001011101",
50136 => "1111110001011101",
50137 => "1111110001011101",
50138 => "1111110001011110",
50139 => "1111110001011110",
50140 => "1111110001011110",
50141 => "1111110001011110",
50142 => "1111110001011110",
50143 => "1111110001011111",
50144 => "1111110001011111",
50145 => "1111110001011111",
50146 => "1111110001011111",
50147 => "1111110001100000",
50148 => "1111110001100000",
50149 => "1111110001100000",
50150 => "1111110001100000",
50151 => "1111110001100000",
50152 => "1111110001100001",
50153 => "1111110001100001",
50154 => "1111110001100001",
50155 => "1111110001100001",
50156 => "1111110001100010",
50157 => "1111110001100010",
50158 => "1111110001100010",
50159 => "1111110001100010",
50160 => "1111110001100010",
50161 => "1111110001100011",
50162 => "1111110001100011",
50163 => "1111110001100011",
50164 => "1111110001100011",
50165 => "1111110001100100",
50166 => "1111110001100100",
50167 => "1111110001100100",
50168 => "1111110001100100",
50169 => "1111110001100100",
50170 => "1111110001100101",
50171 => "1111110001100101",
50172 => "1111110001100101",
50173 => "1111110001100101",
50174 => "1111110001100110",
50175 => "1111110001100110",
50176 => "1111110001100110",
50177 => "1111110001100110",
50178 => "1111110001100110",
50179 => "1111110001100111",
50180 => "1111110001100111",
50181 => "1111110001100111",
50182 => "1111110001100111",
50183 => "1111110001101000",
50184 => "1111110001101000",
50185 => "1111110001101000",
50186 => "1111110001101000",
50187 => "1111110001101000",
50188 => "1111110001101001",
50189 => "1111110001101001",
50190 => "1111110001101001",
50191 => "1111110001101001",
50192 => "1111110001101010",
50193 => "1111110001101010",
50194 => "1111110001101010",
50195 => "1111110001101010",
50196 => "1111110001101010",
50197 => "1111110001101011",
50198 => "1111110001101011",
50199 => "1111110001101011",
50200 => "1111110001101011",
50201 => "1111110001101100",
50202 => "1111110001101100",
50203 => "1111110001101100",
50204 => "1111110001101100",
50205 => "1111110001101100",
50206 => "1111110001101101",
50207 => "1111110001101101",
50208 => "1111110001101101",
50209 => "1111110001101101",
50210 => "1111110001101110",
50211 => "1111110001101110",
50212 => "1111110001101110",
50213 => "1111110001101110",
50214 => "1111110001101110",
50215 => "1111110001101111",
50216 => "1111110001101111",
50217 => "1111110001101111",
50218 => "1111110001101111",
50219 => "1111110001101111",
50220 => "1111110001110000",
50221 => "1111110001110000",
50222 => "1111110001110000",
50223 => "1111110001110000",
50224 => "1111110001110001",
50225 => "1111110001110001",
50226 => "1111110001110001",
50227 => "1111110001110001",
50228 => "1111110001110001",
50229 => "1111110001110010",
50230 => "1111110001110010",
50231 => "1111110001110010",
50232 => "1111110001110010",
50233 => "1111110001110011",
50234 => "1111110001110011",
50235 => "1111110001110011",
50236 => "1111110001110011",
50237 => "1111110001110011",
50238 => "1111110001110100",
50239 => "1111110001110100",
50240 => "1111110001110100",
50241 => "1111110001110100",
50242 => "1111110001110101",
50243 => "1111110001110101",
50244 => "1111110001110101",
50245 => "1111110001110101",
50246 => "1111110001110101",
50247 => "1111110001110110",
50248 => "1111110001110110",
50249 => "1111110001110110",
50250 => "1111110001110110",
50251 => "1111110001110110",
50252 => "1111110001110111",
50253 => "1111110001110111",
50254 => "1111110001110111",
50255 => "1111110001110111",
50256 => "1111110001111000",
50257 => "1111110001111000",
50258 => "1111110001111000",
50259 => "1111110001111000",
50260 => "1111110001111000",
50261 => "1111110001111001",
50262 => "1111110001111001",
50263 => "1111110001111001",
50264 => "1111110001111001",
50265 => "1111110001111010",
50266 => "1111110001111010",
50267 => "1111110001111010",
50268 => "1111110001111010",
50269 => "1111110001111010",
50270 => "1111110001111011",
50271 => "1111110001111011",
50272 => "1111110001111011",
50273 => "1111110001111011",
50274 => "1111110001111011",
50275 => "1111110001111100",
50276 => "1111110001111100",
50277 => "1111110001111100",
50278 => "1111110001111100",
50279 => "1111110001111101",
50280 => "1111110001111101",
50281 => "1111110001111101",
50282 => "1111110001111101",
50283 => "1111110001111101",
50284 => "1111110001111110",
50285 => "1111110001111110",
50286 => "1111110001111110",
50287 => "1111110001111110",
50288 => "1111110001111111",
50289 => "1111110001111111",
50290 => "1111110001111111",
50291 => "1111110001111111",
50292 => "1111110001111111",
50293 => "1111110010000000",
50294 => "1111110010000000",
50295 => "1111110010000000",
50296 => "1111110010000000",
50297 => "1111110010000000",
50298 => "1111110010000001",
50299 => "1111110010000001",
50300 => "1111110010000001",
50301 => "1111110010000001",
50302 => "1111110010000010",
50303 => "1111110010000010",
50304 => "1111110010000010",
50305 => "1111110010000010",
50306 => "1111110010000010",
50307 => "1111110010000011",
50308 => "1111110010000011",
50309 => "1111110010000011",
50310 => "1111110010000011",
50311 => "1111110010000011",
50312 => "1111110010000100",
50313 => "1111110010000100",
50314 => "1111110010000100",
50315 => "1111110010000100",
50316 => "1111110010000101",
50317 => "1111110010000101",
50318 => "1111110010000101",
50319 => "1111110010000101",
50320 => "1111110010000101",
50321 => "1111110010000110",
50322 => "1111110010000110",
50323 => "1111110010000110",
50324 => "1111110010000110",
50325 => "1111110010000110",
50326 => "1111110010000111",
50327 => "1111110010000111",
50328 => "1111110010000111",
50329 => "1111110010000111",
50330 => "1111110010001000",
50331 => "1111110010001000",
50332 => "1111110010001000",
50333 => "1111110010001000",
50334 => "1111110010001000",
50335 => "1111110010001001",
50336 => "1111110010001001",
50337 => "1111110010001001",
50338 => "1111110010001001",
50339 => "1111110010001001",
50340 => "1111110010001010",
50341 => "1111110010001010",
50342 => "1111110010001010",
50343 => "1111110010001010",
50344 => "1111110010001011",
50345 => "1111110010001011",
50346 => "1111110010001011",
50347 => "1111110010001011",
50348 => "1111110010001011",
50349 => "1111110010001100",
50350 => "1111110010001100",
50351 => "1111110010001100",
50352 => "1111110010001100",
50353 => "1111110010001100",
50354 => "1111110010001101",
50355 => "1111110010001101",
50356 => "1111110010001101",
50357 => "1111110010001101",
50358 => "1111110010001110",
50359 => "1111110010001110",
50360 => "1111110010001110",
50361 => "1111110010001110",
50362 => "1111110010001110",
50363 => "1111110010001111",
50364 => "1111110010001111",
50365 => "1111110010001111",
50366 => "1111110010001111",
50367 => "1111110010001111",
50368 => "1111110010010000",
50369 => "1111110010010000",
50370 => "1111110010010000",
50371 => "1111110010010000",
50372 => "1111110010010000",
50373 => "1111110010010001",
50374 => "1111110010010001",
50375 => "1111110010010001",
50376 => "1111110010010001",
50377 => "1111110010010010",
50378 => "1111110010010010",
50379 => "1111110010010010",
50380 => "1111110010010010",
50381 => "1111110010010010",
50382 => "1111110010010011",
50383 => "1111110010010011",
50384 => "1111110010010011",
50385 => "1111110010010011",
50386 => "1111110010010011",
50387 => "1111110010010100",
50388 => "1111110010010100",
50389 => "1111110010010100",
50390 => "1111110010010100",
50391 => "1111110010010100",
50392 => "1111110010010101",
50393 => "1111110010010101",
50394 => "1111110010010101",
50395 => "1111110010010101",
50396 => "1111110010010110",
50397 => "1111110010010110",
50398 => "1111110010010110",
50399 => "1111110010010110",
50400 => "1111110010010110",
50401 => "1111110010010111",
50402 => "1111110010010111",
50403 => "1111110010010111",
50404 => "1111110010010111",
50405 => "1111110010010111",
50406 => "1111110010011000",
50407 => "1111110010011000",
50408 => "1111110010011000",
50409 => "1111110010011000",
50410 => "1111110010011000",
50411 => "1111110010011001",
50412 => "1111110010011001",
50413 => "1111110010011001",
50414 => "1111110010011001",
50415 => "1111110010011010",
50416 => "1111110010011010",
50417 => "1111110010011010",
50418 => "1111110010011010",
50419 => "1111110010011010",
50420 => "1111110010011011",
50421 => "1111110010011011",
50422 => "1111110010011011",
50423 => "1111110010011011",
50424 => "1111110010011011",
50425 => "1111110010011100",
50426 => "1111110010011100",
50427 => "1111110010011100",
50428 => "1111110010011100",
50429 => "1111110010011100",
50430 => "1111110010011101",
50431 => "1111110010011101",
50432 => "1111110010011101",
50433 => "1111110010011101",
50434 => "1111110010011110",
50435 => "1111110010011110",
50436 => "1111110010011110",
50437 => "1111110010011110",
50438 => "1111110010011110",
50439 => "1111110010011111",
50440 => "1111110010011111",
50441 => "1111110010011111",
50442 => "1111110010011111",
50443 => "1111110010011111",
50444 => "1111110010100000",
50445 => "1111110010100000",
50446 => "1111110010100000",
50447 => "1111110010100000",
50448 => "1111110010100000",
50449 => "1111110010100001",
50450 => "1111110010100001",
50451 => "1111110010100001",
50452 => "1111110010100001",
50453 => "1111110010100001",
50454 => "1111110010100010",
50455 => "1111110010100010",
50456 => "1111110010100010",
50457 => "1111110010100010",
50458 => "1111110010100011",
50459 => "1111110010100011",
50460 => "1111110010100011",
50461 => "1111110010100011",
50462 => "1111110010100011",
50463 => "1111110010100100",
50464 => "1111110010100100",
50465 => "1111110010100100",
50466 => "1111110010100100",
50467 => "1111110010100100",
50468 => "1111110010100101",
50469 => "1111110010100101",
50470 => "1111110010100101",
50471 => "1111110010100101",
50472 => "1111110010100101",
50473 => "1111110010100110",
50474 => "1111110010100110",
50475 => "1111110010100110",
50476 => "1111110010100110",
50477 => "1111110010100110",
50478 => "1111110010100111",
50479 => "1111110010100111",
50480 => "1111110010100111",
50481 => "1111110010100111",
50482 => "1111110010100111",
50483 => "1111110010101000",
50484 => "1111110010101000",
50485 => "1111110010101000",
50486 => "1111110010101000",
50487 => "1111110010101000",
50488 => "1111110010101001",
50489 => "1111110010101001",
50490 => "1111110010101001",
50491 => "1111110010101001",
50492 => "1111110010101010",
50493 => "1111110010101010",
50494 => "1111110010101010",
50495 => "1111110010101010",
50496 => "1111110010101010",
50497 => "1111110010101011",
50498 => "1111110010101011",
50499 => "1111110010101011",
50500 => "1111110010101011",
50501 => "1111110010101011",
50502 => "1111110010101100",
50503 => "1111110010101100",
50504 => "1111110010101100",
50505 => "1111110010101100",
50506 => "1111110010101100",
50507 => "1111110010101101",
50508 => "1111110010101101",
50509 => "1111110010101101",
50510 => "1111110010101101",
50511 => "1111110010101101",
50512 => "1111110010101110",
50513 => "1111110010101110",
50514 => "1111110010101110",
50515 => "1111110010101110",
50516 => "1111110010101110",
50517 => "1111110010101111",
50518 => "1111110010101111",
50519 => "1111110010101111",
50520 => "1111110010101111",
50521 => "1111110010101111",
50522 => "1111110010110000",
50523 => "1111110010110000",
50524 => "1111110010110000",
50525 => "1111110010110000",
50526 => "1111110010110000",
50527 => "1111110010110001",
50528 => "1111110010110001",
50529 => "1111110010110001",
50530 => "1111110010110001",
50531 => "1111110010110010",
50532 => "1111110010110010",
50533 => "1111110010110010",
50534 => "1111110010110010",
50535 => "1111110010110010",
50536 => "1111110010110011",
50537 => "1111110010110011",
50538 => "1111110010110011",
50539 => "1111110010110011",
50540 => "1111110010110011",
50541 => "1111110010110100",
50542 => "1111110010110100",
50543 => "1111110010110100",
50544 => "1111110010110100",
50545 => "1111110010110100",
50546 => "1111110010110101",
50547 => "1111110010110101",
50548 => "1111110010110101",
50549 => "1111110010110101",
50550 => "1111110010110101",
50551 => "1111110010110110",
50552 => "1111110010110110",
50553 => "1111110010110110",
50554 => "1111110010110110",
50555 => "1111110010110110",
50556 => "1111110010110111",
50557 => "1111110010110111",
50558 => "1111110010110111",
50559 => "1111110010110111",
50560 => "1111110010110111",
50561 => "1111110010111000",
50562 => "1111110010111000",
50563 => "1111110010111000",
50564 => "1111110010111000",
50565 => "1111110010111000",
50566 => "1111110010111001",
50567 => "1111110010111001",
50568 => "1111110010111001",
50569 => "1111110010111001",
50570 => "1111110010111001",
50571 => "1111110010111010",
50572 => "1111110010111010",
50573 => "1111110010111010",
50574 => "1111110010111010",
50575 => "1111110010111010",
50576 => "1111110010111011",
50577 => "1111110010111011",
50578 => "1111110010111011",
50579 => "1111110010111011",
50580 => "1111110010111011",
50581 => "1111110010111100",
50582 => "1111110010111100",
50583 => "1111110010111100",
50584 => "1111110010111100",
50585 => "1111110010111100",
50586 => "1111110010111101",
50587 => "1111110010111101",
50588 => "1111110010111101",
50589 => "1111110010111101",
50590 => "1111110010111101",
50591 => "1111110010111110",
50592 => "1111110010111110",
50593 => "1111110010111110",
50594 => "1111110010111110",
50595 => "1111110010111110",
50596 => "1111110010111111",
50597 => "1111110010111111",
50598 => "1111110010111111",
50599 => "1111110010111111",
50600 => "1111110010111111",
50601 => "1111110011000000",
50602 => "1111110011000000",
50603 => "1111110011000000",
50604 => "1111110011000000",
50605 => "1111110011000000",
50606 => "1111110011000001",
50607 => "1111110011000001",
50608 => "1111110011000001",
50609 => "1111110011000001",
50610 => "1111110011000001",
50611 => "1111110011000010",
50612 => "1111110011000010",
50613 => "1111110011000010",
50614 => "1111110011000010",
50615 => "1111110011000010",
50616 => "1111110011000011",
50617 => "1111110011000011",
50618 => "1111110011000011",
50619 => "1111110011000011",
50620 => "1111110011000011",
50621 => "1111110011000100",
50622 => "1111110011000100",
50623 => "1111110011000100",
50624 => "1111110011000100",
50625 => "1111110011000100",
50626 => "1111110011000101",
50627 => "1111110011000101",
50628 => "1111110011000101",
50629 => "1111110011000101",
50630 => "1111110011000101",
50631 => "1111110011000110",
50632 => "1111110011000110",
50633 => "1111110011000110",
50634 => "1111110011000110",
50635 => "1111110011000110",
50636 => "1111110011000111",
50637 => "1111110011000111",
50638 => "1111110011000111",
50639 => "1111110011000111",
50640 => "1111110011000111",
50641 => "1111110011001000",
50642 => "1111110011001000",
50643 => "1111110011001000",
50644 => "1111110011001000",
50645 => "1111110011001000",
50646 => "1111110011001001",
50647 => "1111110011001001",
50648 => "1111110011001001",
50649 => "1111110011001001",
50650 => "1111110011001001",
50651 => "1111110011001010",
50652 => "1111110011001010",
50653 => "1111110011001010",
50654 => "1111110011001010",
50655 => "1111110011001010",
50656 => "1111110011001011",
50657 => "1111110011001011",
50658 => "1111110011001011",
50659 => "1111110011001011",
50660 => "1111110011001011",
50661 => "1111110011001100",
50662 => "1111110011001100",
50663 => "1111110011001100",
50664 => "1111110011001100",
50665 => "1111110011001100",
50666 => "1111110011001101",
50667 => "1111110011001101",
50668 => "1111110011001101",
50669 => "1111110011001101",
50670 => "1111110011001101",
50671 => "1111110011001110",
50672 => "1111110011001110",
50673 => "1111110011001110",
50674 => "1111110011001110",
50675 => "1111110011001110",
50676 => "1111110011001111",
50677 => "1111110011001111",
50678 => "1111110011001111",
50679 => "1111110011001111",
50680 => "1111110011001111",
50681 => "1111110011010000",
50682 => "1111110011010000",
50683 => "1111110011010000",
50684 => "1111110011010000",
50685 => "1111110011010000",
50686 => "1111110011010001",
50687 => "1111110011010001",
50688 => "1111110011010001",
50689 => "1111110011010001",
50690 => "1111110011010001",
50691 => "1111110011010010",
50692 => "1111110011010010",
50693 => "1111110011010010",
50694 => "1111110011010010",
50695 => "1111110011010010",
50696 => "1111110011010011",
50697 => "1111110011010011",
50698 => "1111110011010011",
50699 => "1111110011010011",
50700 => "1111110011010011",
50701 => "1111110011010011",
50702 => "1111110011010100",
50703 => "1111110011010100",
50704 => "1111110011010100",
50705 => "1111110011010100",
50706 => "1111110011010100",
50707 => "1111110011010101",
50708 => "1111110011010101",
50709 => "1111110011010101",
50710 => "1111110011010101",
50711 => "1111110011010101",
50712 => "1111110011010110",
50713 => "1111110011010110",
50714 => "1111110011010110",
50715 => "1111110011010110",
50716 => "1111110011010110",
50717 => "1111110011010111",
50718 => "1111110011010111",
50719 => "1111110011010111",
50720 => "1111110011010111",
50721 => "1111110011010111",
50722 => "1111110011011000",
50723 => "1111110011011000",
50724 => "1111110011011000",
50725 => "1111110011011000",
50726 => "1111110011011000",
50727 => "1111110011011001",
50728 => "1111110011011001",
50729 => "1111110011011001",
50730 => "1111110011011001",
50731 => "1111110011011001",
50732 => "1111110011011010",
50733 => "1111110011011010",
50734 => "1111110011011010",
50735 => "1111110011011010",
50736 => "1111110011011010",
50737 => "1111110011011010",
50738 => "1111110011011011",
50739 => "1111110011011011",
50740 => "1111110011011011",
50741 => "1111110011011011",
50742 => "1111110011011011",
50743 => "1111110011011100",
50744 => "1111110011011100",
50745 => "1111110011011100",
50746 => "1111110011011100",
50747 => "1111110011011100",
50748 => "1111110011011101",
50749 => "1111110011011101",
50750 => "1111110011011101",
50751 => "1111110011011101",
50752 => "1111110011011101",
50753 => "1111110011011110",
50754 => "1111110011011110",
50755 => "1111110011011110",
50756 => "1111110011011110",
50757 => "1111110011011110",
50758 => "1111110011011111",
50759 => "1111110011011111",
50760 => "1111110011011111",
50761 => "1111110011011111",
50762 => "1111110011011111",
50763 => "1111110011100000",
50764 => "1111110011100000",
50765 => "1111110011100000",
50766 => "1111110011100000",
50767 => "1111110011100000",
50768 => "1111110011100000",
50769 => "1111110011100001",
50770 => "1111110011100001",
50771 => "1111110011100001",
50772 => "1111110011100001",
50773 => "1111110011100001",
50774 => "1111110011100010",
50775 => "1111110011100010",
50776 => "1111110011100010",
50777 => "1111110011100010",
50778 => "1111110011100010",
50779 => "1111110011100011",
50780 => "1111110011100011",
50781 => "1111110011100011",
50782 => "1111110011100011",
50783 => "1111110011100011",
50784 => "1111110011100100",
50785 => "1111110011100100",
50786 => "1111110011100100",
50787 => "1111110011100100",
50788 => "1111110011100100",
50789 => "1111110011100101",
50790 => "1111110011100101",
50791 => "1111110011100101",
50792 => "1111110011100101",
50793 => "1111110011100101",
50794 => "1111110011100101",
50795 => "1111110011100110",
50796 => "1111110011100110",
50797 => "1111110011100110",
50798 => "1111110011100110",
50799 => "1111110011100110",
50800 => "1111110011100111",
50801 => "1111110011100111",
50802 => "1111110011100111",
50803 => "1111110011100111",
50804 => "1111110011100111",
50805 => "1111110011101000",
50806 => "1111110011101000",
50807 => "1111110011101000",
50808 => "1111110011101000",
50809 => "1111110011101000",
50810 => "1111110011101001",
50811 => "1111110011101001",
50812 => "1111110011101001",
50813 => "1111110011101001",
50814 => "1111110011101001",
50815 => "1111110011101010",
50816 => "1111110011101010",
50817 => "1111110011101010",
50818 => "1111110011101010",
50819 => "1111110011101010",
50820 => "1111110011101010",
50821 => "1111110011101011",
50822 => "1111110011101011",
50823 => "1111110011101011",
50824 => "1111110011101011",
50825 => "1111110011101011",
50826 => "1111110011101100",
50827 => "1111110011101100",
50828 => "1111110011101100",
50829 => "1111110011101100",
50830 => "1111110011101100",
50831 => "1111110011101101",
50832 => "1111110011101101",
50833 => "1111110011101101",
50834 => "1111110011101101",
50835 => "1111110011101101",
50836 => "1111110011101101",
50837 => "1111110011101110",
50838 => "1111110011101110",
50839 => "1111110011101110",
50840 => "1111110011101110",
50841 => "1111110011101110",
50842 => "1111110011101111",
50843 => "1111110011101111",
50844 => "1111110011101111",
50845 => "1111110011101111",
50846 => "1111110011101111",
50847 => "1111110011110000",
50848 => "1111110011110000",
50849 => "1111110011110000",
50850 => "1111110011110000",
50851 => "1111110011110000",
50852 => "1111110011110001",
50853 => "1111110011110001",
50854 => "1111110011110001",
50855 => "1111110011110001",
50856 => "1111110011110001",
50857 => "1111110011110001",
50858 => "1111110011110010",
50859 => "1111110011110010",
50860 => "1111110011110010",
50861 => "1111110011110010",
50862 => "1111110011110010",
50863 => "1111110011110011",
50864 => "1111110011110011",
50865 => "1111110011110011",
50866 => "1111110011110011",
50867 => "1111110011110011",
50868 => "1111110011110100",
50869 => "1111110011110100",
50870 => "1111110011110100",
50871 => "1111110011110100",
50872 => "1111110011110100",
50873 => "1111110011110100",
50874 => "1111110011110101",
50875 => "1111110011110101",
50876 => "1111110011110101",
50877 => "1111110011110101",
50878 => "1111110011110101",
50879 => "1111110011110110",
50880 => "1111110011110110",
50881 => "1111110011110110",
50882 => "1111110011110110",
50883 => "1111110011110110",
50884 => "1111110011110111",
50885 => "1111110011110111",
50886 => "1111110011110111",
50887 => "1111110011110111",
50888 => "1111110011110111",
50889 => "1111110011110111",
50890 => "1111110011111000",
50891 => "1111110011111000",
50892 => "1111110011111000",
50893 => "1111110011111000",
50894 => "1111110011111000",
50895 => "1111110011111001",
50896 => "1111110011111001",
50897 => "1111110011111001",
50898 => "1111110011111001",
50899 => "1111110011111001",
50900 => "1111110011111010",
50901 => "1111110011111010",
50902 => "1111110011111010",
50903 => "1111110011111010",
50904 => "1111110011111010",
50905 => "1111110011111010",
50906 => "1111110011111011",
50907 => "1111110011111011",
50908 => "1111110011111011",
50909 => "1111110011111011",
50910 => "1111110011111011",
50911 => "1111110011111100",
50912 => "1111110011111100",
50913 => "1111110011111100",
50914 => "1111110011111100",
50915 => "1111110011111100",
50916 => "1111110011111101",
50917 => "1111110011111101",
50918 => "1111110011111101",
50919 => "1111110011111101",
50920 => "1111110011111101",
50921 => "1111110011111101",
50922 => "1111110011111110",
50923 => "1111110011111110",
50924 => "1111110011111110",
50925 => "1111110011111110",
50926 => "1111110011111110",
50927 => "1111110011111111",
50928 => "1111110011111111",
50929 => "1111110011111111",
50930 => "1111110011111111",
50931 => "1111110011111111",
50932 => "1111110011111111",
50933 => "1111110100000000",
50934 => "1111110100000000",
50935 => "1111110100000000",
50936 => "1111110100000000",
50937 => "1111110100000000",
50938 => "1111110100000001",
50939 => "1111110100000001",
50940 => "1111110100000001",
50941 => "1111110100000001",
50942 => "1111110100000001",
50943 => "1111110100000010",
50944 => "1111110100000010",
50945 => "1111110100000010",
50946 => "1111110100000010",
50947 => "1111110100000010",
50948 => "1111110100000010",
50949 => "1111110100000011",
50950 => "1111110100000011",
50951 => "1111110100000011",
50952 => "1111110100000011",
50953 => "1111110100000011",
50954 => "1111110100000100",
50955 => "1111110100000100",
50956 => "1111110100000100",
50957 => "1111110100000100",
50958 => "1111110100000100",
50959 => "1111110100000100",
50960 => "1111110100000101",
50961 => "1111110100000101",
50962 => "1111110100000101",
50963 => "1111110100000101",
50964 => "1111110100000101",
50965 => "1111110100000110",
50966 => "1111110100000110",
50967 => "1111110100000110",
50968 => "1111110100000110",
50969 => "1111110100000110",
50970 => "1111110100000110",
50971 => "1111110100000111",
50972 => "1111110100000111",
50973 => "1111110100000111",
50974 => "1111110100000111",
50975 => "1111110100000111",
50976 => "1111110100001000",
50977 => "1111110100001000",
50978 => "1111110100001000",
50979 => "1111110100001000",
50980 => "1111110100001000",
50981 => "1111110100001001",
50982 => "1111110100001001",
50983 => "1111110100001001",
50984 => "1111110100001001",
50985 => "1111110100001001",
50986 => "1111110100001001",
50987 => "1111110100001010",
50988 => "1111110100001010",
50989 => "1111110100001010",
50990 => "1111110100001010",
50991 => "1111110100001010",
50992 => "1111110100001011",
50993 => "1111110100001011",
50994 => "1111110100001011",
50995 => "1111110100001011",
50996 => "1111110100001011",
50997 => "1111110100001011",
50998 => "1111110100001100",
50999 => "1111110100001100",
51000 => "1111110100001100",
51001 => "1111110100001100",
51002 => "1111110100001100",
51003 => "1111110100001101",
51004 => "1111110100001101",
51005 => "1111110100001101",
51006 => "1111110100001101",
51007 => "1111110100001101",
51008 => "1111110100001101",
51009 => "1111110100001110",
51010 => "1111110100001110",
51011 => "1111110100001110",
51012 => "1111110100001110",
51013 => "1111110100001110",
51014 => "1111110100001111",
51015 => "1111110100001111",
51016 => "1111110100001111",
51017 => "1111110100001111",
51018 => "1111110100001111",
51019 => "1111110100001111",
51020 => "1111110100010000",
51021 => "1111110100010000",
51022 => "1111110100010000",
51023 => "1111110100010000",
51024 => "1111110100010000",
51025 => "1111110100010001",
51026 => "1111110100010001",
51027 => "1111110100010001",
51028 => "1111110100010001",
51029 => "1111110100010001",
51030 => "1111110100010001",
51031 => "1111110100010010",
51032 => "1111110100010010",
51033 => "1111110100010010",
51034 => "1111110100010010",
51035 => "1111110100010010",
51036 => "1111110100010011",
51037 => "1111110100010011",
51038 => "1111110100010011",
51039 => "1111110100010011",
51040 => "1111110100010011",
51041 => "1111110100010011",
51042 => "1111110100010100",
51043 => "1111110100010100",
51044 => "1111110100010100",
51045 => "1111110100010100",
51046 => "1111110100010100",
51047 => "1111110100010101",
51048 => "1111110100010101",
51049 => "1111110100010101",
51050 => "1111110100010101",
51051 => "1111110100010101",
51052 => "1111110100010101",
51053 => "1111110100010110",
51054 => "1111110100010110",
51055 => "1111110100010110",
51056 => "1111110100010110",
51057 => "1111110100010110",
51058 => "1111110100010110",
51059 => "1111110100010111",
51060 => "1111110100010111",
51061 => "1111110100010111",
51062 => "1111110100010111",
51063 => "1111110100010111",
51064 => "1111110100011000",
51065 => "1111110100011000",
51066 => "1111110100011000",
51067 => "1111110100011000",
51068 => "1111110100011000",
51069 => "1111110100011000",
51070 => "1111110100011001",
51071 => "1111110100011001",
51072 => "1111110100011001",
51073 => "1111110100011001",
51074 => "1111110100011001",
51075 => "1111110100011010",
51076 => "1111110100011010",
51077 => "1111110100011010",
51078 => "1111110100011010",
51079 => "1111110100011010",
51080 => "1111110100011010",
51081 => "1111110100011011",
51082 => "1111110100011011",
51083 => "1111110100011011",
51084 => "1111110100011011",
51085 => "1111110100011011",
51086 => "1111110100011100",
51087 => "1111110100011100",
51088 => "1111110100011100",
51089 => "1111110100011100",
51090 => "1111110100011100",
51091 => "1111110100011100",
51092 => "1111110100011101",
51093 => "1111110100011101",
51094 => "1111110100011101",
51095 => "1111110100011101",
51096 => "1111110100011101",
51097 => "1111110100011101",
51098 => "1111110100011110",
51099 => "1111110100011110",
51100 => "1111110100011110",
51101 => "1111110100011110",
51102 => "1111110100011110",
51103 => "1111110100011111",
51104 => "1111110100011111",
51105 => "1111110100011111",
51106 => "1111110100011111",
51107 => "1111110100011111",
51108 => "1111110100011111",
51109 => "1111110100100000",
51110 => "1111110100100000",
51111 => "1111110100100000",
51112 => "1111110100100000",
51113 => "1111110100100000",
51114 => "1111110100100000",
51115 => "1111110100100001",
51116 => "1111110100100001",
51117 => "1111110100100001",
51118 => "1111110100100001",
51119 => "1111110100100001",
51120 => "1111110100100010",
51121 => "1111110100100010",
51122 => "1111110100100010",
51123 => "1111110100100010",
51124 => "1111110100100010",
51125 => "1111110100100010",
51126 => "1111110100100011",
51127 => "1111110100100011",
51128 => "1111110100100011",
51129 => "1111110100100011",
51130 => "1111110100100011",
51131 => "1111110100100100",
51132 => "1111110100100100",
51133 => "1111110100100100",
51134 => "1111110100100100",
51135 => "1111110100100100",
51136 => "1111110100100100",
51137 => "1111110100100101",
51138 => "1111110100100101",
51139 => "1111110100100101",
51140 => "1111110100100101",
51141 => "1111110100100101",
51142 => "1111110100100101",
51143 => "1111110100100110",
51144 => "1111110100100110",
51145 => "1111110100100110",
51146 => "1111110100100110",
51147 => "1111110100100110",
51148 => "1111110100100111",
51149 => "1111110100100111",
51150 => "1111110100100111",
51151 => "1111110100100111",
51152 => "1111110100100111",
51153 => "1111110100100111",
51154 => "1111110100101000",
51155 => "1111110100101000",
51156 => "1111110100101000",
51157 => "1111110100101000",
51158 => "1111110100101000",
51159 => "1111110100101000",
51160 => "1111110100101001",
51161 => "1111110100101001",
51162 => "1111110100101001",
51163 => "1111110100101001",
51164 => "1111110100101001",
51165 => "1111110100101001",
51166 => "1111110100101010",
51167 => "1111110100101010",
51168 => "1111110100101010",
51169 => "1111110100101010",
51170 => "1111110100101010",
51171 => "1111110100101011",
51172 => "1111110100101011",
51173 => "1111110100101011",
51174 => "1111110100101011",
51175 => "1111110100101011",
51176 => "1111110100101011",
51177 => "1111110100101100",
51178 => "1111110100101100",
51179 => "1111110100101100",
51180 => "1111110100101100",
51181 => "1111110100101100",
51182 => "1111110100101100",
51183 => "1111110100101101",
51184 => "1111110100101101",
51185 => "1111110100101101",
51186 => "1111110100101101",
51187 => "1111110100101101",
51188 => "1111110100101110",
51189 => "1111110100101110",
51190 => "1111110100101110",
51191 => "1111110100101110",
51192 => "1111110100101110",
51193 => "1111110100101110",
51194 => "1111110100101111",
51195 => "1111110100101111",
51196 => "1111110100101111",
51197 => "1111110100101111",
51198 => "1111110100101111",
51199 => "1111110100101111",
51200 => "1111110100110000",
51201 => "1111110100110000",
51202 => "1111110100110000",
51203 => "1111110100110000",
51204 => "1111110100110000",
51205 => "1111110100110000",
51206 => "1111110100110001",
51207 => "1111110100110001",
51208 => "1111110100110001",
51209 => "1111110100110001",
51210 => "1111110100110001",
51211 => "1111110100110010",
51212 => "1111110100110010",
51213 => "1111110100110010",
51214 => "1111110100110010",
51215 => "1111110100110010",
51216 => "1111110100110010",
51217 => "1111110100110011",
51218 => "1111110100110011",
51219 => "1111110100110011",
51220 => "1111110100110011",
51221 => "1111110100110011",
51222 => "1111110100110011",
51223 => "1111110100110100",
51224 => "1111110100110100",
51225 => "1111110100110100",
51226 => "1111110100110100",
51227 => "1111110100110100",
51228 => "1111110100110100",
51229 => "1111110100110101",
51230 => "1111110100110101",
51231 => "1111110100110101",
51232 => "1111110100110101",
51233 => "1111110100110101",
51234 => "1111110100110101",
51235 => "1111110100110110",
51236 => "1111110100110110",
51237 => "1111110100110110",
51238 => "1111110100110110",
51239 => "1111110100110110",
51240 => "1111110100110111",
51241 => "1111110100110111",
51242 => "1111110100110111",
51243 => "1111110100110111",
51244 => "1111110100110111",
51245 => "1111110100110111",
51246 => "1111110100111000",
51247 => "1111110100111000",
51248 => "1111110100111000",
51249 => "1111110100111000",
51250 => "1111110100111000",
51251 => "1111110100111000",
51252 => "1111110100111001",
51253 => "1111110100111001",
51254 => "1111110100111001",
51255 => "1111110100111001",
51256 => "1111110100111001",
51257 => "1111110100111001",
51258 => "1111110100111010",
51259 => "1111110100111010",
51260 => "1111110100111010",
51261 => "1111110100111010",
51262 => "1111110100111010",
51263 => "1111110100111010",
51264 => "1111110100111011",
51265 => "1111110100111011",
51266 => "1111110100111011",
51267 => "1111110100111011",
51268 => "1111110100111011",
51269 => "1111110100111011",
51270 => "1111110100111100",
51271 => "1111110100111100",
51272 => "1111110100111100",
51273 => "1111110100111100",
51274 => "1111110100111100",
51275 => "1111110100111101",
51276 => "1111110100111101",
51277 => "1111110100111101",
51278 => "1111110100111101",
51279 => "1111110100111101",
51280 => "1111110100111101",
51281 => "1111110100111110",
51282 => "1111110100111110",
51283 => "1111110100111110",
51284 => "1111110100111110",
51285 => "1111110100111110",
51286 => "1111110100111110",
51287 => "1111110100111111",
51288 => "1111110100111111",
51289 => "1111110100111111",
51290 => "1111110100111111",
51291 => "1111110100111111",
51292 => "1111110100111111",
51293 => "1111110101000000",
51294 => "1111110101000000",
51295 => "1111110101000000",
51296 => "1111110101000000",
51297 => "1111110101000000",
51298 => "1111110101000000",
51299 => "1111110101000001",
51300 => "1111110101000001",
51301 => "1111110101000001",
51302 => "1111110101000001",
51303 => "1111110101000001",
51304 => "1111110101000001",
51305 => "1111110101000010",
51306 => "1111110101000010",
51307 => "1111110101000010",
51308 => "1111110101000010",
51309 => "1111110101000010",
51310 => "1111110101000010",
51311 => "1111110101000011",
51312 => "1111110101000011",
51313 => "1111110101000011",
51314 => "1111110101000011",
51315 => "1111110101000011",
51316 => "1111110101000011",
51317 => "1111110101000100",
51318 => "1111110101000100",
51319 => "1111110101000100",
51320 => "1111110101000100",
51321 => "1111110101000100",
51322 => "1111110101000100",
51323 => "1111110101000101",
51324 => "1111110101000101",
51325 => "1111110101000101",
51326 => "1111110101000101",
51327 => "1111110101000101",
51328 => "1111110101000110",
51329 => "1111110101000110",
51330 => "1111110101000110",
51331 => "1111110101000110",
51332 => "1111110101000110",
51333 => "1111110101000110",
51334 => "1111110101000111",
51335 => "1111110101000111",
51336 => "1111110101000111",
51337 => "1111110101000111",
51338 => "1111110101000111",
51339 => "1111110101000111",
51340 => "1111110101001000",
51341 => "1111110101001000",
51342 => "1111110101001000",
51343 => "1111110101001000",
51344 => "1111110101001000",
51345 => "1111110101001000",
51346 => "1111110101001001",
51347 => "1111110101001001",
51348 => "1111110101001001",
51349 => "1111110101001001",
51350 => "1111110101001001",
51351 => "1111110101001001",
51352 => "1111110101001010",
51353 => "1111110101001010",
51354 => "1111110101001010",
51355 => "1111110101001010",
51356 => "1111110101001010",
51357 => "1111110101001010",
51358 => "1111110101001011",
51359 => "1111110101001011",
51360 => "1111110101001011",
51361 => "1111110101001011",
51362 => "1111110101001011",
51363 => "1111110101001011",
51364 => "1111110101001100",
51365 => "1111110101001100",
51366 => "1111110101001100",
51367 => "1111110101001100",
51368 => "1111110101001100",
51369 => "1111110101001100",
51370 => "1111110101001101",
51371 => "1111110101001101",
51372 => "1111110101001101",
51373 => "1111110101001101",
51374 => "1111110101001101",
51375 => "1111110101001101",
51376 => "1111110101001110",
51377 => "1111110101001110",
51378 => "1111110101001110",
51379 => "1111110101001110",
51380 => "1111110101001110",
51381 => "1111110101001110",
51382 => "1111110101001111",
51383 => "1111110101001111",
51384 => "1111110101001111",
51385 => "1111110101001111",
51386 => "1111110101001111",
51387 => "1111110101001111",
51388 => "1111110101010000",
51389 => "1111110101010000",
51390 => "1111110101010000",
51391 => "1111110101010000",
51392 => "1111110101010000",
51393 => "1111110101010000",
51394 => "1111110101010001",
51395 => "1111110101010001",
51396 => "1111110101010001",
51397 => "1111110101010001",
51398 => "1111110101010001",
51399 => "1111110101010001",
51400 => "1111110101010010",
51401 => "1111110101010010",
51402 => "1111110101010010",
51403 => "1111110101010010",
51404 => "1111110101010010",
51405 => "1111110101010010",
51406 => "1111110101010011",
51407 => "1111110101010011",
51408 => "1111110101010011",
51409 => "1111110101010011",
51410 => "1111110101010011",
51411 => "1111110101010011",
51412 => "1111110101010100",
51413 => "1111110101010100",
51414 => "1111110101010100",
51415 => "1111110101010100",
51416 => "1111110101010100",
51417 => "1111110101010100",
51418 => "1111110101010101",
51419 => "1111110101010101",
51420 => "1111110101010101",
51421 => "1111110101010101",
51422 => "1111110101010101",
51423 => "1111110101010101",
51424 => "1111110101010110",
51425 => "1111110101010110",
51426 => "1111110101010110",
51427 => "1111110101010110",
51428 => "1111110101010110",
51429 => "1111110101010110",
51430 => "1111110101010110",
51431 => "1111110101010111",
51432 => "1111110101010111",
51433 => "1111110101010111",
51434 => "1111110101010111",
51435 => "1111110101010111",
51436 => "1111110101010111",
51437 => "1111110101011000",
51438 => "1111110101011000",
51439 => "1111110101011000",
51440 => "1111110101011000",
51441 => "1111110101011000",
51442 => "1111110101011000",
51443 => "1111110101011001",
51444 => "1111110101011001",
51445 => "1111110101011001",
51446 => "1111110101011001",
51447 => "1111110101011001",
51448 => "1111110101011001",
51449 => "1111110101011010",
51450 => "1111110101011010",
51451 => "1111110101011010",
51452 => "1111110101011010",
51453 => "1111110101011010",
51454 => "1111110101011010",
51455 => "1111110101011011",
51456 => "1111110101011011",
51457 => "1111110101011011",
51458 => "1111110101011011",
51459 => "1111110101011011",
51460 => "1111110101011011",
51461 => "1111110101011100",
51462 => "1111110101011100",
51463 => "1111110101011100",
51464 => "1111110101011100",
51465 => "1111110101011100",
51466 => "1111110101011100",
51467 => "1111110101011101",
51468 => "1111110101011101",
51469 => "1111110101011101",
51470 => "1111110101011101",
51471 => "1111110101011101",
51472 => "1111110101011101",
51473 => "1111110101011110",
51474 => "1111110101011110",
51475 => "1111110101011110",
51476 => "1111110101011110",
51477 => "1111110101011110",
51478 => "1111110101011110",
51479 => "1111110101011111",
51480 => "1111110101011111",
51481 => "1111110101011111",
51482 => "1111110101011111",
51483 => "1111110101011111",
51484 => "1111110101011111",
51485 => "1111110101011111",
51486 => "1111110101100000",
51487 => "1111110101100000",
51488 => "1111110101100000",
51489 => "1111110101100000",
51490 => "1111110101100000",
51491 => "1111110101100000",
51492 => "1111110101100001",
51493 => "1111110101100001",
51494 => "1111110101100001",
51495 => "1111110101100001",
51496 => "1111110101100001",
51497 => "1111110101100001",
51498 => "1111110101100010",
51499 => "1111110101100010",
51500 => "1111110101100010",
51501 => "1111110101100010",
51502 => "1111110101100010",
51503 => "1111110101100010",
51504 => "1111110101100011",
51505 => "1111110101100011",
51506 => "1111110101100011",
51507 => "1111110101100011",
51508 => "1111110101100011",
51509 => "1111110101100011",
51510 => "1111110101100100",
51511 => "1111110101100100",
51512 => "1111110101100100",
51513 => "1111110101100100",
51514 => "1111110101100100",
51515 => "1111110101100100",
51516 => "1111110101100101",
51517 => "1111110101100101",
51518 => "1111110101100101",
51519 => "1111110101100101",
51520 => "1111110101100101",
51521 => "1111110101100101",
51522 => "1111110101100101",
51523 => "1111110101100110",
51524 => "1111110101100110",
51525 => "1111110101100110",
51526 => "1111110101100110",
51527 => "1111110101100110",
51528 => "1111110101100110",
51529 => "1111110101100111",
51530 => "1111110101100111",
51531 => "1111110101100111",
51532 => "1111110101100111",
51533 => "1111110101100111",
51534 => "1111110101100111",
51535 => "1111110101101000",
51536 => "1111110101101000",
51537 => "1111110101101000",
51538 => "1111110101101000",
51539 => "1111110101101000",
51540 => "1111110101101000",
51541 => "1111110101101001",
51542 => "1111110101101001",
51543 => "1111110101101001",
51544 => "1111110101101001",
51545 => "1111110101101001",
51546 => "1111110101101001",
51547 => "1111110101101001",
51548 => "1111110101101010",
51549 => "1111110101101010",
51550 => "1111110101101010",
51551 => "1111110101101010",
51552 => "1111110101101010",
51553 => "1111110101101010",
51554 => "1111110101101011",
51555 => "1111110101101011",
51556 => "1111110101101011",
51557 => "1111110101101011",
51558 => "1111110101101011",
51559 => "1111110101101011",
51560 => "1111110101101100",
51561 => "1111110101101100",
51562 => "1111110101101100",
51563 => "1111110101101100",
51564 => "1111110101101100",
51565 => "1111110101101100",
51566 => "1111110101101101",
51567 => "1111110101101101",
51568 => "1111110101101101",
51569 => "1111110101101101",
51570 => "1111110101101101",
51571 => "1111110101101101",
51572 => "1111110101101101",
51573 => "1111110101101110",
51574 => "1111110101101110",
51575 => "1111110101101110",
51576 => "1111110101101110",
51577 => "1111110101101110",
51578 => "1111110101101110",
51579 => "1111110101101111",
51580 => "1111110101101111",
51581 => "1111110101101111",
51582 => "1111110101101111",
51583 => "1111110101101111",
51584 => "1111110101101111",
51585 => "1111110101110000",
51586 => "1111110101110000",
51587 => "1111110101110000",
51588 => "1111110101110000",
51589 => "1111110101110000",
51590 => "1111110101110000",
51591 => "1111110101110000",
51592 => "1111110101110001",
51593 => "1111110101110001",
51594 => "1111110101110001",
51595 => "1111110101110001",
51596 => "1111110101110001",
51597 => "1111110101110001",
51598 => "1111110101110010",
51599 => "1111110101110010",
51600 => "1111110101110010",
51601 => "1111110101110010",
51602 => "1111110101110010",
51603 => "1111110101110010",
51604 => "1111110101110011",
51605 => "1111110101110011",
51606 => "1111110101110011",
51607 => "1111110101110011",
51608 => "1111110101110011",
51609 => "1111110101110011",
51610 => "1111110101110011",
51611 => "1111110101110100",
51612 => "1111110101110100",
51613 => "1111110101110100",
51614 => "1111110101110100",
51615 => "1111110101110100",
51616 => "1111110101110100",
51617 => "1111110101110101",
51618 => "1111110101110101",
51619 => "1111110101110101",
51620 => "1111110101110101",
51621 => "1111110101110101",
51622 => "1111110101110101",
51623 => "1111110101110110",
51624 => "1111110101110110",
51625 => "1111110101110110",
51626 => "1111110101110110",
51627 => "1111110101110110",
51628 => "1111110101110110",
51629 => "1111110101110110",
51630 => "1111110101110111",
51631 => "1111110101110111",
51632 => "1111110101110111",
51633 => "1111110101110111",
51634 => "1111110101110111",
51635 => "1111110101110111",
51636 => "1111110101111000",
51637 => "1111110101111000",
51638 => "1111110101111000",
51639 => "1111110101111000",
51640 => "1111110101111000",
51641 => "1111110101111000",
51642 => "1111110101111001",
51643 => "1111110101111001",
51644 => "1111110101111001",
51645 => "1111110101111001",
51646 => "1111110101111001",
51647 => "1111110101111001",
51648 => "1111110101111001",
51649 => "1111110101111010",
51650 => "1111110101111010",
51651 => "1111110101111010",
51652 => "1111110101111010",
51653 => "1111110101111010",
51654 => "1111110101111010",
51655 => "1111110101111011",
51656 => "1111110101111011",
51657 => "1111110101111011",
51658 => "1111110101111011",
51659 => "1111110101111011",
51660 => "1111110101111011",
51661 => "1111110101111011",
51662 => "1111110101111100",
51663 => "1111110101111100",
51664 => "1111110101111100",
51665 => "1111110101111100",
51666 => "1111110101111100",
51667 => "1111110101111100",
51668 => "1111110101111101",
51669 => "1111110101111101",
51670 => "1111110101111101",
51671 => "1111110101111101",
51672 => "1111110101111101",
51673 => "1111110101111101",
51674 => "1111110101111101",
51675 => "1111110101111110",
51676 => "1111110101111110",
51677 => "1111110101111110",
51678 => "1111110101111110",
51679 => "1111110101111110",
51680 => "1111110101111110",
51681 => "1111110101111111",
51682 => "1111110101111111",
51683 => "1111110101111111",
51684 => "1111110101111111",
51685 => "1111110101111111",
51686 => "1111110101111111",
51687 => "1111110110000000",
51688 => "1111110110000000",
51689 => "1111110110000000",
51690 => "1111110110000000",
51691 => "1111110110000000",
51692 => "1111110110000000",
51693 => "1111110110000000",
51694 => "1111110110000001",
51695 => "1111110110000001",
51696 => "1111110110000001",
51697 => "1111110110000001",
51698 => "1111110110000001",
51699 => "1111110110000001",
51700 => "1111110110000010",
51701 => "1111110110000010",
51702 => "1111110110000010",
51703 => "1111110110000010",
51704 => "1111110110000010",
51705 => "1111110110000010",
51706 => "1111110110000010",
51707 => "1111110110000011",
51708 => "1111110110000011",
51709 => "1111110110000011",
51710 => "1111110110000011",
51711 => "1111110110000011",
51712 => "1111110110000011",
51713 => "1111110110000100",
51714 => "1111110110000100",
51715 => "1111110110000100",
51716 => "1111110110000100",
51717 => "1111110110000100",
51718 => "1111110110000100",
51719 => "1111110110000100",
51720 => "1111110110000101",
51721 => "1111110110000101",
51722 => "1111110110000101",
51723 => "1111110110000101",
51724 => "1111110110000101",
51725 => "1111110110000101",
51726 => "1111110110000110",
51727 => "1111110110000110",
51728 => "1111110110000110",
51729 => "1111110110000110",
51730 => "1111110110000110",
51731 => "1111110110000110",
51732 => "1111110110000110",
51733 => "1111110110000111",
51734 => "1111110110000111",
51735 => "1111110110000111",
51736 => "1111110110000111",
51737 => "1111110110000111",
51738 => "1111110110000111",
51739 => "1111110110001000",
51740 => "1111110110001000",
51741 => "1111110110001000",
51742 => "1111110110001000",
51743 => "1111110110001000",
51744 => "1111110110001000",
51745 => "1111110110001000",
51746 => "1111110110001001",
51747 => "1111110110001001",
51748 => "1111110110001001",
51749 => "1111110110001001",
51750 => "1111110110001001",
51751 => "1111110110001001",
51752 => "1111110110001001",
51753 => "1111110110001010",
51754 => "1111110110001010",
51755 => "1111110110001010",
51756 => "1111110110001010",
51757 => "1111110110001010",
51758 => "1111110110001010",
51759 => "1111110110001011",
51760 => "1111110110001011",
51761 => "1111110110001011",
51762 => "1111110110001011",
51763 => "1111110110001011",
51764 => "1111110110001011",
51765 => "1111110110001011",
51766 => "1111110110001100",
51767 => "1111110110001100",
51768 => "1111110110001100",
51769 => "1111110110001100",
51770 => "1111110110001100",
51771 => "1111110110001100",
51772 => "1111110110001101",
51773 => "1111110110001101",
51774 => "1111110110001101",
51775 => "1111110110001101",
51776 => "1111110110001101",
51777 => "1111110110001101",
51778 => "1111110110001101",
51779 => "1111110110001110",
51780 => "1111110110001110",
51781 => "1111110110001110",
51782 => "1111110110001110",
51783 => "1111110110001110",
51784 => "1111110110001110",
51785 => "1111110110001110",
51786 => "1111110110001111",
51787 => "1111110110001111",
51788 => "1111110110001111",
51789 => "1111110110001111",
51790 => "1111110110001111",
51791 => "1111110110001111",
51792 => "1111110110010000",
51793 => "1111110110010000",
51794 => "1111110110010000",
51795 => "1111110110010000",
51796 => "1111110110010000",
51797 => "1111110110010000",
51798 => "1111110110010000",
51799 => "1111110110010001",
51800 => "1111110110010001",
51801 => "1111110110010001",
51802 => "1111110110010001",
51803 => "1111110110010001",
51804 => "1111110110010001",
51805 => "1111110110010010",
51806 => "1111110110010010",
51807 => "1111110110010010",
51808 => "1111110110010010",
51809 => "1111110110010010",
51810 => "1111110110010010",
51811 => "1111110110010010",
51812 => "1111110110010011",
51813 => "1111110110010011",
51814 => "1111110110010011",
51815 => "1111110110010011",
51816 => "1111110110010011",
51817 => "1111110110010011",
51818 => "1111110110010011",
51819 => "1111110110010100",
51820 => "1111110110010100",
51821 => "1111110110010100",
51822 => "1111110110010100",
51823 => "1111110110010100",
51824 => "1111110110010100",
51825 => "1111110110010101",
51826 => "1111110110010101",
51827 => "1111110110010101",
51828 => "1111110110010101",
51829 => "1111110110010101",
51830 => "1111110110010101",
51831 => "1111110110010101",
51832 => "1111110110010110",
51833 => "1111110110010110",
51834 => "1111110110010110",
51835 => "1111110110010110",
51836 => "1111110110010110",
51837 => "1111110110010110",
51838 => "1111110110010110",
51839 => "1111110110010111",
51840 => "1111110110010111",
51841 => "1111110110010111",
51842 => "1111110110010111",
51843 => "1111110110010111",
51844 => "1111110110010111",
51845 => "1111110110010111",
51846 => "1111110110011000",
51847 => "1111110110011000",
51848 => "1111110110011000",
51849 => "1111110110011000",
51850 => "1111110110011000",
51851 => "1111110110011000",
51852 => "1111110110011001",
51853 => "1111110110011001",
51854 => "1111110110011001",
51855 => "1111110110011001",
51856 => "1111110110011001",
51857 => "1111110110011001",
51858 => "1111110110011001",
51859 => "1111110110011010",
51860 => "1111110110011010",
51861 => "1111110110011010",
51862 => "1111110110011010",
51863 => "1111110110011010",
51864 => "1111110110011010",
51865 => "1111110110011010",
51866 => "1111110110011011",
51867 => "1111110110011011",
51868 => "1111110110011011",
51869 => "1111110110011011",
51870 => "1111110110011011",
51871 => "1111110110011011",
51872 => "1111110110011100",
51873 => "1111110110011100",
51874 => "1111110110011100",
51875 => "1111110110011100",
51876 => "1111110110011100",
51877 => "1111110110011100",
51878 => "1111110110011100",
51879 => "1111110110011101",
51880 => "1111110110011101",
51881 => "1111110110011101",
51882 => "1111110110011101",
51883 => "1111110110011101",
51884 => "1111110110011101",
51885 => "1111110110011101",
51886 => "1111110110011110",
51887 => "1111110110011110",
51888 => "1111110110011110",
51889 => "1111110110011110",
51890 => "1111110110011110",
51891 => "1111110110011110",
51892 => "1111110110011110",
51893 => "1111110110011111",
51894 => "1111110110011111",
51895 => "1111110110011111",
51896 => "1111110110011111",
51897 => "1111110110011111",
51898 => "1111110110011111",
51899 => "1111110110011111",
51900 => "1111110110100000",
51901 => "1111110110100000",
51902 => "1111110110100000",
51903 => "1111110110100000",
51904 => "1111110110100000",
51905 => "1111110110100000",
51906 => "1111110110100001",
51907 => "1111110110100001",
51908 => "1111110110100001",
51909 => "1111110110100001",
51910 => "1111110110100001",
51911 => "1111110110100001",
51912 => "1111110110100001",
51913 => "1111110110100010",
51914 => "1111110110100010",
51915 => "1111110110100010",
51916 => "1111110110100010",
51917 => "1111110110100010",
51918 => "1111110110100010",
51919 => "1111110110100010",
51920 => "1111110110100011",
51921 => "1111110110100011",
51922 => "1111110110100011",
51923 => "1111110110100011",
51924 => "1111110110100011",
51925 => "1111110110100011",
51926 => "1111110110100011",
51927 => "1111110110100100",
51928 => "1111110110100100",
51929 => "1111110110100100",
51930 => "1111110110100100",
51931 => "1111110110100100",
51932 => "1111110110100100",
51933 => "1111110110100100",
51934 => "1111110110100101",
51935 => "1111110110100101",
51936 => "1111110110100101",
51937 => "1111110110100101",
51938 => "1111110110100101",
51939 => "1111110110100101",
51940 => "1111110110100101",
51941 => "1111110110100110",
51942 => "1111110110100110",
51943 => "1111110110100110",
51944 => "1111110110100110",
51945 => "1111110110100110",
51946 => "1111110110100110",
51947 => "1111110110100111",
51948 => "1111110110100111",
51949 => "1111110110100111",
51950 => "1111110110100111",
51951 => "1111110110100111",
51952 => "1111110110100111",
51953 => "1111110110100111",
51954 => "1111110110101000",
51955 => "1111110110101000",
51956 => "1111110110101000",
51957 => "1111110110101000",
51958 => "1111110110101000",
51959 => "1111110110101000",
51960 => "1111110110101000",
51961 => "1111110110101001",
51962 => "1111110110101001",
51963 => "1111110110101001",
51964 => "1111110110101001",
51965 => "1111110110101001",
51966 => "1111110110101001",
51967 => "1111110110101001",
51968 => "1111110110101010",
51969 => "1111110110101010",
51970 => "1111110110101010",
51971 => "1111110110101010",
51972 => "1111110110101010",
51973 => "1111110110101010",
51974 => "1111110110101010",
51975 => "1111110110101011",
51976 => "1111110110101011",
51977 => "1111110110101011",
51978 => "1111110110101011",
51979 => "1111110110101011",
51980 => "1111110110101011",
51981 => "1111110110101011",
51982 => "1111110110101100",
51983 => "1111110110101100",
51984 => "1111110110101100",
51985 => "1111110110101100",
51986 => "1111110110101100",
51987 => "1111110110101100",
51988 => "1111110110101100",
51989 => "1111110110101101",
51990 => "1111110110101101",
51991 => "1111110110101101",
51992 => "1111110110101101",
51993 => "1111110110101101",
51994 => "1111110110101101",
51995 => "1111110110101101",
51996 => "1111110110101110",
51997 => "1111110110101110",
51998 => "1111110110101110",
51999 => "1111110110101110",
52000 => "1111110110101110",
52001 => "1111110110101110",
52002 => "1111110110101110",
52003 => "1111110110101111",
52004 => "1111110110101111",
52005 => "1111110110101111",
52006 => "1111110110101111",
52007 => "1111110110101111",
52008 => "1111110110101111",
52009 => "1111110110101111",
52010 => "1111110110110000",
52011 => "1111110110110000",
52012 => "1111110110110000",
52013 => "1111110110110000",
52014 => "1111110110110000",
52015 => "1111110110110000",
52016 => "1111110110110000",
52017 => "1111110110110001",
52018 => "1111110110110001",
52019 => "1111110110110001",
52020 => "1111110110110001",
52021 => "1111110110110001",
52022 => "1111110110110001",
52023 => "1111110110110001",
52024 => "1111110110110010",
52025 => "1111110110110010",
52026 => "1111110110110010",
52027 => "1111110110110010",
52028 => "1111110110110010",
52029 => "1111110110110010",
52030 => "1111110110110010",
52031 => "1111110110110011",
52032 => "1111110110110011",
52033 => "1111110110110011",
52034 => "1111110110110011",
52035 => "1111110110110011",
52036 => "1111110110110011",
52037 => "1111110110110011",
52038 => "1111110110110100",
52039 => "1111110110110100",
52040 => "1111110110110100",
52041 => "1111110110110100",
52042 => "1111110110110100",
52043 => "1111110110110100",
52044 => "1111110110110100",
52045 => "1111110110110101",
52046 => "1111110110110101",
52047 => "1111110110110101",
52048 => "1111110110110101",
52049 => "1111110110110101",
52050 => "1111110110110101",
52051 => "1111110110110101",
52052 => "1111110110110110",
52053 => "1111110110110110",
52054 => "1111110110110110",
52055 => "1111110110110110",
52056 => "1111110110110110",
52057 => "1111110110110110",
52058 => "1111110110110110",
52059 => "1111110110110111",
52060 => "1111110110110111",
52061 => "1111110110110111",
52062 => "1111110110110111",
52063 => "1111110110110111",
52064 => "1111110110110111",
52065 => "1111110110110111",
52066 => "1111110110111000",
52067 => "1111110110111000",
52068 => "1111110110111000",
52069 => "1111110110111000",
52070 => "1111110110111000",
52071 => "1111110110111000",
52072 => "1111110110111000",
52073 => "1111110110111001",
52074 => "1111110110111001",
52075 => "1111110110111001",
52076 => "1111110110111001",
52077 => "1111110110111001",
52078 => "1111110110111001",
52079 => "1111110110111001",
52080 => "1111110110111010",
52081 => "1111110110111010",
52082 => "1111110110111010",
52083 => "1111110110111010",
52084 => "1111110110111010",
52085 => "1111110110111010",
52086 => "1111110110111010",
52087 => "1111110110111011",
52088 => "1111110110111011",
52089 => "1111110110111011",
52090 => "1111110110111011",
52091 => "1111110110111011",
52092 => "1111110110111011",
52093 => "1111110110111011",
52094 => "1111110110111100",
52095 => "1111110110111100",
52096 => "1111110110111100",
52097 => "1111110110111100",
52098 => "1111110110111100",
52099 => "1111110110111100",
52100 => "1111110110111100",
52101 => "1111110110111100",
52102 => "1111110110111101",
52103 => "1111110110111101",
52104 => "1111110110111101",
52105 => "1111110110111101",
52106 => "1111110110111101",
52107 => "1111110110111101",
52108 => "1111110110111101",
52109 => "1111110110111110",
52110 => "1111110110111110",
52111 => "1111110110111110",
52112 => "1111110110111110",
52113 => "1111110110111110",
52114 => "1111110110111110",
52115 => "1111110110111110",
52116 => "1111110110111111",
52117 => "1111110110111111",
52118 => "1111110110111111",
52119 => "1111110110111111",
52120 => "1111110110111111",
52121 => "1111110110111111",
52122 => "1111110110111111",
52123 => "1111110111000000",
52124 => "1111110111000000",
52125 => "1111110111000000",
52126 => "1111110111000000",
52127 => "1111110111000000",
52128 => "1111110111000000",
52129 => "1111110111000000",
52130 => "1111110111000001",
52131 => "1111110111000001",
52132 => "1111110111000001",
52133 => "1111110111000001",
52134 => "1111110111000001",
52135 => "1111110111000001",
52136 => "1111110111000001",
52137 => "1111110111000010",
52138 => "1111110111000010",
52139 => "1111110111000010",
52140 => "1111110111000010",
52141 => "1111110111000010",
52142 => "1111110111000010",
52143 => "1111110111000010",
52144 => "1111110111000010",
52145 => "1111110111000011",
52146 => "1111110111000011",
52147 => "1111110111000011",
52148 => "1111110111000011",
52149 => "1111110111000011",
52150 => "1111110111000011",
52151 => "1111110111000011",
52152 => "1111110111000100",
52153 => "1111110111000100",
52154 => "1111110111000100",
52155 => "1111110111000100",
52156 => "1111110111000100",
52157 => "1111110111000100",
52158 => "1111110111000100",
52159 => "1111110111000101",
52160 => "1111110111000101",
52161 => "1111110111000101",
52162 => "1111110111000101",
52163 => "1111110111000101",
52164 => "1111110111000101",
52165 => "1111110111000101",
52166 => "1111110111000110",
52167 => "1111110111000110",
52168 => "1111110111000110",
52169 => "1111110111000110",
52170 => "1111110111000110",
52171 => "1111110111000110",
52172 => "1111110111000110",
52173 => "1111110111000110",
52174 => "1111110111000111",
52175 => "1111110111000111",
52176 => "1111110111000111",
52177 => "1111110111000111",
52178 => "1111110111000111",
52179 => "1111110111000111",
52180 => "1111110111000111",
52181 => "1111110111001000",
52182 => "1111110111001000",
52183 => "1111110111001000",
52184 => "1111110111001000",
52185 => "1111110111001000",
52186 => "1111110111001000",
52187 => "1111110111001000",
52188 => "1111110111001001",
52189 => "1111110111001001",
52190 => "1111110111001001",
52191 => "1111110111001001",
52192 => "1111110111001001",
52193 => "1111110111001001",
52194 => "1111110111001001",
52195 => "1111110111001010",
52196 => "1111110111001010",
52197 => "1111110111001010",
52198 => "1111110111001010",
52199 => "1111110111001010",
52200 => "1111110111001010",
52201 => "1111110111001010",
52202 => "1111110111001010",
52203 => "1111110111001011",
52204 => "1111110111001011",
52205 => "1111110111001011",
52206 => "1111110111001011",
52207 => "1111110111001011",
52208 => "1111110111001011",
52209 => "1111110111001011",
52210 => "1111110111001100",
52211 => "1111110111001100",
52212 => "1111110111001100",
52213 => "1111110111001100",
52214 => "1111110111001100",
52215 => "1111110111001100",
52216 => "1111110111001100",
52217 => "1111110111001101",
52218 => "1111110111001101",
52219 => "1111110111001101",
52220 => "1111110111001101",
52221 => "1111110111001101",
52222 => "1111110111001101",
52223 => "1111110111001101",
52224 => "1111110111001101",
52225 => "1111110111001110",
52226 => "1111110111001110",
52227 => "1111110111001110",
52228 => "1111110111001110",
52229 => "1111110111001110",
52230 => "1111110111001110",
52231 => "1111110111001110",
52232 => "1111110111001111",
52233 => "1111110111001111",
52234 => "1111110111001111",
52235 => "1111110111001111",
52236 => "1111110111001111",
52237 => "1111110111001111",
52238 => "1111110111001111",
52239 => "1111110111010000",
52240 => "1111110111010000",
52241 => "1111110111010000",
52242 => "1111110111010000",
52243 => "1111110111010000",
52244 => "1111110111010000",
52245 => "1111110111010000",
52246 => "1111110111010000",
52247 => "1111110111010001",
52248 => "1111110111010001",
52249 => "1111110111010001",
52250 => "1111110111010001",
52251 => "1111110111010001",
52252 => "1111110111010001",
52253 => "1111110111010001",
52254 => "1111110111010010",
52255 => "1111110111010010",
52256 => "1111110111010010",
52257 => "1111110111010010",
52258 => "1111110111010010",
52259 => "1111110111010010",
52260 => "1111110111010010",
52261 => "1111110111010010",
52262 => "1111110111010011",
52263 => "1111110111010011",
52264 => "1111110111010011",
52265 => "1111110111010011",
52266 => "1111110111010011",
52267 => "1111110111010011",
52268 => "1111110111010011",
52269 => "1111110111010100",
52270 => "1111110111010100",
52271 => "1111110111010100",
52272 => "1111110111010100",
52273 => "1111110111010100",
52274 => "1111110111010100",
52275 => "1111110111010100",
52276 => "1111110111010101",
52277 => "1111110111010101",
52278 => "1111110111010101",
52279 => "1111110111010101",
52280 => "1111110111010101",
52281 => "1111110111010101",
52282 => "1111110111010101",
52283 => "1111110111010101",
52284 => "1111110111010110",
52285 => "1111110111010110",
52286 => "1111110111010110",
52287 => "1111110111010110",
52288 => "1111110111010110",
52289 => "1111110111010110",
52290 => "1111110111010110",
52291 => "1111110111010111",
52292 => "1111110111010111",
52293 => "1111110111010111",
52294 => "1111110111010111",
52295 => "1111110111010111",
52296 => "1111110111010111",
52297 => "1111110111010111",
52298 => "1111110111010111",
52299 => "1111110111011000",
52300 => "1111110111011000",
52301 => "1111110111011000",
52302 => "1111110111011000",
52303 => "1111110111011000",
52304 => "1111110111011000",
52305 => "1111110111011000",
52306 => "1111110111011001",
52307 => "1111110111011001",
52308 => "1111110111011001",
52309 => "1111110111011001",
52310 => "1111110111011001",
52311 => "1111110111011001",
52312 => "1111110111011001",
52313 => "1111110111011001",
52314 => "1111110111011010",
52315 => "1111110111011010",
52316 => "1111110111011010",
52317 => "1111110111011010",
52318 => "1111110111011010",
52319 => "1111110111011010",
52320 => "1111110111011010",
52321 => "1111110111011011",
52322 => "1111110111011011",
52323 => "1111110111011011",
52324 => "1111110111011011",
52325 => "1111110111011011",
52326 => "1111110111011011",
52327 => "1111110111011011",
52328 => "1111110111011011",
52329 => "1111110111011100",
52330 => "1111110111011100",
52331 => "1111110111011100",
52332 => "1111110111011100",
52333 => "1111110111011100",
52334 => "1111110111011100",
52335 => "1111110111011100",
52336 => "1111110111011101",
52337 => "1111110111011101",
52338 => "1111110111011101",
52339 => "1111110111011101",
52340 => "1111110111011101",
52341 => "1111110111011101",
52342 => "1111110111011101",
52343 => "1111110111011101",
52344 => "1111110111011110",
52345 => "1111110111011110",
52346 => "1111110111011110",
52347 => "1111110111011110",
52348 => "1111110111011110",
52349 => "1111110111011110",
52350 => "1111110111011110",
52351 => "1111110111011110",
52352 => "1111110111011111",
52353 => "1111110111011111",
52354 => "1111110111011111",
52355 => "1111110111011111",
52356 => "1111110111011111",
52357 => "1111110111011111",
52358 => "1111110111011111",
52359 => "1111110111100000",
52360 => "1111110111100000",
52361 => "1111110111100000",
52362 => "1111110111100000",
52363 => "1111110111100000",
52364 => "1111110111100000",
52365 => "1111110111100000",
52366 => "1111110111100000",
52367 => "1111110111100001",
52368 => "1111110111100001",
52369 => "1111110111100001",
52370 => "1111110111100001",
52371 => "1111110111100001",
52372 => "1111110111100001",
52373 => "1111110111100001",
52374 => "1111110111100010",
52375 => "1111110111100010",
52376 => "1111110111100010",
52377 => "1111110111100010",
52378 => "1111110111100010",
52379 => "1111110111100010",
52380 => "1111110111100010",
52381 => "1111110111100010",
52382 => "1111110111100011",
52383 => "1111110111100011",
52384 => "1111110111100011",
52385 => "1111110111100011",
52386 => "1111110111100011",
52387 => "1111110111100011",
52388 => "1111110111100011",
52389 => "1111110111100011",
52390 => "1111110111100100",
52391 => "1111110111100100",
52392 => "1111110111100100",
52393 => "1111110111100100",
52394 => "1111110111100100",
52395 => "1111110111100100",
52396 => "1111110111100100",
52397 => "1111110111100101",
52398 => "1111110111100101",
52399 => "1111110111100101",
52400 => "1111110111100101",
52401 => "1111110111100101",
52402 => "1111110111100101",
52403 => "1111110111100101",
52404 => "1111110111100101",
52405 => "1111110111100110",
52406 => "1111110111100110",
52407 => "1111110111100110",
52408 => "1111110111100110",
52409 => "1111110111100110",
52410 => "1111110111100110",
52411 => "1111110111100110",
52412 => "1111110111100110",
52413 => "1111110111100111",
52414 => "1111110111100111",
52415 => "1111110111100111",
52416 => "1111110111100111",
52417 => "1111110111100111",
52418 => "1111110111100111",
52419 => "1111110111100111",
52420 => "1111110111101000",
52421 => "1111110111101000",
52422 => "1111110111101000",
52423 => "1111110111101000",
52424 => "1111110111101000",
52425 => "1111110111101000",
52426 => "1111110111101000",
52427 => "1111110111101000",
52428 => "1111110111101001",
52429 => "1111110111101001",
52430 => "1111110111101001",
52431 => "1111110111101001",
52432 => "1111110111101001",
52433 => "1111110111101001",
52434 => "1111110111101001",
52435 => "1111110111101001",
52436 => "1111110111101010",
52437 => "1111110111101010",
52438 => "1111110111101010",
52439 => "1111110111101010",
52440 => "1111110111101010",
52441 => "1111110111101010",
52442 => "1111110111101010",
52443 => "1111110111101010",
52444 => "1111110111101011",
52445 => "1111110111101011",
52446 => "1111110111101011",
52447 => "1111110111101011",
52448 => "1111110111101011",
52449 => "1111110111101011",
52450 => "1111110111101011",
52451 => "1111110111101100",
52452 => "1111110111101100",
52453 => "1111110111101100",
52454 => "1111110111101100",
52455 => "1111110111101100",
52456 => "1111110111101100",
52457 => "1111110111101100",
52458 => "1111110111101100",
52459 => "1111110111101101",
52460 => "1111110111101101",
52461 => "1111110111101101",
52462 => "1111110111101101",
52463 => "1111110111101101",
52464 => "1111110111101101",
52465 => "1111110111101101",
52466 => "1111110111101101",
52467 => "1111110111101110",
52468 => "1111110111101110",
52469 => "1111110111101110",
52470 => "1111110111101110",
52471 => "1111110111101110",
52472 => "1111110111101110",
52473 => "1111110111101110",
52474 => "1111110111101110",
52475 => "1111110111101111",
52476 => "1111110111101111",
52477 => "1111110111101111",
52478 => "1111110111101111",
52479 => "1111110111101111",
52480 => "1111110111101111",
52481 => "1111110111101111",
52482 => "1111110111110000",
52483 => "1111110111110000",
52484 => "1111110111110000",
52485 => "1111110111110000",
52486 => "1111110111110000",
52487 => "1111110111110000",
52488 => "1111110111110000",
52489 => "1111110111110000",
52490 => "1111110111110001",
52491 => "1111110111110001",
52492 => "1111110111110001",
52493 => "1111110111110001",
52494 => "1111110111110001",
52495 => "1111110111110001",
52496 => "1111110111110001",
52497 => "1111110111110001",
52498 => "1111110111110010",
52499 => "1111110111110010",
52500 => "1111110111110010",
52501 => "1111110111110010",
52502 => "1111110111110010",
52503 => "1111110111110010",
52504 => "1111110111110010",
52505 => "1111110111110010",
52506 => "1111110111110011",
52507 => "1111110111110011",
52508 => "1111110111110011",
52509 => "1111110111110011",
52510 => "1111110111110011",
52511 => "1111110111110011",
52512 => "1111110111110011",
52513 => "1111110111110011",
52514 => "1111110111110100",
52515 => "1111110111110100",
52516 => "1111110111110100",
52517 => "1111110111110100",
52518 => "1111110111110100",
52519 => "1111110111110100",
52520 => "1111110111110100",
52521 => "1111110111110100",
52522 => "1111110111110101",
52523 => "1111110111110101",
52524 => "1111110111110101",
52525 => "1111110111110101",
52526 => "1111110111110101",
52527 => "1111110111110101",
52528 => "1111110111110101",
52529 => "1111110111110101",
52530 => "1111110111110110",
52531 => "1111110111110110",
52532 => "1111110111110110",
52533 => "1111110111110110",
52534 => "1111110111110110",
52535 => "1111110111110110",
52536 => "1111110111110110",
52537 => "1111110111110110",
52538 => "1111110111110111",
52539 => "1111110111110111",
52540 => "1111110111110111",
52541 => "1111110111110111",
52542 => "1111110111110111",
52543 => "1111110111110111",
52544 => "1111110111110111",
52545 => "1111110111111000",
52546 => "1111110111111000",
52547 => "1111110111111000",
52548 => "1111110111111000",
52549 => "1111110111111000",
52550 => "1111110111111000",
52551 => "1111110111111000",
52552 => "1111110111111000",
52553 => "1111110111111001",
52554 => "1111110111111001",
52555 => "1111110111111001",
52556 => "1111110111111001",
52557 => "1111110111111001",
52558 => "1111110111111001",
52559 => "1111110111111001",
52560 => "1111110111111001",
52561 => "1111110111111010",
52562 => "1111110111111010",
52563 => "1111110111111010",
52564 => "1111110111111010",
52565 => "1111110111111010",
52566 => "1111110111111010",
52567 => "1111110111111010",
52568 => "1111110111111010",
52569 => "1111110111111011",
52570 => "1111110111111011",
52571 => "1111110111111011",
52572 => "1111110111111011",
52573 => "1111110111111011",
52574 => "1111110111111011",
52575 => "1111110111111011",
52576 => "1111110111111011",
52577 => "1111110111111100",
52578 => "1111110111111100",
52579 => "1111110111111100",
52580 => "1111110111111100",
52581 => "1111110111111100",
52582 => "1111110111111100",
52583 => "1111110111111100",
52584 => "1111110111111100",
52585 => "1111110111111101",
52586 => "1111110111111101",
52587 => "1111110111111101",
52588 => "1111110111111101",
52589 => "1111110111111101",
52590 => "1111110111111101",
52591 => "1111110111111101",
52592 => "1111110111111101",
52593 => "1111110111111110",
52594 => "1111110111111110",
52595 => "1111110111111110",
52596 => "1111110111111110",
52597 => "1111110111111110",
52598 => "1111110111111110",
52599 => "1111110111111110",
52600 => "1111110111111110",
52601 => "1111110111111111",
52602 => "1111110111111111",
52603 => "1111110111111111",
52604 => "1111110111111111",
52605 => "1111110111111111",
52606 => "1111110111111111",
52607 => "1111110111111111",
52608 => "1111110111111111",
52609 => "1111111000000000",
52610 => "1111111000000000",
52611 => "1111111000000000",
52612 => "1111111000000000",
52613 => "1111111000000000",
52614 => "1111111000000000",
52615 => "1111111000000000",
52616 => "1111111000000000",
52617 => "1111111000000000",
52618 => "1111111000000001",
52619 => "1111111000000001",
52620 => "1111111000000001",
52621 => "1111111000000001",
52622 => "1111111000000001",
52623 => "1111111000000001",
52624 => "1111111000000001",
52625 => "1111111000000001",
52626 => "1111111000000010",
52627 => "1111111000000010",
52628 => "1111111000000010",
52629 => "1111111000000010",
52630 => "1111111000000010",
52631 => "1111111000000010",
52632 => "1111111000000010",
52633 => "1111111000000010",
52634 => "1111111000000011",
52635 => "1111111000000011",
52636 => "1111111000000011",
52637 => "1111111000000011",
52638 => "1111111000000011",
52639 => "1111111000000011",
52640 => "1111111000000011",
52641 => "1111111000000011",
52642 => "1111111000000100",
52643 => "1111111000000100",
52644 => "1111111000000100",
52645 => "1111111000000100",
52646 => "1111111000000100",
52647 => "1111111000000100",
52648 => "1111111000000100",
52649 => "1111111000000100",
52650 => "1111111000000101",
52651 => "1111111000000101",
52652 => "1111111000000101",
52653 => "1111111000000101",
52654 => "1111111000000101",
52655 => "1111111000000101",
52656 => "1111111000000101",
52657 => "1111111000000101",
52658 => "1111111000000110",
52659 => "1111111000000110",
52660 => "1111111000000110",
52661 => "1111111000000110",
52662 => "1111111000000110",
52663 => "1111111000000110",
52664 => "1111111000000110",
52665 => "1111111000000110",
52666 => "1111111000000111",
52667 => "1111111000000111",
52668 => "1111111000000111",
52669 => "1111111000000111",
52670 => "1111111000000111",
52671 => "1111111000000111",
52672 => "1111111000000111",
52673 => "1111111000000111",
52674 => "1111111000001000",
52675 => "1111111000001000",
52676 => "1111111000001000",
52677 => "1111111000001000",
52678 => "1111111000001000",
52679 => "1111111000001000",
52680 => "1111111000001000",
52681 => "1111111000001000",
52682 => "1111111000001000",
52683 => "1111111000001001",
52684 => "1111111000001001",
52685 => "1111111000001001",
52686 => "1111111000001001",
52687 => "1111111000001001",
52688 => "1111111000001001",
52689 => "1111111000001001",
52690 => "1111111000001001",
52691 => "1111111000001010",
52692 => "1111111000001010",
52693 => "1111111000001010",
52694 => "1111111000001010",
52695 => "1111111000001010",
52696 => "1111111000001010",
52697 => "1111111000001010",
52698 => "1111111000001010",
52699 => "1111111000001011",
52700 => "1111111000001011",
52701 => "1111111000001011",
52702 => "1111111000001011",
52703 => "1111111000001011",
52704 => "1111111000001011",
52705 => "1111111000001011",
52706 => "1111111000001011",
52707 => "1111111000001100",
52708 => "1111111000001100",
52709 => "1111111000001100",
52710 => "1111111000001100",
52711 => "1111111000001100",
52712 => "1111111000001100",
52713 => "1111111000001100",
52714 => "1111111000001100",
52715 => "1111111000001100",
52716 => "1111111000001101",
52717 => "1111111000001101",
52718 => "1111111000001101",
52719 => "1111111000001101",
52720 => "1111111000001101",
52721 => "1111111000001101",
52722 => "1111111000001101",
52723 => "1111111000001101",
52724 => "1111111000001110",
52725 => "1111111000001110",
52726 => "1111111000001110",
52727 => "1111111000001110",
52728 => "1111111000001110",
52729 => "1111111000001110",
52730 => "1111111000001110",
52731 => "1111111000001110",
52732 => "1111111000001111",
52733 => "1111111000001111",
52734 => "1111111000001111",
52735 => "1111111000001111",
52736 => "1111111000001111",
52737 => "1111111000001111",
52738 => "1111111000001111",
52739 => "1111111000001111",
52740 => "1111111000001111",
52741 => "1111111000010000",
52742 => "1111111000010000",
52743 => "1111111000010000",
52744 => "1111111000010000",
52745 => "1111111000010000",
52746 => "1111111000010000",
52747 => "1111111000010000",
52748 => "1111111000010000",
52749 => "1111111000010001",
52750 => "1111111000010001",
52751 => "1111111000010001",
52752 => "1111111000010001",
52753 => "1111111000010001",
52754 => "1111111000010001",
52755 => "1111111000010001",
52756 => "1111111000010001",
52757 => "1111111000010010",
52758 => "1111111000010010",
52759 => "1111111000010010",
52760 => "1111111000010010",
52761 => "1111111000010010",
52762 => "1111111000010010",
52763 => "1111111000010010",
52764 => "1111111000010010",
52765 => "1111111000010010",
52766 => "1111111000010011",
52767 => "1111111000010011",
52768 => "1111111000010011",
52769 => "1111111000010011",
52770 => "1111111000010011",
52771 => "1111111000010011",
52772 => "1111111000010011",
52773 => "1111111000010011",
52774 => "1111111000010100",
52775 => "1111111000010100",
52776 => "1111111000010100",
52777 => "1111111000010100",
52778 => "1111111000010100",
52779 => "1111111000010100",
52780 => "1111111000010100",
52781 => "1111111000010100",
52782 => "1111111000010101",
52783 => "1111111000010101",
52784 => "1111111000010101",
52785 => "1111111000010101",
52786 => "1111111000010101",
52787 => "1111111000010101",
52788 => "1111111000010101",
52789 => "1111111000010101",
52790 => "1111111000010101",
52791 => "1111111000010110",
52792 => "1111111000010110",
52793 => "1111111000010110",
52794 => "1111111000010110",
52795 => "1111111000010110",
52796 => "1111111000010110",
52797 => "1111111000010110",
52798 => "1111111000010110",
52799 => "1111111000010111",
52800 => "1111111000010111",
52801 => "1111111000010111",
52802 => "1111111000010111",
52803 => "1111111000010111",
52804 => "1111111000010111",
52805 => "1111111000010111",
52806 => "1111111000010111",
52807 => "1111111000010111",
52808 => "1111111000011000",
52809 => "1111111000011000",
52810 => "1111111000011000",
52811 => "1111111000011000",
52812 => "1111111000011000",
52813 => "1111111000011000",
52814 => "1111111000011000",
52815 => "1111111000011000",
52816 => "1111111000011001",
52817 => "1111111000011001",
52818 => "1111111000011001",
52819 => "1111111000011001",
52820 => "1111111000011001",
52821 => "1111111000011001",
52822 => "1111111000011001",
52823 => "1111111000011001",
52824 => "1111111000011001",
52825 => "1111111000011010",
52826 => "1111111000011010",
52827 => "1111111000011010",
52828 => "1111111000011010",
52829 => "1111111000011010",
52830 => "1111111000011010",
52831 => "1111111000011010",
52832 => "1111111000011010",
52833 => "1111111000011011",
52834 => "1111111000011011",
52835 => "1111111000011011",
52836 => "1111111000011011",
52837 => "1111111000011011",
52838 => "1111111000011011",
52839 => "1111111000011011",
52840 => "1111111000011011",
52841 => "1111111000011011",
52842 => "1111111000011100",
52843 => "1111111000011100",
52844 => "1111111000011100",
52845 => "1111111000011100",
52846 => "1111111000011100",
52847 => "1111111000011100",
52848 => "1111111000011100",
52849 => "1111111000011100",
52850 => "1111111000011101",
52851 => "1111111000011101",
52852 => "1111111000011101",
52853 => "1111111000011101",
52854 => "1111111000011101",
52855 => "1111111000011101",
52856 => "1111111000011101",
52857 => "1111111000011101",
52858 => "1111111000011101",
52859 => "1111111000011110",
52860 => "1111111000011110",
52861 => "1111111000011110",
52862 => "1111111000011110",
52863 => "1111111000011110",
52864 => "1111111000011110",
52865 => "1111111000011110",
52866 => "1111111000011110",
52867 => "1111111000011111",
52868 => "1111111000011111",
52869 => "1111111000011111",
52870 => "1111111000011111",
52871 => "1111111000011111",
52872 => "1111111000011111",
52873 => "1111111000011111",
52874 => "1111111000011111",
52875 => "1111111000011111",
52876 => "1111111000100000",
52877 => "1111111000100000",
52878 => "1111111000100000",
52879 => "1111111000100000",
52880 => "1111111000100000",
52881 => "1111111000100000",
52882 => "1111111000100000",
52883 => "1111111000100000",
52884 => "1111111000100001",
52885 => "1111111000100001",
52886 => "1111111000100001",
52887 => "1111111000100001",
52888 => "1111111000100001",
52889 => "1111111000100001",
52890 => "1111111000100001",
52891 => "1111111000100001",
52892 => "1111111000100001",
52893 => "1111111000100010",
52894 => "1111111000100010",
52895 => "1111111000100010",
52896 => "1111111000100010",
52897 => "1111111000100010",
52898 => "1111111000100010",
52899 => "1111111000100010",
52900 => "1111111000100010",
52901 => "1111111000100010",
52902 => "1111111000100011",
52903 => "1111111000100011",
52904 => "1111111000100011",
52905 => "1111111000100011",
52906 => "1111111000100011",
52907 => "1111111000100011",
52908 => "1111111000100011",
52909 => "1111111000100011",
52910 => "1111111000100100",
52911 => "1111111000100100",
52912 => "1111111000100100",
52913 => "1111111000100100",
52914 => "1111111000100100",
52915 => "1111111000100100",
52916 => "1111111000100100",
52917 => "1111111000100100",
52918 => "1111111000100100",
52919 => "1111111000100101",
52920 => "1111111000100101",
52921 => "1111111000100101",
52922 => "1111111000100101",
52923 => "1111111000100101",
52924 => "1111111000100101",
52925 => "1111111000100101",
52926 => "1111111000100101",
52927 => "1111111000100101",
52928 => "1111111000100110",
52929 => "1111111000100110",
52930 => "1111111000100110",
52931 => "1111111000100110",
52932 => "1111111000100110",
52933 => "1111111000100110",
52934 => "1111111000100110",
52935 => "1111111000100110",
52936 => "1111111000100111",
52937 => "1111111000100111",
52938 => "1111111000100111",
52939 => "1111111000100111",
52940 => "1111111000100111",
52941 => "1111111000100111",
52942 => "1111111000100111",
52943 => "1111111000100111",
52944 => "1111111000100111",
52945 => "1111111000101000",
52946 => "1111111000101000",
52947 => "1111111000101000",
52948 => "1111111000101000",
52949 => "1111111000101000",
52950 => "1111111000101000",
52951 => "1111111000101000",
52952 => "1111111000101000",
52953 => "1111111000101000",
52954 => "1111111000101001",
52955 => "1111111000101001",
52956 => "1111111000101001",
52957 => "1111111000101001",
52958 => "1111111000101001",
52959 => "1111111000101001",
52960 => "1111111000101001",
52961 => "1111111000101001",
52962 => "1111111000101001",
52963 => "1111111000101010",
52964 => "1111111000101010",
52965 => "1111111000101010",
52966 => "1111111000101010",
52967 => "1111111000101010",
52968 => "1111111000101010",
52969 => "1111111000101010",
52970 => "1111111000101010",
52971 => "1111111000101011",
52972 => "1111111000101011",
52973 => "1111111000101011",
52974 => "1111111000101011",
52975 => "1111111000101011",
52976 => "1111111000101011",
52977 => "1111111000101011",
52978 => "1111111000101011",
52979 => "1111111000101011",
52980 => "1111111000101100",
52981 => "1111111000101100",
52982 => "1111111000101100",
52983 => "1111111000101100",
52984 => "1111111000101100",
52985 => "1111111000101100",
52986 => "1111111000101100",
52987 => "1111111000101100",
52988 => "1111111000101100",
52989 => "1111111000101101",
52990 => "1111111000101101",
52991 => "1111111000101101",
52992 => "1111111000101101",
52993 => "1111111000101101",
52994 => "1111111000101101",
52995 => "1111111000101101",
52996 => "1111111000101101",
52997 => "1111111000101101",
52998 => "1111111000101110",
52999 => "1111111000101110",
53000 => "1111111000101110",
53001 => "1111111000101110",
53002 => "1111111000101110",
53003 => "1111111000101110",
53004 => "1111111000101110",
53005 => "1111111000101110",
53006 => "1111111000101110",
53007 => "1111111000101111",
53008 => "1111111000101111",
53009 => "1111111000101111",
53010 => "1111111000101111",
53011 => "1111111000101111",
53012 => "1111111000101111",
53013 => "1111111000101111",
53014 => "1111111000101111",
53015 => "1111111000101111",
53016 => "1111111000110000",
53017 => "1111111000110000",
53018 => "1111111000110000",
53019 => "1111111000110000",
53020 => "1111111000110000",
53021 => "1111111000110000",
53022 => "1111111000110000",
53023 => "1111111000110000",
53024 => "1111111000110000",
53025 => "1111111000110001",
53026 => "1111111000110001",
53027 => "1111111000110001",
53028 => "1111111000110001",
53029 => "1111111000110001",
53030 => "1111111000110001",
53031 => "1111111000110001",
53032 => "1111111000110001",
53033 => "1111111000110001",
53034 => "1111111000110010",
53035 => "1111111000110010",
53036 => "1111111000110010",
53037 => "1111111000110010",
53038 => "1111111000110010",
53039 => "1111111000110010",
53040 => "1111111000110010",
53041 => "1111111000110010",
53042 => "1111111000110011",
53043 => "1111111000110011",
53044 => "1111111000110011",
53045 => "1111111000110011",
53046 => "1111111000110011",
53047 => "1111111000110011",
53048 => "1111111000110011",
53049 => "1111111000110011",
53050 => "1111111000110011",
53051 => "1111111000110100",
53052 => "1111111000110100",
53053 => "1111111000110100",
53054 => "1111111000110100",
53055 => "1111111000110100",
53056 => "1111111000110100",
53057 => "1111111000110100",
53058 => "1111111000110100",
53059 => "1111111000110100",
53060 => "1111111000110101",
53061 => "1111111000110101",
53062 => "1111111000110101",
53063 => "1111111000110101",
53064 => "1111111000110101",
53065 => "1111111000110101",
53066 => "1111111000110101",
53067 => "1111111000110101",
53068 => "1111111000110101",
53069 => "1111111000110110",
53070 => "1111111000110110",
53071 => "1111111000110110",
53072 => "1111111000110110",
53073 => "1111111000110110",
53074 => "1111111000110110",
53075 => "1111111000110110",
53076 => "1111111000110110",
53077 => "1111111000110110",
53078 => "1111111000110111",
53079 => "1111111000110111",
53080 => "1111111000110111",
53081 => "1111111000110111",
53082 => "1111111000110111",
53083 => "1111111000110111",
53084 => "1111111000110111",
53085 => "1111111000110111",
53086 => "1111111000110111",
53087 => "1111111000111000",
53088 => "1111111000111000",
53089 => "1111111000111000",
53090 => "1111111000111000",
53091 => "1111111000111000",
53092 => "1111111000111000",
53093 => "1111111000111000",
53094 => "1111111000111000",
53095 => "1111111000111000",
53096 => "1111111000111000",
53097 => "1111111000111001",
53098 => "1111111000111001",
53099 => "1111111000111001",
53100 => "1111111000111001",
53101 => "1111111000111001",
53102 => "1111111000111001",
53103 => "1111111000111001",
53104 => "1111111000111001",
53105 => "1111111000111001",
53106 => "1111111000111010",
53107 => "1111111000111010",
53108 => "1111111000111010",
53109 => "1111111000111010",
53110 => "1111111000111010",
53111 => "1111111000111010",
53112 => "1111111000111010",
53113 => "1111111000111010",
53114 => "1111111000111010",
53115 => "1111111000111011",
53116 => "1111111000111011",
53117 => "1111111000111011",
53118 => "1111111000111011",
53119 => "1111111000111011",
53120 => "1111111000111011",
53121 => "1111111000111011",
53122 => "1111111000111011",
53123 => "1111111000111011",
53124 => "1111111000111100",
53125 => "1111111000111100",
53126 => "1111111000111100",
53127 => "1111111000111100",
53128 => "1111111000111100",
53129 => "1111111000111100",
53130 => "1111111000111100",
53131 => "1111111000111100",
53132 => "1111111000111100",
53133 => "1111111000111101",
53134 => "1111111000111101",
53135 => "1111111000111101",
53136 => "1111111000111101",
53137 => "1111111000111101",
53138 => "1111111000111101",
53139 => "1111111000111101",
53140 => "1111111000111101",
53141 => "1111111000111101",
53142 => "1111111000111110",
53143 => "1111111000111110",
53144 => "1111111000111110",
53145 => "1111111000111110",
53146 => "1111111000111110",
53147 => "1111111000111110",
53148 => "1111111000111110",
53149 => "1111111000111110",
53150 => "1111111000111110",
53151 => "1111111000111111",
53152 => "1111111000111111",
53153 => "1111111000111111",
53154 => "1111111000111111",
53155 => "1111111000111111",
53156 => "1111111000111111",
53157 => "1111111000111111",
53158 => "1111111000111111",
53159 => "1111111000111111",
53160 => "1111111001000000",
53161 => "1111111001000000",
53162 => "1111111001000000",
53163 => "1111111001000000",
53164 => "1111111001000000",
53165 => "1111111001000000",
53166 => "1111111001000000",
53167 => "1111111001000000",
53168 => "1111111001000000",
53169 => "1111111001000000",
53170 => "1111111001000001",
53171 => "1111111001000001",
53172 => "1111111001000001",
53173 => "1111111001000001",
53174 => "1111111001000001",
53175 => "1111111001000001",
53176 => "1111111001000001",
53177 => "1111111001000001",
53178 => "1111111001000001",
53179 => "1111111001000010",
53180 => "1111111001000010",
53181 => "1111111001000010",
53182 => "1111111001000010",
53183 => "1111111001000010",
53184 => "1111111001000010",
53185 => "1111111001000010",
53186 => "1111111001000010",
53187 => "1111111001000010",
53188 => "1111111001000011",
53189 => "1111111001000011",
53190 => "1111111001000011",
53191 => "1111111001000011",
53192 => "1111111001000011",
53193 => "1111111001000011",
53194 => "1111111001000011",
53195 => "1111111001000011",
53196 => "1111111001000011",
53197 => "1111111001000100",
53198 => "1111111001000100",
53199 => "1111111001000100",
53200 => "1111111001000100",
53201 => "1111111001000100",
53202 => "1111111001000100",
53203 => "1111111001000100",
53204 => "1111111001000100",
53205 => "1111111001000100",
53206 => "1111111001000100",
53207 => "1111111001000101",
53208 => "1111111001000101",
53209 => "1111111001000101",
53210 => "1111111001000101",
53211 => "1111111001000101",
53212 => "1111111001000101",
53213 => "1111111001000101",
53214 => "1111111001000101",
53215 => "1111111001000101",
53216 => "1111111001000110",
53217 => "1111111001000110",
53218 => "1111111001000110",
53219 => "1111111001000110",
53220 => "1111111001000110",
53221 => "1111111001000110",
53222 => "1111111001000110",
53223 => "1111111001000110",
53224 => "1111111001000110",
53225 => "1111111001000111",
53226 => "1111111001000111",
53227 => "1111111001000111",
53228 => "1111111001000111",
53229 => "1111111001000111",
53230 => "1111111001000111",
53231 => "1111111001000111",
53232 => "1111111001000111",
53233 => "1111111001000111",
53234 => "1111111001000111",
53235 => "1111111001001000",
53236 => "1111111001001000",
53237 => "1111111001001000",
53238 => "1111111001001000",
53239 => "1111111001001000",
53240 => "1111111001001000",
53241 => "1111111001001000",
53242 => "1111111001001000",
53243 => "1111111001001000",
53244 => "1111111001001001",
53245 => "1111111001001001",
53246 => "1111111001001001",
53247 => "1111111001001001",
53248 => "1111111001001001",
53249 => "1111111001001001",
53250 => "1111111001001001",
53251 => "1111111001001001",
53252 => "1111111001001001",
53253 => "1111111001001001",
53254 => "1111111001001010",
53255 => "1111111001001010",
53256 => "1111111001001010",
53257 => "1111111001001010",
53258 => "1111111001001010",
53259 => "1111111001001010",
53260 => "1111111001001010",
53261 => "1111111001001010",
53262 => "1111111001001010",
53263 => "1111111001001011",
53264 => "1111111001001011",
53265 => "1111111001001011",
53266 => "1111111001001011",
53267 => "1111111001001011",
53268 => "1111111001001011",
53269 => "1111111001001011",
53270 => "1111111001001011",
53271 => "1111111001001011",
53272 => "1111111001001100",
53273 => "1111111001001100",
53274 => "1111111001001100",
53275 => "1111111001001100",
53276 => "1111111001001100",
53277 => "1111111001001100",
53278 => "1111111001001100",
53279 => "1111111001001100",
53280 => "1111111001001100",
53281 => "1111111001001100",
53282 => "1111111001001101",
53283 => "1111111001001101",
53284 => "1111111001001101",
53285 => "1111111001001101",
53286 => "1111111001001101",
53287 => "1111111001001101",
53288 => "1111111001001101",
53289 => "1111111001001101",
53290 => "1111111001001101",
53291 => "1111111001001110",
53292 => "1111111001001110",
53293 => "1111111001001110",
53294 => "1111111001001110",
53295 => "1111111001001110",
53296 => "1111111001001110",
53297 => "1111111001001110",
53298 => "1111111001001110",
53299 => "1111111001001110",
53300 => "1111111001001110",
53301 => "1111111001001111",
53302 => "1111111001001111",
53303 => "1111111001001111",
53304 => "1111111001001111",
53305 => "1111111001001111",
53306 => "1111111001001111",
53307 => "1111111001001111",
53308 => "1111111001001111",
53309 => "1111111001001111",
53310 => "1111111001010000",
53311 => "1111111001010000",
53312 => "1111111001010000",
53313 => "1111111001010000",
53314 => "1111111001010000",
53315 => "1111111001010000",
53316 => "1111111001010000",
53317 => "1111111001010000",
53318 => "1111111001010000",
53319 => "1111111001010000",
53320 => "1111111001010001",
53321 => "1111111001010001",
53322 => "1111111001010001",
53323 => "1111111001010001",
53324 => "1111111001010001",
53325 => "1111111001010001",
53326 => "1111111001010001",
53327 => "1111111001010001",
53328 => "1111111001010001",
53329 => "1111111001010001",
53330 => "1111111001010010",
53331 => "1111111001010010",
53332 => "1111111001010010",
53333 => "1111111001010010",
53334 => "1111111001010010",
53335 => "1111111001010010",
53336 => "1111111001010010",
53337 => "1111111001010010",
53338 => "1111111001010010",
53339 => "1111111001010011",
53340 => "1111111001010011",
53341 => "1111111001010011",
53342 => "1111111001010011",
53343 => "1111111001010011",
53344 => "1111111001010011",
53345 => "1111111001010011",
53346 => "1111111001010011",
53347 => "1111111001010011",
53348 => "1111111001010011",
53349 => "1111111001010100",
53350 => "1111111001010100",
53351 => "1111111001010100",
53352 => "1111111001010100",
53353 => "1111111001010100",
53354 => "1111111001010100",
53355 => "1111111001010100",
53356 => "1111111001010100",
53357 => "1111111001010100",
53358 => "1111111001010101",
53359 => "1111111001010101",
53360 => "1111111001010101",
53361 => "1111111001010101",
53362 => "1111111001010101",
53363 => "1111111001010101",
53364 => "1111111001010101",
53365 => "1111111001010101",
53366 => "1111111001010101",
53367 => "1111111001010101",
53368 => "1111111001010110",
53369 => "1111111001010110",
53370 => "1111111001010110",
53371 => "1111111001010110",
53372 => "1111111001010110",
53373 => "1111111001010110",
53374 => "1111111001010110",
53375 => "1111111001010110",
53376 => "1111111001010110",
53377 => "1111111001010110",
53378 => "1111111001010111",
53379 => "1111111001010111",
53380 => "1111111001010111",
53381 => "1111111001010111",
53382 => "1111111001010111",
53383 => "1111111001010111",
53384 => "1111111001010111",
53385 => "1111111001010111",
53386 => "1111111001010111",
53387 => "1111111001011000",
53388 => "1111111001011000",
53389 => "1111111001011000",
53390 => "1111111001011000",
53391 => "1111111001011000",
53392 => "1111111001011000",
53393 => "1111111001011000",
53394 => "1111111001011000",
53395 => "1111111001011000",
53396 => "1111111001011000",
53397 => "1111111001011001",
53398 => "1111111001011001",
53399 => "1111111001011001",
53400 => "1111111001011001",
53401 => "1111111001011001",
53402 => "1111111001011001",
53403 => "1111111001011001",
53404 => "1111111001011001",
53405 => "1111111001011001",
53406 => "1111111001011001",
53407 => "1111111001011010",
53408 => "1111111001011010",
53409 => "1111111001011010",
53410 => "1111111001011010",
53411 => "1111111001011010",
53412 => "1111111001011010",
53413 => "1111111001011010",
53414 => "1111111001011010",
53415 => "1111111001011010",
53416 => "1111111001011010",
53417 => "1111111001011011",
53418 => "1111111001011011",
53419 => "1111111001011011",
53420 => "1111111001011011",
53421 => "1111111001011011",
53422 => "1111111001011011",
53423 => "1111111001011011",
53424 => "1111111001011011",
53425 => "1111111001011011",
53426 => "1111111001011011",
53427 => "1111111001011100",
53428 => "1111111001011100",
53429 => "1111111001011100",
53430 => "1111111001011100",
53431 => "1111111001011100",
53432 => "1111111001011100",
53433 => "1111111001011100",
53434 => "1111111001011100",
53435 => "1111111001011100",
53436 => "1111111001011101",
53437 => "1111111001011101",
53438 => "1111111001011101",
53439 => "1111111001011101",
53440 => "1111111001011101",
53441 => "1111111001011101",
53442 => "1111111001011101",
53443 => "1111111001011101",
53444 => "1111111001011101",
53445 => "1111111001011101",
53446 => "1111111001011110",
53447 => "1111111001011110",
53448 => "1111111001011110",
53449 => "1111111001011110",
53450 => "1111111001011110",
53451 => "1111111001011110",
53452 => "1111111001011110",
53453 => "1111111001011110",
53454 => "1111111001011110",
53455 => "1111111001011110",
53456 => "1111111001011111",
53457 => "1111111001011111",
53458 => "1111111001011111",
53459 => "1111111001011111",
53460 => "1111111001011111",
53461 => "1111111001011111",
53462 => "1111111001011111",
53463 => "1111111001011111",
53464 => "1111111001011111",
53465 => "1111111001011111",
53466 => "1111111001100000",
53467 => "1111111001100000",
53468 => "1111111001100000",
53469 => "1111111001100000",
53470 => "1111111001100000",
53471 => "1111111001100000",
53472 => "1111111001100000",
53473 => "1111111001100000",
53474 => "1111111001100000",
53475 => "1111111001100000",
53476 => "1111111001100001",
53477 => "1111111001100001",
53478 => "1111111001100001",
53479 => "1111111001100001",
53480 => "1111111001100001",
53481 => "1111111001100001",
53482 => "1111111001100001",
53483 => "1111111001100001",
53484 => "1111111001100001",
53485 => "1111111001100001",
53486 => "1111111001100010",
53487 => "1111111001100010",
53488 => "1111111001100010",
53489 => "1111111001100010",
53490 => "1111111001100010",
53491 => "1111111001100010",
53492 => "1111111001100010",
53493 => "1111111001100010",
53494 => "1111111001100010",
53495 => "1111111001100010",
53496 => "1111111001100011",
53497 => "1111111001100011",
53498 => "1111111001100011",
53499 => "1111111001100011",
53500 => "1111111001100011",
53501 => "1111111001100011",
53502 => "1111111001100011",
53503 => "1111111001100011",
53504 => "1111111001100011",
53505 => "1111111001100011",
53506 => "1111111001100100",
53507 => "1111111001100100",
53508 => "1111111001100100",
53509 => "1111111001100100",
53510 => "1111111001100100",
53511 => "1111111001100100",
53512 => "1111111001100100",
53513 => "1111111001100100",
53514 => "1111111001100100",
53515 => "1111111001100100",
53516 => "1111111001100101",
53517 => "1111111001100101",
53518 => "1111111001100101",
53519 => "1111111001100101",
53520 => "1111111001100101",
53521 => "1111111001100101",
53522 => "1111111001100101",
53523 => "1111111001100101",
53524 => "1111111001100101",
53525 => "1111111001100101",
53526 => "1111111001100110",
53527 => "1111111001100110",
53528 => "1111111001100110",
53529 => "1111111001100110",
53530 => "1111111001100110",
53531 => "1111111001100110",
53532 => "1111111001100110",
53533 => "1111111001100110",
53534 => "1111111001100110",
53535 => "1111111001100110",
53536 => "1111111001100111",
53537 => "1111111001100111",
53538 => "1111111001100111",
53539 => "1111111001100111",
53540 => "1111111001100111",
53541 => "1111111001100111",
53542 => "1111111001100111",
53543 => "1111111001100111",
53544 => "1111111001100111",
53545 => "1111111001100111",
53546 => "1111111001101000",
53547 => "1111111001101000",
53548 => "1111111001101000",
53549 => "1111111001101000",
53550 => "1111111001101000",
53551 => "1111111001101000",
53552 => "1111111001101000",
53553 => "1111111001101000",
53554 => "1111111001101000",
53555 => "1111111001101000",
53556 => "1111111001101001",
53557 => "1111111001101001",
53558 => "1111111001101001",
53559 => "1111111001101001",
53560 => "1111111001101001",
53561 => "1111111001101001",
53562 => "1111111001101001",
53563 => "1111111001101001",
53564 => "1111111001101001",
53565 => "1111111001101001",
53566 => "1111111001101010",
53567 => "1111111001101010",
53568 => "1111111001101010",
53569 => "1111111001101010",
53570 => "1111111001101010",
53571 => "1111111001101010",
53572 => "1111111001101010",
53573 => "1111111001101010",
53574 => "1111111001101010",
53575 => "1111111001101010",
53576 => "1111111001101011",
53577 => "1111111001101011",
53578 => "1111111001101011",
53579 => "1111111001101011",
53580 => "1111111001101011",
53581 => "1111111001101011",
53582 => "1111111001101011",
53583 => "1111111001101011",
53584 => "1111111001101011",
53585 => "1111111001101011",
53586 => "1111111001101011",
53587 => "1111111001101100",
53588 => "1111111001101100",
53589 => "1111111001101100",
53590 => "1111111001101100",
53591 => "1111111001101100",
53592 => "1111111001101100",
53593 => "1111111001101100",
53594 => "1111111001101100",
53595 => "1111111001101100",
53596 => "1111111001101100",
53597 => "1111111001101101",
53598 => "1111111001101101",
53599 => "1111111001101101",
53600 => "1111111001101101",
53601 => "1111111001101101",
53602 => "1111111001101101",
53603 => "1111111001101101",
53604 => "1111111001101101",
53605 => "1111111001101101",
53606 => "1111111001101101",
53607 => "1111111001101110",
53608 => "1111111001101110",
53609 => "1111111001101110",
53610 => "1111111001101110",
53611 => "1111111001101110",
53612 => "1111111001101110",
53613 => "1111111001101110",
53614 => "1111111001101110",
53615 => "1111111001101110",
53616 => "1111111001101110",
53617 => "1111111001101111",
53618 => "1111111001101111",
53619 => "1111111001101111",
53620 => "1111111001101111",
53621 => "1111111001101111",
53622 => "1111111001101111",
53623 => "1111111001101111",
53624 => "1111111001101111",
53625 => "1111111001101111",
53626 => "1111111001101111",
53627 => "1111111001101111",
53628 => "1111111001110000",
53629 => "1111111001110000",
53630 => "1111111001110000",
53631 => "1111111001110000",
53632 => "1111111001110000",
53633 => "1111111001110000",
53634 => "1111111001110000",
53635 => "1111111001110000",
53636 => "1111111001110000",
53637 => "1111111001110000",
53638 => "1111111001110001",
53639 => "1111111001110001",
53640 => "1111111001110001",
53641 => "1111111001110001",
53642 => "1111111001110001",
53643 => "1111111001110001",
53644 => "1111111001110001",
53645 => "1111111001110001",
53646 => "1111111001110001",
53647 => "1111111001110001",
53648 => "1111111001110010",
53649 => "1111111001110010",
53650 => "1111111001110010",
53651 => "1111111001110010",
53652 => "1111111001110010",
53653 => "1111111001110010",
53654 => "1111111001110010",
53655 => "1111111001110010",
53656 => "1111111001110010",
53657 => "1111111001110010",
53658 => "1111111001110010",
53659 => "1111111001110011",
53660 => "1111111001110011",
53661 => "1111111001110011",
53662 => "1111111001110011",
53663 => "1111111001110011",
53664 => "1111111001110011",
53665 => "1111111001110011",
53666 => "1111111001110011",
53667 => "1111111001110011",
53668 => "1111111001110011",
53669 => "1111111001110100",
53670 => "1111111001110100",
53671 => "1111111001110100",
53672 => "1111111001110100",
53673 => "1111111001110100",
53674 => "1111111001110100",
53675 => "1111111001110100",
53676 => "1111111001110100",
53677 => "1111111001110100",
53678 => "1111111001110100",
53679 => "1111111001110101",
53680 => "1111111001110101",
53681 => "1111111001110101",
53682 => "1111111001110101",
53683 => "1111111001110101",
53684 => "1111111001110101",
53685 => "1111111001110101",
53686 => "1111111001110101",
53687 => "1111111001110101",
53688 => "1111111001110101",
53689 => "1111111001110101",
53690 => "1111111001110110",
53691 => "1111111001110110",
53692 => "1111111001110110",
53693 => "1111111001110110",
53694 => "1111111001110110",
53695 => "1111111001110110",
53696 => "1111111001110110",
53697 => "1111111001110110",
53698 => "1111111001110110",
53699 => "1111111001110110",
53700 => "1111111001110111",
53701 => "1111111001110111",
53702 => "1111111001110111",
53703 => "1111111001110111",
53704 => "1111111001110111",
53705 => "1111111001110111",
53706 => "1111111001110111",
53707 => "1111111001110111",
53708 => "1111111001110111",
53709 => "1111111001110111",
53710 => "1111111001110111",
53711 => "1111111001111000",
53712 => "1111111001111000",
53713 => "1111111001111000",
53714 => "1111111001111000",
53715 => "1111111001111000",
53716 => "1111111001111000",
53717 => "1111111001111000",
53718 => "1111111001111000",
53719 => "1111111001111000",
53720 => "1111111001111000",
53721 => "1111111001111001",
53722 => "1111111001111001",
53723 => "1111111001111001",
53724 => "1111111001111001",
53725 => "1111111001111001",
53726 => "1111111001111001",
53727 => "1111111001111001",
53728 => "1111111001111001",
53729 => "1111111001111001",
53730 => "1111111001111001",
53731 => "1111111001111001",
53732 => "1111111001111010",
53733 => "1111111001111010",
53734 => "1111111001111010",
53735 => "1111111001111010",
53736 => "1111111001111010",
53737 => "1111111001111010",
53738 => "1111111001111010",
53739 => "1111111001111010",
53740 => "1111111001111010",
53741 => "1111111001111010",
53742 => "1111111001111010",
53743 => "1111111001111011",
53744 => "1111111001111011",
53745 => "1111111001111011",
53746 => "1111111001111011",
53747 => "1111111001111011",
53748 => "1111111001111011",
53749 => "1111111001111011",
53750 => "1111111001111011",
53751 => "1111111001111011",
53752 => "1111111001111011",
53753 => "1111111001111100",
53754 => "1111111001111100",
53755 => "1111111001111100",
53756 => "1111111001111100",
53757 => "1111111001111100",
53758 => "1111111001111100",
53759 => "1111111001111100",
53760 => "1111111001111100",
53761 => "1111111001111100",
53762 => "1111111001111100",
53763 => "1111111001111100",
53764 => "1111111001111101",
53765 => "1111111001111101",
53766 => "1111111001111101",
53767 => "1111111001111101",
53768 => "1111111001111101",
53769 => "1111111001111101",
53770 => "1111111001111101",
53771 => "1111111001111101",
53772 => "1111111001111101",
53773 => "1111111001111101",
53774 => "1111111001111110",
53775 => "1111111001111110",
53776 => "1111111001111110",
53777 => "1111111001111110",
53778 => "1111111001111110",
53779 => "1111111001111110",
53780 => "1111111001111110",
53781 => "1111111001111110",
53782 => "1111111001111110",
53783 => "1111111001111110",
53784 => "1111111001111110",
53785 => "1111111001111111",
53786 => "1111111001111111",
53787 => "1111111001111111",
53788 => "1111111001111111",
53789 => "1111111001111111",
53790 => "1111111001111111",
53791 => "1111111001111111",
53792 => "1111111001111111",
53793 => "1111111001111111",
53794 => "1111111001111111",
53795 => "1111111001111111",
53796 => "1111111010000000",
53797 => "1111111010000000",
53798 => "1111111010000000",
53799 => "1111111010000000",
53800 => "1111111010000000",
53801 => "1111111010000000",
53802 => "1111111010000000",
53803 => "1111111010000000",
53804 => "1111111010000000",
53805 => "1111111010000000",
53806 => "1111111010000000",
53807 => "1111111010000001",
53808 => "1111111010000001",
53809 => "1111111010000001",
53810 => "1111111010000001",
53811 => "1111111010000001",
53812 => "1111111010000001",
53813 => "1111111010000001",
53814 => "1111111010000001",
53815 => "1111111010000001",
53816 => "1111111010000001",
53817 => "1111111010000010",
53818 => "1111111010000010",
53819 => "1111111010000010",
53820 => "1111111010000010",
53821 => "1111111010000010",
53822 => "1111111010000010",
53823 => "1111111010000010",
53824 => "1111111010000010",
53825 => "1111111010000010",
53826 => "1111111010000010",
53827 => "1111111010000010",
53828 => "1111111010000011",
53829 => "1111111010000011",
53830 => "1111111010000011",
53831 => "1111111010000011",
53832 => "1111111010000011",
53833 => "1111111010000011",
53834 => "1111111010000011",
53835 => "1111111010000011",
53836 => "1111111010000011",
53837 => "1111111010000011",
53838 => "1111111010000011",
53839 => "1111111010000100",
53840 => "1111111010000100",
53841 => "1111111010000100",
53842 => "1111111010000100",
53843 => "1111111010000100",
53844 => "1111111010000100",
53845 => "1111111010000100",
53846 => "1111111010000100",
53847 => "1111111010000100",
53848 => "1111111010000100",
53849 => "1111111010000100",
53850 => "1111111010000101",
53851 => "1111111010000101",
53852 => "1111111010000101",
53853 => "1111111010000101",
53854 => "1111111010000101",
53855 => "1111111010000101",
53856 => "1111111010000101",
53857 => "1111111010000101",
53858 => "1111111010000101",
53859 => "1111111010000101",
53860 => "1111111010000101",
53861 => "1111111010000110",
53862 => "1111111010000110",
53863 => "1111111010000110",
53864 => "1111111010000110",
53865 => "1111111010000110",
53866 => "1111111010000110",
53867 => "1111111010000110",
53868 => "1111111010000110",
53869 => "1111111010000110",
53870 => "1111111010000110",
53871 => "1111111010000110",
53872 => "1111111010000111",
53873 => "1111111010000111",
53874 => "1111111010000111",
53875 => "1111111010000111",
53876 => "1111111010000111",
53877 => "1111111010000111",
53878 => "1111111010000111",
53879 => "1111111010000111",
53880 => "1111111010000111",
53881 => "1111111010000111",
53882 => "1111111010000111",
53883 => "1111111010001000",
53884 => "1111111010001000",
53885 => "1111111010001000",
53886 => "1111111010001000",
53887 => "1111111010001000",
53888 => "1111111010001000",
53889 => "1111111010001000",
53890 => "1111111010001000",
53891 => "1111111010001000",
53892 => "1111111010001000",
53893 => "1111111010001000",
53894 => "1111111010001001",
53895 => "1111111010001001",
53896 => "1111111010001001",
53897 => "1111111010001001",
53898 => "1111111010001001",
53899 => "1111111010001001",
53900 => "1111111010001001",
53901 => "1111111010001001",
53902 => "1111111010001001",
53903 => "1111111010001001",
53904 => "1111111010001001",
53905 => "1111111010001010",
53906 => "1111111010001010",
53907 => "1111111010001010",
53908 => "1111111010001010",
53909 => "1111111010001010",
53910 => "1111111010001010",
53911 => "1111111010001010",
53912 => "1111111010001010",
53913 => "1111111010001010",
53914 => "1111111010001010",
53915 => "1111111010001010",
53916 => "1111111010001011",
53917 => "1111111010001011",
53918 => "1111111010001011",
53919 => "1111111010001011",
53920 => "1111111010001011",
53921 => "1111111010001011",
53922 => "1111111010001011",
53923 => "1111111010001011",
53924 => "1111111010001011",
53925 => "1111111010001011",
53926 => "1111111010001011",
53927 => "1111111010001100",
53928 => "1111111010001100",
53929 => "1111111010001100",
53930 => "1111111010001100",
53931 => "1111111010001100",
53932 => "1111111010001100",
53933 => "1111111010001100",
53934 => "1111111010001100",
53935 => "1111111010001100",
53936 => "1111111010001100",
53937 => "1111111010001100",
53938 => "1111111010001101",
53939 => "1111111010001101",
53940 => "1111111010001101",
53941 => "1111111010001101",
53942 => "1111111010001101",
53943 => "1111111010001101",
53944 => "1111111010001101",
53945 => "1111111010001101",
53946 => "1111111010001101",
53947 => "1111111010001101",
53948 => "1111111010001101",
53949 => "1111111010001110",
53950 => "1111111010001110",
53951 => "1111111010001110",
53952 => "1111111010001110",
53953 => "1111111010001110",
53954 => "1111111010001110",
53955 => "1111111010001110",
53956 => "1111111010001110",
53957 => "1111111010001110",
53958 => "1111111010001110",
53959 => "1111111010001110",
53960 => "1111111010001111",
53961 => "1111111010001111",
53962 => "1111111010001111",
53963 => "1111111010001111",
53964 => "1111111010001111",
53965 => "1111111010001111",
53966 => "1111111010001111",
53967 => "1111111010001111",
53968 => "1111111010001111",
53969 => "1111111010001111",
53970 => "1111111010001111",
53971 => "1111111010010000",
53972 => "1111111010010000",
53973 => "1111111010010000",
53974 => "1111111010010000",
53975 => "1111111010010000",
53976 => "1111111010010000",
53977 => "1111111010010000",
53978 => "1111111010010000",
53979 => "1111111010010000",
53980 => "1111111010010000",
53981 => "1111111010010000",
53982 => "1111111010010001",
53983 => "1111111010010001",
53984 => "1111111010010001",
53985 => "1111111010010001",
53986 => "1111111010010001",
53987 => "1111111010010001",
53988 => "1111111010010001",
53989 => "1111111010010001",
53990 => "1111111010010001",
53991 => "1111111010010001",
53992 => "1111111010010001",
53993 => "1111111010010001",
53994 => "1111111010010010",
53995 => "1111111010010010",
53996 => "1111111010010010",
53997 => "1111111010010010",
53998 => "1111111010010010",
53999 => "1111111010010010",
54000 => "1111111010010010",
54001 => "1111111010010010",
54002 => "1111111010010010",
54003 => "1111111010010010",
54004 => "1111111010010010",
54005 => "1111111010010011",
54006 => "1111111010010011",
54007 => "1111111010010011",
54008 => "1111111010010011",
54009 => "1111111010010011",
54010 => "1111111010010011",
54011 => "1111111010010011",
54012 => "1111111010010011",
54013 => "1111111010010011",
54014 => "1111111010010011",
54015 => "1111111010010011",
54016 => "1111111010010100",
54017 => "1111111010010100",
54018 => "1111111010010100",
54019 => "1111111010010100",
54020 => "1111111010010100",
54021 => "1111111010010100",
54022 => "1111111010010100",
54023 => "1111111010010100",
54024 => "1111111010010100",
54025 => "1111111010010100",
54026 => "1111111010010100",
54027 => "1111111010010100",
54028 => "1111111010010101",
54029 => "1111111010010101",
54030 => "1111111010010101",
54031 => "1111111010010101",
54032 => "1111111010010101",
54033 => "1111111010010101",
54034 => "1111111010010101",
54035 => "1111111010010101",
54036 => "1111111010010101",
54037 => "1111111010010101",
54038 => "1111111010010101",
54039 => "1111111010010110",
54040 => "1111111010010110",
54041 => "1111111010010110",
54042 => "1111111010010110",
54043 => "1111111010010110",
54044 => "1111111010010110",
54045 => "1111111010010110",
54046 => "1111111010010110",
54047 => "1111111010010110",
54048 => "1111111010010110",
54049 => "1111111010010110",
54050 => "1111111010010111",
54051 => "1111111010010111",
54052 => "1111111010010111",
54053 => "1111111010010111",
54054 => "1111111010010111",
54055 => "1111111010010111",
54056 => "1111111010010111",
54057 => "1111111010010111",
54058 => "1111111010010111",
54059 => "1111111010010111",
54060 => "1111111010010111",
54061 => "1111111010010111",
54062 => "1111111010011000",
54063 => "1111111010011000",
54064 => "1111111010011000",
54065 => "1111111010011000",
54066 => "1111111010011000",
54067 => "1111111010011000",
54068 => "1111111010011000",
54069 => "1111111010011000",
54070 => "1111111010011000",
54071 => "1111111010011000",
54072 => "1111111010011000",
54073 => "1111111010011001",
54074 => "1111111010011001",
54075 => "1111111010011001",
54076 => "1111111010011001",
54077 => "1111111010011001",
54078 => "1111111010011001",
54079 => "1111111010011001",
54080 => "1111111010011001",
54081 => "1111111010011001",
54082 => "1111111010011001",
54083 => "1111111010011001",
54084 => "1111111010011001",
54085 => "1111111010011010",
54086 => "1111111010011010",
54087 => "1111111010011010",
54088 => "1111111010011010",
54089 => "1111111010011010",
54090 => "1111111010011010",
54091 => "1111111010011010",
54092 => "1111111010011010",
54093 => "1111111010011010",
54094 => "1111111010011010",
54095 => "1111111010011010",
54096 => "1111111010011011",
54097 => "1111111010011011",
54098 => "1111111010011011",
54099 => "1111111010011011",
54100 => "1111111010011011",
54101 => "1111111010011011",
54102 => "1111111010011011",
54103 => "1111111010011011",
54104 => "1111111010011011",
54105 => "1111111010011011",
54106 => "1111111010011011",
54107 => "1111111010011011",
54108 => "1111111010011100",
54109 => "1111111010011100",
54110 => "1111111010011100",
54111 => "1111111010011100",
54112 => "1111111010011100",
54113 => "1111111010011100",
54114 => "1111111010011100",
54115 => "1111111010011100",
54116 => "1111111010011100",
54117 => "1111111010011100",
54118 => "1111111010011100",
54119 => "1111111010011101",
54120 => "1111111010011101",
54121 => "1111111010011101",
54122 => "1111111010011101",
54123 => "1111111010011101",
54124 => "1111111010011101",
54125 => "1111111010011101",
54126 => "1111111010011101",
54127 => "1111111010011101",
54128 => "1111111010011101",
54129 => "1111111010011101",
54130 => "1111111010011101",
54131 => "1111111010011110",
54132 => "1111111010011110",
54133 => "1111111010011110",
54134 => "1111111010011110",
54135 => "1111111010011110",
54136 => "1111111010011110",
54137 => "1111111010011110",
54138 => "1111111010011110",
54139 => "1111111010011110",
54140 => "1111111010011110",
54141 => "1111111010011110",
54142 => "1111111010011110",
54143 => "1111111010011111",
54144 => "1111111010011111",
54145 => "1111111010011111",
54146 => "1111111010011111",
54147 => "1111111010011111",
54148 => "1111111010011111",
54149 => "1111111010011111",
54150 => "1111111010011111",
54151 => "1111111010011111",
54152 => "1111111010011111",
54153 => "1111111010011111",
54154 => "1111111010100000",
54155 => "1111111010100000",
54156 => "1111111010100000",
54157 => "1111111010100000",
54158 => "1111111010100000",
54159 => "1111111010100000",
54160 => "1111111010100000",
54161 => "1111111010100000",
54162 => "1111111010100000",
54163 => "1111111010100000",
54164 => "1111111010100000",
54165 => "1111111010100000",
54166 => "1111111010100001",
54167 => "1111111010100001",
54168 => "1111111010100001",
54169 => "1111111010100001",
54170 => "1111111010100001",
54171 => "1111111010100001",
54172 => "1111111010100001",
54173 => "1111111010100001",
54174 => "1111111010100001",
54175 => "1111111010100001",
54176 => "1111111010100001",
54177 => "1111111010100001",
54178 => "1111111010100010",
54179 => "1111111010100010",
54180 => "1111111010100010",
54181 => "1111111010100010",
54182 => "1111111010100010",
54183 => "1111111010100010",
54184 => "1111111010100010",
54185 => "1111111010100010",
54186 => "1111111010100010",
54187 => "1111111010100010",
54188 => "1111111010100010",
54189 => "1111111010100010",
54190 => "1111111010100011",
54191 => "1111111010100011",
54192 => "1111111010100011",
54193 => "1111111010100011",
54194 => "1111111010100011",
54195 => "1111111010100011",
54196 => "1111111010100011",
54197 => "1111111010100011",
54198 => "1111111010100011",
54199 => "1111111010100011",
54200 => "1111111010100011",
54201 => "1111111010100100",
54202 => "1111111010100100",
54203 => "1111111010100100",
54204 => "1111111010100100",
54205 => "1111111010100100",
54206 => "1111111010100100",
54207 => "1111111010100100",
54208 => "1111111010100100",
54209 => "1111111010100100",
54210 => "1111111010100100",
54211 => "1111111010100100",
54212 => "1111111010100100",
54213 => "1111111010100101",
54214 => "1111111010100101",
54215 => "1111111010100101",
54216 => "1111111010100101",
54217 => "1111111010100101",
54218 => "1111111010100101",
54219 => "1111111010100101",
54220 => "1111111010100101",
54221 => "1111111010100101",
54222 => "1111111010100101",
54223 => "1111111010100101",
54224 => "1111111010100101",
54225 => "1111111010100110",
54226 => "1111111010100110",
54227 => "1111111010100110",
54228 => "1111111010100110",
54229 => "1111111010100110",
54230 => "1111111010100110",
54231 => "1111111010100110",
54232 => "1111111010100110",
54233 => "1111111010100110",
54234 => "1111111010100110",
54235 => "1111111010100110",
54236 => "1111111010100110",
54237 => "1111111010100111",
54238 => "1111111010100111",
54239 => "1111111010100111",
54240 => "1111111010100111",
54241 => "1111111010100111",
54242 => "1111111010100111",
54243 => "1111111010100111",
54244 => "1111111010100111",
54245 => "1111111010100111",
54246 => "1111111010100111",
54247 => "1111111010100111",
54248 => "1111111010100111",
54249 => "1111111010101000",
54250 => "1111111010101000",
54251 => "1111111010101000",
54252 => "1111111010101000",
54253 => "1111111010101000",
54254 => "1111111010101000",
54255 => "1111111010101000",
54256 => "1111111010101000",
54257 => "1111111010101000",
54258 => "1111111010101000",
54259 => "1111111010101000",
54260 => "1111111010101000",
54261 => "1111111010101001",
54262 => "1111111010101001",
54263 => "1111111010101001",
54264 => "1111111010101001",
54265 => "1111111010101001",
54266 => "1111111010101001",
54267 => "1111111010101001",
54268 => "1111111010101001",
54269 => "1111111010101001",
54270 => "1111111010101001",
54271 => "1111111010101001",
54272 => "1111111010101001",
54273 => "1111111010101010",
54274 => "1111111010101010",
54275 => "1111111010101010",
54276 => "1111111010101010",
54277 => "1111111010101010",
54278 => "1111111010101010",
54279 => "1111111010101010",
54280 => "1111111010101010",
54281 => "1111111010101010",
54282 => "1111111010101010",
54283 => "1111111010101010",
54284 => "1111111010101010",
54285 => "1111111010101011",
54286 => "1111111010101011",
54287 => "1111111010101011",
54288 => "1111111010101011",
54289 => "1111111010101011",
54290 => "1111111010101011",
54291 => "1111111010101011",
54292 => "1111111010101011",
54293 => "1111111010101011",
54294 => "1111111010101011",
54295 => "1111111010101011",
54296 => "1111111010101011",
54297 => "1111111010101100",
54298 => "1111111010101100",
54299 => "1111111010101100",
54300 => "1111111010101100",
54301 => "1111111010101100",
54302 => "1111111010101100",
54303 => "1111111010101100",
54304 => "1111111010101100",
54305 => "1111111010101100",
54306 => "1111111010101100",
54307 => "1111111010101100",
54308 => "1111111010101100",
54309 => "1111111010101101",
54310 => "1111111010101101",
54311 => "1111111010101101",
54312 => "1111111010101101",
54313 => "1111111010101101",
54314 => "1111111010101101",
54315 => "1111111010101101",
54316 => "1111111010101101",
54317 => "1111111010101101",
54318 => "1111111010101101",
54319 => "1111111010101101",
54320 => "1111111010101101",
54321 => "1111111010101110",
54322 => "1111111010101110",
54323 => "1111111010101110",
54324 => "1111111010101110",
54325 => "1111111010101110",
54326 => "1111111010101110",
54327 => "1111111010101110",
54328 => "1111111010101110",
54329 => "1111111010101110",
54330 => "1111111010101110",
54331 => "1111111010101110",
54332 => "1111111010101110",
54333 => "1111111010101110",
54334 => "1111111010101111",
54335 => "1111111010101111",
54336 => "1111111010101111",
54337 => "1111111010101111",
54338 => "1111111010101111",
54339 => "1111111010101111",
54340 => "1111111010101111",
54341 => "1111111010101111",
54342 => "1111111010101111",
54343 => "1111111010101111",
54344 => "1111111010101111",
54345 => "1111111010101111",
54346 => "1111111010110000",
54347 => "1111111010110000",
54348 => "1111111010110000",
54349 => "1111111010110000",
54350 => "1111111010110000",
54351 => "1111111010110000",
54352 => "1111111010110000",
54353 => "1111111010110000",
54354 => "1111111010110000",
54355 => "1111111010110000",
54356 => "1111111010110000",
54357 => "1111111010110000",
54358 => "1111111010110001",
54359 => "1111111010110001",
54360 => "1111111010110001",
54361 => "1111111010110001",
54362 => "1111111010110001",
54363 => "1111111010110001",
54364 => "1111111010110001",
54365 => "1111111010110001",
54366 => "1111111010110001",
54367 => "1111111010110001",
54368 => "1111111010110001",
54369 => "1111111010110001",
54370 => "1111111010110010",
54371 => "1111111010110010",
54372 => "1111111010110010",
54373 => "1111111010110010",
54374 => "1111111010110010",
54375 => "1111111010110010",
54376 => "1111111010110010",
54377 => "1111111010110010",
54378 => "1111111010110010",
54379 => "1111111010110010",
54380 => "1111111010110010",
54381 => "1111111010110010",
54382 => "1111111010110010",
54383 => "1111111010110011",
54384 => "1111111010110011",
54385 => "1111111010110011",
54386 => "1111111010110011",
54387 => "1111111010110011",
54388 => "1111111010110011",
54389 => "1111111010110011",
54390 => "1111111010110011",
54391 => "1111111010110011",
54392 => "1111111010110011",
54393 => "1111111010110011",
54394 => "1111111010110011",
54395 => "1111111010110100",
54396 => "1111111010110100",
54397 => "1111111010110100",
54398 => "1111111010110100",
54399 => "1111111010110100",
54400 => "1111111010110100",
54401 => "1111111010110100",
54402 => "1111111010110100",
54403 => "1111111010110100",
54404 => "1111111010110100",
54405 => "1111111010110100",
54406 => "1111111010110100",
54407 => "1111111010110100",
54408 => "1111111010110101",
54409 => "1111111010110101",
54410 => "1111111010110101",
54411 => "1111111010110101",
54412 => "1111111010110101",
54413 => "1111111010110101",
54414 => "1111111010110101",
54415 => "1111111010110101",
54416 => "1111111010110101",
54417 => "1111111010110101",
54418 => "1111111010110101",
54419 => "1111111010110101",
54420 => "1111111010110110",
54421 => "1111111010110110",
54422 => "1111111010110110",
54423 => "1111111010110110",
54424 => "1111111010110110",
54425 => "1111111010110110",
54426 => "1111111010110110",
54427 => "1111111010110110",
54428 => "1111111010110110",
54429 => "1111111010110110",
54430 => "1111111010110110",
54431 => "1111111010110110",
54432 => "1111111010110111",
54433 => "1111111010110111",
54434 => "1111111010110111",
54435 => "1111111010110111",
54436 => "1111111010110111",
54437 => "1111111010110111",
54438 => "1111111010110111",
54439 => "1111111010110111",
54440 => "1111111010110111",
54441 => "1111111010110111",
54442 => "1111111010110111",
54443 => "1111111010110111",
54444 => "1111111010110111",
54445 => "1111111010111000",
54446 => "1111111010111000",
54447 => "1111111010111000",
54448 => "1111111010111000",
54449 => "1111111010111000",
54450 => "1111111010111000",
54451 => "1111111010111000",
54452 => "1111111010111000",
54453 => "1111111010111000",
54454 => "1111111010111000",
54455 => "1111111010111000",
54456 => "1111111010111000",
54457 => "1111111010111000",
54458 => "1111111010111001",
54459 => "1111111010111001",
54460 => "1111111010111001",
54461 => "1111111010111001",
54462 => "1111111010111001",
54463 => "1111111010111001",
54464 => "1111111010111001",
54465 => "1111111010111001",
54466 => "1111111010111001",
54467 => "1111111010111001",
54468 => "1111111010111001",
54469 => "1111111010111001",
54470 => "1111111010111010",
54471 => "1111111010111010",
54472 => "1111111010111010",
54473 => "1111111010111010",
54474 => "1111111010111010",
54475 => "1111111010111010",
54476 => "1111111010111010",
54477 => "1111111010111010",
54478 => "1111111010111010",
54479 => "1111111010111010",
54480 => "1111111010111010",
54481 => "1111111010111010",
54482 => "1111111010111010",
54483 => "1111111010111011",
54484 => "1111111010111011",
54485 => "1111111010111011",
54486 => "1111111010111011",
54487 => "1111111010111011",
54488 => "1111111010111011",
54489 => "1111111010111011",
54490 => "1111111010111011",
54491 => "1111111010111011",
54492 => "1111111010111011",
54493 => "1111111010111011",
54494 => "1111111010111011",
54495 => "1111111010111011",
54496 => "1111111010111100",
54497 => "1111111010111100",
54498 => "1111111010111100",
54499 => "1111111010111100",
54500 => "1111111010111100",
54501 => "1111111010111100",
54502 => "1111111010111100",
54503 => "1111111010111100",
54504 => "1111111010111100",
54505 => "1111111010111100",
54506 => "1111111010111100",
54507 => "1111111010111100",
54508 => "1111111010111101",
54509 => "1111111010111101",
54510 => "1111111010111101",
54511 => "1111111010111101",
54512 => "1111111010111101",
54513 => "1111111010111101",
54514 => "1111111010111101",
54515 => "1111111010111101",
54516 => "1111111010111101",
54517 => "1111111010111101",
54518 => "1111111010111101",
54519 => "1111111010111101",
54520 => "1111111010111101",
54521 => "1111111010111110",
54522 => "1111111010111110",
54523 => "1111111010111110",
54524 => "1111111010111110",
54525 => "1111111010111110",
54526 => "1111111010111110",
54527 => "1111111010111110",
54528 => "1111111010111110",
54529 => "1111111010111110",
54530 => "1111111010111110",
54531 => "1111111010111110",
54532 => "1111111010111110",
54533 => "1111111010111110",
54534 => "1111111010111111",
54535 => "1111111010111111",
54536 => "1111111010111111",
54537 => "1111111010111111",
54538 => "1111111010111111",
54539 => "1111111010111111",
54540 => "1111111010111111",
54541 => "1111111010111111",
54542 => "1111111010111111",
54543 => "1111111010111111",
54544 => "1111111010111111",
54545 => "1111111010111111",
54546 => "1111111010111111",
54547 => "1111111011000000",
54548 => "1111111011000000",
54549 => "1111111011000000",
54550 => "1111111011000000",
54551 => "1111111011000000",
54552 => "1111111011000000",
54553 => "1111111011000000",
54554 => "1111111011000000",
54555 => "1111111011000000",
54556 => "1111111011000000",
54557 => "1111111011000000",
54558 => "1111111011000000",
54559 => "1111111011000000",
54560 => "1111111011000001",
54561 => "1111111011000001",
54562 => "1111111011000001",
54563 => "1111111011000001",
54564 => "1111111011000001",
54565 => "1111111011000001",
54566 => "1111111011000001",
54567 => "1111111011000001",
54568 => "1111111011000001",
54569 => "1111111011000001",
54570 => "1111111011000001",
54571 => "1111111011000001",
54572 => "1111111011000010",
54573 => "1111111011000010",
54574 => "1111111011000010",
54575 => "1111111011000010",
54576 => "1111111011000010",
54577 => "1111111011000010",
54578 => "1111111011000010",
54579 => "1111111011000010",
54580 => "1111111011000010",
54581 => "1111111011000010",
54582 => "1111111011000010",
54583 => "1111111011000010",
54584 => "1111111011000010",
54585 => "1111111011000011",
54586 => "1111111011000011",
54587 => "1111111011000011",
54588 => "1111111011000011",
54589 => "1111111011000011",
54590 => "1111111011000011",
54591 => "1111111011000011",
54592 => "1111111011000011",
54593 => "1111111011000011",
54594 => "1111111011000011",
54595 => "1111111011000011",
54596 => "1111111011000011",
54597 => "1111111011000011",
54598 => "1111111011000100",
54599 => "1111111011000100",
54600 => "1111111011000100",
54601 => "1111111011000100",
54602 => "1111111011000100",
54603 => "1111111011000100",
54604 => "1111111011000100",
54605 => "1111111011000100",
54606 => "1111111011000100",
54607 => "1111111011000100",
54608 => "1111111011000100",
54609 => "1111111011000100",
54610 => "1111111011000100",
54611 => "1111111011000101",
54612 => "1111111011000101",
54613 => "1111111011000101",
54614 => "1111111011000101",
54615 => "1111111011000101",
54616 => "1111111011000101",
54617 => "1111111011000101",
54618 => "1111111011000101",
54619 => "1111111011000101",
54620 => "1111111011000101",
54621 => "1111111011000101",
54622 => "1111111011000101",
54623 => "1111111011000101",
54624 => "1111111011000101",
54625 => "1111111011000110",
54626 => "1111111011000110",
54627 => "1111111011000110",
54628 => "1111111011000110",
54629 => "1111111011000110",
54630 => "1111111011000110",
54631 => "1111111011000110",
54632 => "1111111011000110",
54633 => "1111111011000110",
54634 => "1111111011000110",
54635 => "1111111011000110",
54636 => "1111111011000110",
54637 => "1111111011000110",
54638 => "1111111011000111",
54639 => "1111111011000111",
54640 => "1111111011000111",
54641 => "1111111011000111",
54642 => "1111111011000111",
54643 => "1111111011000111",
54644 => "1111111011000111",
54645 => "1111111011000111",
54646 => "1111111011000111",
54647 => "1111111011000111",
54648 => "1111111011000111",
54649 => "1111111011000111",
54650 => "1111111011000111",
54651 => "1111111011001000",
54652 => "1111111011001000",
54653 => "1111111011001000",
54654 => "1111111011001000",
54655 => "1111111011001000",
54656 => "1111111011001000",
54657 => "1111111011001000",
54658 => "1111111011001000",
54659 => "1111111011001000",
54660 => "1111111011001000",
54661 => "1111111011001000",
54662 => "1111111011001000",
54663 => "1111111011001000",
54664 => "1111111011001001",
54665 => "1111111011001001",
54666 => "1111111011001001",
54667 => "1111111011001001",
54668 => "1111111011001001",
54669 => "1111111011001001",
54670 => "1111111011001001",
54671 => "1111111011001001",
54672 => "1111111011001001",
54673 => "1111111011001001",
54674 => "1111111011001001",
54675 => "1111111011001001",
54676 => "1111111011001001",
54677 => "1111111011001010",
54678 => "1111111011001010",
54679 => "1111111011001010",
54680 => "1111111011001010",
54681 => "1111111011001010",
54682 => "1111111011001010",
54683 => "1111111011001010",
54684 => "1111111011001010",
54685 => "1111111011001010",
54686 => "1111111011001010",
54687 => "1111111011001010",
54688 => "1111111011001010",
54689 => "1111111011001010",
54690 => "1111111011001010",
54691 => "1111111011001011",
54692 => "1111111011001011",
54693 => "1111111011001011",
54694 => "1111111011001011",
54695 => "1111111011001011",
54696 => "1111111011001011",
54697 => "1111111011001011",
54698 => "1111111011001011",
54699 => "1111111011001011",
54700 => "1111111011001011",
54701 => "1111111011001011",
54702 => "1111111011001011",
54703 => "1111111011001011",
54704 => "1111111011001100",
54705 => "1111111011001100",
54706 => "1111111011001100",
54707 => "1111111011001100",
54708 => "1111111011001100",
54709 => "1111111011001100",
54710 => "1111111011001100",
54711 => "1111111011001100",
54712 => "1111111011001100",
54713 => "1111111011001100",
54714 => "1111111011001100",
54715 => "1111111011001100",
54716 => "1111111011001100",
54717 => "1111111011001101",
54718 => "1111111011001101",
54719 => "1111111011001101",
54720 => "1111111011001101",
54721 => "1111111011001101",
54722 => "1111111011001101",
54723 => "1111111011001101",
54724 => "1111111011001101",
54725 => "1111111011001101",
54726 => "1111111011001101",
54727 => "1111111011001101",
54728 => "1111111011001101",
54729 => "1111111011001101",
54730 => "1111111011001101",
54731 => "1111111011001110",
54732 => "1111111011001110",
54733 => "1111111011001110",
54734 => "1111111011001110",
54735 => "1111111011001110",
54736 => "1111111011001110",
54737 => "1111111011001110",
54738 => "1111111011001110",
54739 => "1111111011001110",
54740 => "1111111011001110",
54741 => "1111111011001110",
54742 => "1111111011001110",
54743 => "1111111011001110",
54744 => "1111111011001111",
54745 => "1111111011001111",
54746 => "1111111011001111",
54747 => "1111111011001111",
54748 => "1111111011001111",
54749 => "1111111011001111",
54750 => "1111111011001111",
54751 => "1111111011001111",
54752 => "1111111011001111",
54753 => "1111111011001111",
54754 => "1111111011001111",
54755 => "1111111011001111",
54756 => "1111111011001111",
54757 => "1111111011001111",
54758 => "1111111011010000",
54759 => "1111111011010000",
54760 => "1111111011010000",
54761 => "1111111011010000",
54762 => "1111111011010000",
54763 => "1111111011010000",
54764 => "1111111011010000",
54765 => "1111111011010000",
54766 => "1111111011010000",
54767 => "1111111011010000",
54768 => "1111111011010000",
54769 => "1111111011010000",
54770 => "1111111011010000",
54771 => "1111111011010001",
54772 => "1111111011010001",
54773 => "1111111011010001",
54774 => "1111111011010001",
54775 => "1111111011010001",
54776 => "1111111011010001",
54777 => "1111111011010001",
54778 => "1111111011010001",
54779 => "1111111011010001",
54780 => "1111111011010001",
54781 => "1111111011010001",
54782 => "1111111011010001",
54783 => "1111111011010001",
54784 => "1111111011010001",
54785 => "1111111011010010",
54786 => "1111111011010010",
54787 => "1111111011010010",
54788 => "1111111011010010",
54789 => "1111111011010010",
54790 => "1111111011010010",
54791 => "1111111011010010",
54792 => "1111111011010010",
54793 => "1111111011010010",
54794 => "1111111011010010",
54795 => "1111111011010010",
54796 => "1111111011010010",
54797 => "1111111011010010",
54798 => "1111111011010010",
54799 => "1111111011010011",
54800 => "1111111011010011",
54801 => "1111111011010011",
54802 => "1111111011010011",
54803 => "1111111011010011",
54804 => "1111111011010011",
54805 => "1111111011010011",
54806 => "1111111011010011",
54807 => "1111111011010011",
54808 => "1111111011010011",
54809 => "1111111011010011",
54810 => "1111111011010011",
54811 => "1111111011010011",
54812 => "1111111011010100",
54813 => "1111111011010100",
54814 => "1111111011010100",
54815 => "1111111011010100",
54816 => "1111111011010100",
54817 => "1111111011010100",
54818 => "1111111011010100",
54819 => "1111111011010100",
54820 => "1111111011010100",
54821 => "1111111011010100",
54822 => "1111111011010100",
54823 => "1111111011010100",
54824 => "1111111011010100",
54825 => "1111111011010100",
54826 => "1111111011010101",
54827 => "1111111011010101",
54828 => "1111111011010101",
54829 => "1111111011010101",
54830 => "1111111011010101",
54831 => "1111111011010101",
54832 => "1111111011010101",
54833 => "1111111011010101",
54834 => "1111111011010101",
54835 => "1111111011010101",
54836 => "1111111011010101",
54837 => "1111111011010101",
54838 => "1111111011010101",
54839 => "1111111011010101",
54840 => "1111111011010110",
54841 => "1111111011010110",
54842 => "1111111011010110",
54843 => "1111111011010110",
54844 => "1111111011010110",
54845 => "1111111011010110",
54846 => "1111111011010110",
54847 => "1111111011010110",
54848 => "1111111011010110",
54849 => "1111111011010110",
54850 => "1111111011010110",
54851 => "1111111011010110",
54852 => "1111111011010110",
54853 => "1111111011010110",
54854 => "1111111011010111",
54855 => "1111111011010111",
54856 => "1111111011010111",
54857 => "1111111011010111",
54858 => "1111111011010111",
54859 => "1111111011010111",
54860 => "1111111011010111",
54861 => "1111111011010111",
54862 => "1111111011010111",
54863 => "1111111011010111",
54864 => "1111111011010111",
54865 => "1111111011010111",
54866 => "1111111011010111",
54867 => "1111111011010111",
54868 => "1111111011011000",
54869 => "1111111011011000",
54870 => "1111111011011000",
54871 => "1111111011011000",
54872 => "1111111011011000",
54873 => "1111111011011000",
54874 => "1111111011011000",
54875 => "1111111011011000",
54876 => "1111111011011000",
54877 => "1111111011011000",
54878 => "1111111011011000",
54879 => "1111111011011000",
54880 => "1111111011011000",
54881 => "1111111011011001",
54882 => "1111111011011001",
54883 => "1111111011011001",
54884 => "1111111011011001",
54885 => "1111111011011001",
54886 => "1111111011011001",
54887 => "1111111011011001",
54888 => "1111111011011001",
54889 => "1111111011011001",
54890 => "1111111011011001",
54891 => "1111111011011001",
54892 => "1111111011011001",
54893 => "1111111011011001",
54894 => "1111111011011001",
54895 => "1111111011011010",
54896 => "1111111011011010",
54897 => "1111111011011010",
54898 => "1111111011011010",
54899 => "1111111011011010",
54900 => "1111111011011010",
54901 => "1111111011011010",
54902 => "1111111011011010",
54903 => "1111111011011010",
54904 => "1111111011011010",
54905 => "1111111011011010",
54906 => "1111111011011010",
54907 => "1111111011011010",
54908 => "1111111011011010",
54909 => "1111111011011011",
54910 => "1111111011011011",
54911 => "1111111011011011",
54912 => "1111111011011011",
54913 => "1111111011011011",
54914 => "1111111011011011",
54915 => "1111111011011011",
54916 => "1111111011011011",
54917 => "1111111011011011",
54918 => "1111111011011011",
54919 => "1111111011011011",
54920 => "1111111011011011",
54921 => "1111111011011011",
54922 => "1111111011011011",
54923 => "1111111011011100",
54924 => "1111111011011100",
54925 => "1111111011011100",
54926 => "1111111011011100",
54927 => "1111111011011100",
54928 => "1111111011011100",
54929 => "1111111011011100",
54930 => "1111111011011100",
54931 => "1111111011011100",
54932 => "1111111011011100",
54933 => "1111111011011100",
54934 => "1111111011011100",
54935 => "1111111011011100",
54936 => "1111111011011100",
54937 => "1111111011011100",
54938 => "1111111011011101",
54939 => "1111111011011101",
54940 => "1111111011011101",
54941 => "1111111011011101",
54942 => "1111111011011101",
54943 => "1111111011011101",
54944 => "1111111011011101",
54945 => "1111111011011101",
54946 => "1111111011011101",
54947 => "1111111011011101",
54948 => "1111111011011101",
54949 => "1111111011011101",
54950 => "1111111011011101",
54951 => "1111111011011101",
54952 => "1111111011011110",
54953 => "1111111011011110",
54954 => "1111111011011110",
54955 => "1111111011011110",
54956 => "1111111011011110",
54957 => "1111111011011110",
54958 => "1111111011011110",
54959 => "1111111011011110",
54960 => "1111111011011110",
54961 => "1111111011011110",
54962 => "1111111011011110",
54963 => "1111111011011110",
54964 => "1111111011011110",
54965 => "1111111011011110",
54966 => "1111111011011111",
54967 => "1111111011011111",
54968 => "1111111011011111",
54969 => "1111111011011111",
54970 => "1111111011011111",
54971 => "1111111011011111",
54972 => "1111111011011111",
54973 => "1111111011011111",
54974 => "1111111011011111",
54975 => "1111111011011111",
54976 => "1111111011011111",
54977 => "1111111011011111",
54978 => "1111111011011111",
54979 => "1111111011011111",
54980 => "1111111011100000",
54981 => "1111111011100000",
54982 => "1111111011100000",
54983 => "1111111011100000",
54984 => "1111111011100000",
54985 => "1111111011100000",
54986 => "1111111011100000",
54987 => "1111111011100000",
54988 => "1111111011100000",
54989 => "1111111011100000",
54990 => "1111111011100000",
54991 => "1111111011100000",
54992 => "1111111011100000",
54993 => "1111111011100000",
54994 => "1111111011100000",
54995 => "1111111011100001",
54996 => "1111111011100001",
54997 => "1111111011100001",
54998 => "1111111011100001",
54999 => "1111111011100001",
55000 => "1111111011100001",
55001 => "1111111011100001",
55002 => "1111111011100001",
55003 => "1111111011100001",
55004 => "1111111011100001",
55005 => "1111111011100001",
55006 => "1111111011100001",
55007 => "1111111011100001",
55008 => "1111111011100001",
55009 => "1111111011100010",
55010 => "1111111011100010",
55011 => "1111111011100010",
55012 => "1111111011100010",
55013 => "1111111011100010",
55014 => "1111111011100010",
55015 => "1111111011100010",
55016 => "1111111011100010",
55017 => "1111111011100010",
55018 => "1111111011100010",
55019 => "1111111011100010",
55020 => "1111111011100010",
55021 => "1111111011100010",
55022 => "1111111011100010",
55023 => "1111111011100011",
55024 => "1111111011100011",
55025 => "1111111011100011",
55026 => "1111111011100011",
55027 => "1111111011100011",
55028 => "1111111011100011",
55029 => "1111111011100011",
55030 => "1111111011100011",
55031 => "1111111011100011",
55032 => "1111111011100011",
55033 => "1111111011100011",
55034 => "1111111011100011",
55035 => "1111111011100011",
55036 => "1111111011100011",
55037 => "1111111011100011",
55038 => "1111111011100100",
55039 => "1111111011100100",
55040 => "1111111011100100",
55041 => "1111111011100100",
55042 => "1111111011100100",
55043 => "1111111011100100",
55044 => "1111111011100100",
55045 => "1111111011100100",
55046 => "1111111011100100",
55047 => "1111111011100100",
55048 => "1111111011100100",
55049 => "1111111011100100",
55050 => "1111111011100100",
55051 => "1111111011100100",
55052 => "1111111011100101",
55053 => "1111111011100101",
55054 => "1111111011100101",
55055 => "1111111011100101",
55056 => "1111111011100101",
55057 => "1111111011100101",
55058 => "1111111011100101",
55059 => "1111111011100101",
55060 => "1111111011100101",
55061 => "1111111011100101",
55062 => "1111111011100101",
55063 => "1111111011100101",
55064 => "1111111011100101",
55065 => "1111111011100101",
55066 => "1111111011100101",
55067 => "1111111011100110",
55068 => "1111111011100110",
55069 => "1111111011100110",
55070 => "1111111011100110",
55071 => "1111111011100110",
55072 => "1111111011100110",
55073 => "1111111011100110",
55074 => "1111111011100110",
55075 => "1111111011100110",
55076 => "1111111011100110",
55077 => "1111111011100110",
55078 => "1111111011100110",
55079 => "1111111011100110",
55080 => "1111111011100110",
55081 => "1111111011100111",
55082 => "1111111011100111",
55083 => "1111111011100111",
55084 => "1111111011100111",
55085 => "1111111011100111",
55086 => "1111111011100111",
55087 => "1111111011100111",
55088 => "1111111011100111",
55089 => "1111111011100111",
55090 => "1111111011100111",
55091 => "1111111011100111",
55092 => "1111111011100111",
55093 => "1111111011100111",
55094 => "1111111011100111",
55095 => "1111111011100111",
55096 => "1111111011101000",
55097 => "1111111011101000",
55098 => "1111111011101000",
55099 => "1111111011101000",
55100 => "1111111011101000",
55101 => "1111111011101000",
55102 => "1111111011101000",
55103 => "1111111011101000",
55104 => "1111111011101000",
55105 => "1111111011101000",
55106 => "1111111011101000",
55107 => "1111111011101000",
55108 => "1111111011101000",
55109 => "1111111011101000",
55110 => "1111111011101000",
55111 => "1111111011101001",
55112 => "1111111011101001",
55113 => "1111111011101001",
55114 => "1111111011101001",
55115 => "1111111011101001",
55116 => "1111111011101001",
55117 => "1111111011101001",
55118 => "1111111011101001",
55119 => "1111111011101001",
55120 => "1111111011101001",
55121 => "1111111011101001",
55122 => "1111111011101001",
55123 => "1111111011101001",
55124 => "1111111011101001",
55125 => "1111111011101001",
55126 => "1111111011101010",
55127 => "1111111011101010",
55128 => "1111111011101010",
55129 => "1111111011101010",
55130 => "1111111011101010",
55131 => "1111111011101010",
55132 => "1111111011101010",
55133 => "1111111011101010",
55134 => "1111111011101010",
55135 => "1111111011101010",
55136 => "1111111011101010",
55137 => "1111111011101010",
55138 => "1111111011101010",
55139 => "1111111011101010",
55140 => "1111111011101011",
55141 => "1111111011101011",
55142 => "1111111011101011",
55143 => "1111111011101011",
55144 => "1111111011101011",
55145 => "1111111011101011",
55146 => "1111111011101011",
55147 => "1111111011101011",
55148 => "1111111011101011",
55149 => "1111111011101011",
55150 => "1111111011101011",
55151 => "1111111011101011",
55152 => "1111111011101011",
55153 => "1111111011101011",
55154 => "1111111011101011",
55155 => "1111111011101100",
55156 => "1111111011101100",
55157 => "1111111011101100",
55158 => "1111111011101100",
55159 => "1111111011101100",
55160 => "1111111011101100",
55161 => "1111111011101100",
55162 => "1111111011101100",
55163 => "1111111011101100",
55164 => "1111111011101100",
55165 => "1111111011101100",
55166 => "1111111011101100",
55167 => "1111111011101100",
55168 => "1111111011101100",
55169 => "1111111011101100",
55170 => "1111111011101101",
55171 => "1111111011101101",
55172 => "1111111011101101",
55173 => "1111111011101101",
55174 => "1111111011101101",
55175 => "1111111011101101",
55176 => "1111111011101101",
55177 => "1111111011101101",
55178 => "1111111011101101",
55179 => "1111111011101101",
55180 => "1111111011101101",
55181 => "1111111011101101",
55182 => "1111111011101101",
55183 => "1111111011101101",
55184 => "1111111011101101",
55185 => "1111111011101110",
55186 => "1111111011101110",
55187 => "1111111011101110",
55188 => "1111111011101110",
55189 => "1111111011101110",
55190 => "1111111011101110",
55191 => "1111111011101110",
55192 => "1111111011101110",
55193 => "1111111011101110",
55194 => "1111111011101110",
55195 => "1111111011101110",
55196 => "1111111011101110",
55197 => "1111111011101110",
55198 => "1111111011101110",
55199 => "1111111011101110",
55200 => "1111111011101111",
55201 => "1111111011101111",
55202 => "1111111011101111",
55203 => "1111111011101111",
55204 => "1111111011101111",
55205 => "1111111011101111",
55206 => "1111111011101111",
55207 => "1111111011101111",
55208 => "1111111011101111",
55209 => "1111111011101111",
55210 => "1111111011101111",
55211 => "1111111011101111",
55212 => "1111111011101111",
55213 => "1111111011101111",
55214 => "1111111011101111",
55215 => "1111111011110000",
55216 => "1111111011110000",
55217 => "1111111011110000",
55218 => "1111111011110000",
55219 => "1111111011110000",
55220 => "1111111011110000",
55221 => "1111111011110000",
55222 => "1111111011110000",
55223 => "1111111011110000",
55224 => "1111111011110000",
55225 => "1111111011110000",
55226 => "1111111011110000",
55227 => "1111111011110000",
55228 => "1111111011110000",
55229 => "1111111011110000",
55230 => "1111111011110001",
55231 => "1111111011110001",
55232 => "1111111011110001",
55233 => "1111111011110001",
55234 => "1111111011110001",
55235 => "1111111011110001",
55236 => "1111111011110001",
55237 => "1111111011110001",
55238 => "1111111011110001",
55239 => "1111111011110001",
55240 => "1111111011110001",
55241 => "1111111011110001",
55242 => "1111111011110001",
55243 => "1111111011110001",
55244 => "1111111011110001",
55245 => "1111111011110001",
55246 => "1111111011110010",
55247 => "1111111011110010",
55248 => "1111111011110010",
55249 => "1111111011110010",
55250 => "1111111011110010",
55251 => "1111111011110010",
55252 => "1111111011110010",
55253 => "1111111011110010",
55254 => "1111111011110010",
55255 => "1111111011110010",
55256 => "1111111011110010",
55257 => "1111111011110010",
55258 => "1111111011110010",
55259 => "1111111011110010",
55260 => "1111111011110010",
55261 => "1111111011110011",
55262 => "1111111011110011",
55263 => "1111111011110011",
55264 => "1111111011110011",
55265 => "1111111011110011",
55266 => "1111111011110011",
55267 => "1111111011110011",
55268 => "1111111011110011",
55269 => "1111111011110011",
55270 => "1111111011110011",
55271 => "1111111011110011",
55272 => "1111111011110011",
55273 => "1111111011110011",
55274 => "1111111011110011",
55275 => "1111111011110011",
55276 => "1111111011110100",
55277 => "1111111011110100",
55278 => "1111111011110100",
55279 => "1111111011110100",
55280 => "1111111011110100",
55281 => "1111111011110100",
55282 => "1111111011110100",
55283 => "1111111011110100",
55284 => "1111111011110100",
55285 => "1111111011110100",
55286 => "1111111011110100",
55287 => "1111111011110100",
55288 => "1111111011110100",
55289 => "1111111011110100",
55290 => "1111111011110100",
55291 => "1111111011110100",
55292 => "1111111011110101",
55293 => "1111111011110101",
55294 => "1111111011110101",
55295 => "1111111011110101",
55296 => "1111111011110101",
55297 => "1111111011110101",
55298 => "1111111011110101",
55299 => "1111111011110101",
55300 => "1111111011110101",
55301 => "1111111011110101",
55302 => "1111111011110101",
55303 => "1111111011110101",
55304 => "1111111011110101",
55305 => "1111111011110101",
55306 => "1111111011110101",
55307 => "1111111011110110",
55308 => "1111111011110110",
55309 => "1111111011110110",
55310 => "1111111011110110",
55311 => "1111111011110110",
55312 => "1111111011110110",
55313 => "1111111011110110",
55314 => "1111111011110110",
55315 => "1111111011110110",
55316 => "1111111011110110",
55317 => "1111111011110110",
55318 => "1111111011110110",
55319 => "1111111011110110",
55320 => "1111111011110110",
55321 => "1111111011110110",
55322 => "1111111011110110",
55323 => "1111111011110111",
55324 => "1111111011110111",
55325 => "1111111011110111",
55326 => "1111111011110111",
55327 => "1111111011110111",
55328 => "1111111011110111",
55329 => "1111111011110111",
55330 => "1111111011110111",
55331 => "1111111011110111",
55332 => "1111111011110111",
55333 => "1111111011110111",
55334 => "1111111011110111",
55335 => "1111111011110111",
55336 => "1111111011110111",
55337 => "1111111011110111",
55338 => "1111111011111000",
55339 => "1111111011111000",
55340 => "1111111011111000",
55341 => "1111111011111000",
55342 => "1111111011111000",
55343 => "1111111011111000",
55344 => "1111111011111000",
55345 => "1111111011111000",
55346 => "1111111011111000",
55347 => "1111111011111000",
55348 => "1111111011111000",
55349 => "1111111011111000",
55350 => "1111111011111000",
55351 => "1111111011111000",
55352 => "1111111011111000",
55353 => "1111111011111000",
55354 => "1111111011111001",
55355 => "1111111011111001",
55356 => "1111111011111001",
55357 => "1111111011111001",
55358 => "1111111011111001",
55359 => "1111111011111001",
55360 => "1111111011111001",
55361 => "1111111011111001",
55362 => "1111111011111001",
55363 => "1111111011111001",
55364 => "1111111011111001",
55365 => "1111111011111001",
55366 => "1111111011111001",
55367 => "1111111011111001",
55368 => "1111111011111001",
55369 => "1111111011111010",
55370 => "1111111011111010",
55371 => "1111111011111010",
55372 => "1111111011111010",
55373 => "1111111011111010",
55374 => "1111111011111010",
55375 => "1111111011111010",
55376 => "1111111011111010",
55377 => "1111111011111010",
55378 => "1111111011111010",
55379 => "1111111011111010",
55380 => "1111111011111010",
55381 => "1111111011111010",
55382 => "1111111011111010",
55383 => "1111111011111010",
55384 => "1111111011111010",
55385 => "1111111011111011",
55386 => "1111111011111011",
55387 => "1111111011111011",
55388 => "1111111011111011",
55389 => "1111111011111011",
55390 => "1111111011111011",
55391 => "1111111011111011",
55392 => "1111111011111011",
55393 => "1111111011111011",
55394 => "1111111011111011",
55395 => "1111111011111011",
55396 => "1111111011111011",
55397 => "1111111011111011",
55398 => "1111111011111011",
55399 => "1111111011111011",
55400 => "1111111011111011",
55401 => "1111111011111100",
55402 => "1111111011111100",
55403 => "1111111011111100",
55404 => "1111111011111100",
55405 => "1111111011111100",
55406 => "1111111011111100",
55407 => "1111111011111100",
55408 => "1111111011111100",
55409 => "1111111011111100",
55410 => "1111111011111100",
55411 => "1111111011111100",
55412 => "1111111011111100",
55413 => "1111111011111100",
55414 => "1111111011111100",
55415 => "1111111011111100",
55416 => "1111111011111100",
55417 => "1111111011111101",
55418 => "1111111011111101",
55419 => "1111111011111101",
55420 => "1111111011111101",
55421 => "1111111011111101",
55422 => "1111111011111101",
55423 => "1111111011111101",
55424 => "1111111011111101",
55425 => "1111111011111101",
55426 => "1111111011111101",
55427 => "1111111011111101",
55428 => "1111111011111101",
55429 => "1111111011111101",
55430 => "1111111011111101",
55431 => "1111111011111101",
55432 => "1111111011111101",
55433 => "1111111011111110",
55434 => "1111111011111110",
55435 => "1111111011111110",
55436 => "1111111011111110",
55437 => "1111111011111110",
55438 => "1111111011111110",
55439 => "1111111011111110",
55440 => "1111111011111110",
55441 => "1111111011111110",
55442 => "1111111011111110",
55443 => "1111111011111110",
55444 => "1111111011111110",
55445 => "1111111011111110",
55446 => "1111111011111110",
55447 => "1111111011111110",
55448 => "1111111011111110",
55449 => "1111111011111111",
55450 => "1111111011111111",
55451 => "1111111011111111",
55452 => "1111111011111111",
55453 => "1111111011111111",
55454 => "1111111011111111",
55455 => "1111111011111111",
55456 => "1111111011111111",
55457 => "1111111011111111",
55458 => "1111111011111111",
55459 => "1111111011111111",
55460 => "1111111011111111",
55461 => "1111111011111111",
55462 => "1111111011111111",
55463 => "1111111011111111",
55464 => "1111111011111111",
55465 => "1111111100000000",
55466 => "1111111100000000",
55467 => "1111111100000000",
55468 => "1111111100000000",
55469 => "1111111100000000",
55470 => "1111111100000000",
55471 => "1111111100000000",
55472 => "1111111100000000",
55473 => "1111111100000000",
55474 => "1111111100000000",
55475 => "1111111100000000",
55476 => "1111111100000000",
55477 => "1111111100000000",
55478 => "1111111100000000",
55479 => "1111111100000000",
55480 => "1111111100000000",
55481 => "1111111100000001",
55482 => "1111111100000001",
55483 => "1111111100000001",
55484 => "1111111100000001",
55485 => "1111111100000001",
55486 => "1111111100000001",
55487 => "1111111100000001",
55488 => "1111111100000001",
55489 => "1111111100000001",
55490 => "1111111100000001",
55491 => "1111111100000001",
55492 => "1111111100000001",
55493 => "1111111100000001",
55494 => "1111111100000001",
55495 => "1111111100000001",
55496 => "1111111100000001",
55497 => "1111111100000010",
55498 => "1111111100000010",
55499 => "1111111100000010",
55500 => "1111111100000010",
55501 => "1111111100000010",
55502 => "1111111100000010",
55503 => "1111111100000010",
55504 => "1111111100000010",
55505 => "1111111100000010",
55506 => "1111111100000010",
55507 => "1111111100000010",
55508 => "1111111100000010",
55509 => "1111111100000010",
55510 => "1111111100000010",
55511 => "1111111100000010",
55512 => "1111111100000010",
55513 => "1111111100000011",
55514 => "1111111100000011",
55515 => "1111111100000011",
55516 => "1111111100000011",
55517 => "1111111100000011",
55518 => "1111111100000011",
55519 => "1111111100000011",
55520 => "1111111100000011",
55521 => "1111111100000011",
55522 => "1111111100000011",
55523 => "1111111100000011",
55524 => "1111111100000011",
55525 => "1111111100000011",
55526 => "1111111100000011",
55527 => "1111111100000011",
55528 => "1111111100000011",
55529 => "1111111100000100",
55530 => "1111111100000100",
55531 => "1111111100000100",
55532 => "1111111100000100",
55533 => "1111111100000100",
55534 => "1111111100000100",
55535 => "1111111100000100",
55536 => "1111111100000100",
55537 => "1111111100000100",
55538 => "1111111100000100",
55539 => "1111111100000100",
55540 => "1111111100000100",
55541 => "1111111100000100",
55542 => "1111111100000100",
55543 => "1111111100000100",
55544 => "1111111100000100",
55545 => "1111111100000100",
55546 => "1111111100000101",
55547 => "1111111100000101",
55548 => "1111111100000101",
55549 => "1111111100000101",
55550 => "1111111100000101",
55551 => "1111111100000101",
55552 => "1111111100000101",
55553 => "1111111100000101",
55554 => "1111111100000101",
55555 => "1111111100000101",
55556 => "1111111100000101",
55557 => "1111111100000101",
55558 => "1111111100000101",
55559 => "1111111100000101",
55560 => "1111111100000101",
55561 => "1111111100000101",
55562 => "1111111100000110",
55563 => "1111111100000110",
55564 => "1111111100000110",
55565 => "1111111100000110",
55566 => "1111111100000110",
55567 => "1111111100000110",
55568 => "1111111100000110",
55569 => "1111111100000110",
55570 => "1111111100000110",
55571 => "1111111100000110",
55572 => "1111111100000110",
55573 => "1111111100000110",
55574 => "1111111100000110",
55575 => "1111111100000110",
55576 => "1111111100000110",
55577 => "1111111100000110",
55578 => "1111111100000110",
55579 => "1111111100000111",
55580 => "1111111100000111",
55581 => "1111111100000111",
55582 => "1111111100000111",
55583 => "1111111100000111",
55584 => "1111111100000111",
55585 => "1111111100000111",
55586 => "1111111100000111",
55587 => "1111111100000111",
55588 => "1111111100000111",
55589 => "1111111100000111",
55590 => "1111111100000111",
55591 => "1111111100000111",
55592 => "1111111100000111",
55593 => "1111111100000111",
55594 => "1111111100000111",
55595 => "1111111100001000",
55596 => "1111111100001000",
55597 => "1111111100001000",
55598 => "1111111100001000",
55599 => "1111111100001000",
55600 => "1111111100001000",
55601 => "1111111100001000",
55602 => "1111111100001000",
55603 => "1111111100001000",
55604 => "1111111100001000",
55605 => "1111111100001000",
55606 => "1111111100001000",
55607 => "1111111100001000",
55608 => "1111111100001000",
55609 => "1111111100001000",
55610 => "1111111100001000",
55611 => "1111111100001000",
55612 => "1111111100001001",
55613 => "1111111100001001",
55614 => "1111111100001001",
55615 => "1111111100001001",
55616 => "1111111100001001",
55617 => "1111111100001001",
55618 => "1111111100001001",
55619 => "1111111100001001",
55620 => "1111111100001001",
55621 => "1111111100001001",
55622 => "1111111100001001",
55623 => "1111111100001001",
55624 => "1111111100001001",
55625 => "1111111100001001",
55626 => "1111111100001001",
55627 => "1111111100001001",
55628 => "1111111100001001",
55629 => "1111111100001010",
55630 => "1111111100001010",
55631 => "1111111100001010",
55632 => "1111111100001010",
55633 => "1111111100001010",
55634 => "1111111100001010",
55635 => "1111111100001010",
55636 => "1111111100001010",
55637 => "1111111100001010",
55638 => "1111111100001010",
55639 => "1111111100001010",
55640 => "1111111100001010",
55641 => "1111111100001010",
55642 => "1111111100001010",
55643 => "1111111100001010",
55644 => "1111111100001010",
55645 => "1111111100001011",
55646 => "1111111100001011",
55647 => "1111111100001011",
55648 => "1111111100001011",
55649 => "1111111100001011",
55650 => "1111111100001011",
55651 => "1111111100001011",
55652 => "1111111100001011",
55653 => "1111111100001011",
55654 => "1111111100001011",
55655 => "1111111100001011",
55656 => "1111111100001011",
55657 => "1111111100001011",
55658 => "1111111100001011",
55659 => "1111111100001011",
55660 => "1111111100001011",
55661 => "1111111100001011",
55662 => "1111111100001100",
55663 => "1111111100001100",
55664 => "1111111100001100",
55665 => "1111111100001100",
55666 => "1111111100001100",
55667 => "1111111100001100",
55668 => "1111111100001100",
55669 => "1111111100001100",
55670 => "1111111100001100",
55671 => "1111111100001100",
55672 => "1111111100001100",
55673 => "1111111100001100",
55674 => "1111111100001100",
55675 => "1111111100001100",
55676 => "1111111100001100",
55677 => "1111111100001100",
55678 => "1111111100001100",
55679 => "1111111100001101",
55680 => "1111111100001101",
55681 => "1111111100001101",
55682 => "1111111100001101",
55683 => "1111111100001101",
55684 => "1111111100001101",
55685 => "1111111100001101",
55686 => "1111111100001101",
55687 => "1111111100001101",
55688 => "1111111100001101",
55689 => "1111111100001101",
55690 => "1111111100001101",
55691 => "1111111100001101",
55692 => "1111111100001101",
55693 => "1111111100001101",
55694 => "1111111100001101",
55695 => "1111111100001101",
55696 => "1111111100001110",
55697 => "1111111100001110",
55698 => "1111111100001110",
55699 => "1111111100001110",
55700 => "1111111100001110",
55701 => "1111111100001110",
55702 => "1111111100001110",
55703 => "1111111100001110",
55704 => "1111111100001110",
55705 => "1111111100001110",
55706 => "1111111100001110",
55707 => "1111111100001110",
55708 => "1111111100001110",
55709 => "1111111100001110",
55710 => "1111111100001110",
55711 => "1111111100001110",
55712 => "1111111100001110",
55713 => "1111111100001111",
55714 => "1111111100001111",
55715 => "1111111100001111",
55716 => "1111111100001111",
55717 => "1111111100001111",
55718 => "1111111100001111",
55719 => "1111111100001111",
55720 => "1111111100001111",
55721 => "1111111100001111",
55722 => "1111111100001111",
55723 => "1111111100001111",
55724 => "1111111100001111",
55725 => "1111111100001111",
55726 => "1111111100001111",
55727 => "1111111100001111",
55728 => "1111111100001111",
55729 => "1111111100001111",
55730 => "1111111100010000",
55731 => "1111111100010000",
55732 => "1111111100010000",
55733 => "1111111100010000",
55734 => "1111111100010000",
55735 => "1111111100010000",
55736 => "1111111100010000",
55737 => "1111111100010000",
55738 => "1111111100010000",
55739 => "1111111100010000",
55740 => "1111111100010000",
55741 => "1111111100010000",
55742 => "1111111100010000",
55743 => "1111111100010000",
55744 => "1111111100010000",
55745 => "1111111100010000",
55746 => "1111111100010000",
55747 => "1111111100010001",
55748 => "1111111100010001",
55749 => "1111111100010001",
55750 => "1111111100010001",
55751 => "1111111100010001",
55752 => "1111111100010001",
55753 => "1111111100010001",
55754 => "1111111100010001",
55755 => "1111111100010001",
55756 => "1111111100010001",
55757 => "1111111100010001",
55758 => "1111111100010001",
55759 => "1111111100010001",
55760 => "1111111100010001",
55761 => "1111111100010001",
55762 => "1111111100010001",
55763 => "1111111100010001",
55764 => "1111111100010010",
55765 => "1111111100010010",
55766 => "1111111100010010",
55767 => "1111111100010010",
55768 => "1111111100010010",
55769 => "1111111100010010",
55770 => "1111111100010010",
55771 => "1111111100010010",
55772 => "1111111100010010",
55773 => "1111111100010010",
55774 => "1111111100010010",
55775 => "1111111100010010",
55776 => "1111111100010010",
55777 => "1111111100010010",
55778 => "1111111100010010",
55779 => "1111111100010010",
55780 => "1111111100010010",
55781 => "1111111100010010",
55782 => "1111111100010011",
55783 => "1111111100010011",
55784 => "1111111100010011",
55785 => "1111111100010011",
55786 => "1111111100010011",
55787 => "1111111100010011",
55788 => "1111111100010011",
55789 => "1111111100010011",
55790 => "1111111100010011",
55791 => "1111111100010011",
55792 => "1111111100010011",
55793 => "1111111100010011",
55794 => "1111111100010011",
55795 => "1111111100010011",
55796 => "1111111100010011",
55797 => "1111111100010011",
55798 => "1111111100010011",
55799 => "1111111100010100",
55800 => "1111111100010100",
55801 => "1111111100010100",
55802 => "1111111100010100",
55803 => "1111111100010100",
55804 => "1111111100010100",
55805 => "1111111100010100",
55806 => "1111111100010100",
55807 => "1111111100010100",
55808 => "1111111100010100",
55809 => "1111111100010100",
55810 => "1111111100010100",
55811 => "1111111100010100",
55812 => "1111111100010100",
55813 => "1111111100010100",
55814 => "1111111100010100",
55815 => "1111111100010100",
55816 => "1111111100010100",
55817 => "1111111100010101",
55818 => "1111111100010101",
55819 => "1111111100010101",
55820 => "1111111100010101",
55821 => "1111111100010101",
55822 => "1111111100010101",
55823 => "1111111100010101",
55824 => "1111111100010101",
55825 => "1111111100010101",
55826 => "1111111100010101",
55827 => "1111111100010101",
55828 => "1111111100010101",
55829 => "1111111100010101",
55830 => "1111111100010101",
55831 => "1111111100010101",
55832 => "1111111100010101",
55833 => "1111111100010101",
55834 => "1111111100010110",
55835 => "1111111100010110",
55836 => "1111111100010110",
55837 => "1111111100010110",
55838 => "1111111100010110",
55839 => "1111111100010110",
55840 => "1111111100010110",
55841 => "1111111100010110",
55842 => "1111111100010110",
55843 => "1111111100010110",
55844 => "1111111100010110",
55845 => "1111111100010110",
55846 => "1111111100010110",
55847 => "1111111100010110",
55848 => "1111111100010110",
55849 => "1111111100010110",
55850 => "1111111100010110",
55851 => "1111111100010110",
55852 => "1111111100010111",
55853 => "1111111100010111",
55854 => "1111111100010111",
55855 => "1111111100010111",
55856 => "1111111100010111",
55857 => "1111111100010111",
55858 => "1111111100010111",
55859 => "1111111100010111",
55860 => "1111111100010111",
55861 => "1111111100010111",
55862 => "1111111100010111",
55863 => "1111111100010111",
55864 => "1111111100010111",
55865 => "1111111100010111",
55866 => "1111111100010111",
55867 => "1111111100010111",
55868 => "1111111100010111",
55869 => "1111111100011000",
55870 => "1111111100011000",
55871 => "1111111100011000",
55872 => "1111111100011000",
55873 => "1111111100011000",
55874 => "1111111100011000",
55875 => "1111111100011000",
55876 => "1111111100011000",
55877 => "1111111100011000",
55878 => "1111111100011000",
55879 => "1111111100011000",
55880 => "1111111100011000",
55881 => "1111111100011000",
55882 => "1111111100011000",
55883 => "1111111100011000",
55884 => "1111111100011000",
55885 => "1111111100011000",
55886 => "1111111100011000",
55887 => "1111111100011001",
55888 => "1111111100011001",
55889 => "1111111100011001",
55890 => "1111111100011001",
55891 => "1111111100011001",
55892 => "1111111100011001",
55893 => "1111111100011001",
55894 => "1111111100011001",
55895 => "1111111100011001",
55896 => "1111111100011001",
55897 => "1111111100011001",
55898 => "1111111100011001",
55899 => "1111111100011001",
55900 => "1111111100011001",
55901 => "1111111100011001",
55902 => "1111111100011001",
55903 => "1111111100011001",
55904 => "1111111100011001",
55905 => "1111111100011010",
55906 => "1111111100011010",
55907 => "1111111100011010",
55908 => "1111111100011010",
55909 => "1111111100011010",
55910 => "1111111100011010",
55911 => "1111111100011010",
55912 => "1111111100011010",
55913 => "1111111100011010",
55914 => "1111111100011010",
55915 => "1111111100011010",
55916 => "1111111100011010",
55917 => "1111111100011010",
55918 => "1111111100011010",
55919 => "1111111100011010",
55920 => "1111111100011010",
55921 => "1111111100011010",
55922 => "1111111100011010",
55923 => "1111111100011011",
55924 => "1111111100011011",
55925 => "1111111100011011",
55926 => "1111111100011011",
55927 => "1111111100011011",
55928 => "1111111100011011",
55929 => "1111111100011011",
55930 => "1111111100011011",
55931 => "1111111100011011",
55932 => "1111111100011011",
55933 => "1111111100011011",
55934 => "1111111100011011",
55935 => "1111111100011011",
55936 => "1111111100011011",
55937 => "1111111100011011",
55938 => "1111111100011011",
55939 => "1111111100011011",
55940 => "1111111100011011",
55941 => "1111111100011100",
55942 => "1111111100011100",
55943 => "1111111100011100",
55944 => "1111111100011100",
55945 => "1111111100011100",
55946 => "1111111100011100",
55947 => "1111111100011100",
55948 => "1111111100011100",
55949 => "1111111100011100",
55950 => "1111111100011100",
55951 => "1111111100011100",
55952 => "1111111100011100",
55953 => "1111111100011100",
55954 => "1111111100011100",
55955 => "1111111100011100",
55956 => "1111111100011100",
55957 => "1111111100011100",
55958 => "1111111100011100",
55959 => "1111111100011101",
55960 => "1111111100011101",
55961 => "1111111100011101",
55962 => "1111111100011101",
55963 => "1111111100011101",
55964 => "1111111100011101",
55965 => "1111111100011101",
55966 => "1111111100011101",
55967 => "1111111100011101",
55968 => "1111111100011101",
55969 => "1111111100011101",
55970 => "1111111100011101",
55971 => "1111111100011101",
55972 => "1111111100011101",
55973 => "1111111100011101",
55974 => "1111111100011101",
55975 => "1111111100011101",
55976 => "1111111100011101",
55977 => "1111111100011110",
55978 => "1111111100011110",
55979 => "1111111100011110",
55980 => "1111111100011110",
55981 => "1111111100011110",
55982 => "1111111100011110",
55983 => "1111111100011110",
55984 => "1111111100011110",
55985 => "1111111100011110",
55986 => "1111111100011110",
55987 => "1111111100011110",
55988 => "1111111100011110",
55989 => "1111111100011110",
55990 => "1111111100011110",
55991 => "1111111100011110",
55992 => "1111111100011110",
55993 => "1111111100011110",
55994 => "1111111100011110",
55995 => "1111111100011111",
55996 => "1111111100011111",
55997 => "1111111100011111",
55998 => "1111111100011111",
55999 => "1111111100011111",
56000 => "1111111100011111",
56001 => "1111111100011111",
56002 => "1111111100011111",
56003 => "1111111100011111",
56004 => "1111111100011111",
56005 => "1111111100011111",
56006 => "1111111100011111",
56007 => "1111111100011111",
56008 => "1111111100011111",
56009 => "1111111100011111",
56010 => "1111111100011111",
56011 => "1111111100011111",
56012 => "1111111100011111",
56013 => "1111111100011111",
56014 => "1111111100100000",
56015 => "1111111100100000",
56016 => "1111111100100000",
56017 => "1111111100100000",
56018 => "1111111100100000",
56019 => "1111111100100000",
56020 => "1111111100100000",
56021 => "1111111100100000",
56022 => "1111111100100000",
56023 => "1111111100100000",
56024 => "1111111100100000",
56025 => "1111111100100000",
56026 => "1111111100100000",
56027 => "1111111100100000",
56028 => "1111111100100000",
56029 => "1111111100100000",
56030 => "1111111100100000",
56031 => "1111111100100000",
56032 => "1111111100100001",
56033 => "1111111100100001",
56034 => "1111111100100001",
56035 => "1111111100100001",
56036 => "1111111100100001",
56037 => "1111111100100001",
56038 => "1111111100100001",
56039 => "1111111100100001",
56040 => "1111111100100001",
56041 => "1111111100100001",
56042 => "1111111100100001",
56043 => "1111111100100001",
56044 => "1111111100100001",
56045 => "1111111100100001",
56046 => "1111111100100001",
56047 => "1111111100100001",
56048 => "1111111100100001",
56049 => "1111111100100001",
56050 => "1111111100100010",
56051 => "1111111100100010",
56052 => "1111111100100010",
56053 => "1111111100100010",
56054 => "1111111100100010",
56055 => "1111111100100010",
56056 => "1111111100100010",
56057 => "1111111100100010",
56058 => "1111111100100010",
56059 => "1111111100100010",
56060 => "1111111100100010",
56061 => "1111111100100010",
56062 => "1111111100100010",
56063 => "1111111100100010",
56064 => "1111111100100010",
56065 => "1111111100100010",
56066 => "1111111100100010",
56067 => "1111111100100010",
56068 => "1111111100100010",
56069 => "1111111100100011",
56070 => "1111111100100011",
56071 => "1111111100100011",
56072 => "1111111100100011",
56073 => "1111111100100011",
56074 => "1111111100100011",
56075 => "1111111100100011",
56076 => "1111111100100011",
56077 => "1111111100100011",
56078 => "1111111100100011",
56079 => "1111111100100011",
56080 => "1111111100100011",
56081 => "1111111100100011",
56082 => "1111111100100011",
56083 => "1111111100100011",
56084 => "1111111100100011",
56085 => "1111111100100011",
56086 => "1111111100100011",
56087 => "1111111100100011",
56088 => "1111111100100100",
56089 => "1111111100100100",
56090 => "1111111100100100",
56091 => "1111111100100100",
56092 => "1111111100100100",
56093 => "1111111100100100",
56094 => "1111111100100100",
56095 => "1111111100100100",
56096 => "1111111100100100",
56097 => "1111111100100100",
56098 => "1111111100100100",
56099 => "1111111100100100",
56100 => "1111111100100100",
56101 => "1111111100100100",
56102 => "1111111100100100",
56103 => "1111111100100100",
56104 => "1111111100100100",
56105 => "1111111100100100",
56106 => "1111111100100101",
56107 => "1111111100100101",
56108 => "1111111100100101",
56109 => "1111111100100101",
56110 => "1111111100100101",
56111 => "1111111100100101",
56112 => "1111111100100101",
56113 => "1111111100100101",
56114 => "1111111100100101",
56115 => "1111111100100101",
56116 => "1111111100100101",
56117 => "1111111100100101",
56118 => "1111111100100101",
56119 => "1111111100100101",
56120 => "1111111100100101",
56121 => "1111111100100101",
56122 => "1111111100100101",
56123 => "1111111100100101",
56124 => "1111111100100101",
56125 => "1111111100100110",
56126 => "1111111100100110",
56127 => "1111111100100110",
56128 => "1111111100100110",
56129 => "1111111100100110",
56130 => "1111111100100110",
56131 => "1111111100100110",
56132 => "1111111100100110",
56133 => "1111111100100110",
56134 => "1111111100100110",
56135 => "1111111100100110",
56136 => "1111111100100110",
56137 => "1111111100100110",
56138 => "1111111100100110",
56139 => "1111111100100110",
56140 => "1111111100100110",
56141 => "1111111100100110",
56142 => "1111111100100110",
56143 => "1111111100100110",
56144 => "1111111100100111",
56145 => "1111111100100111",
56146 => "1111111100100111",
56147 => "1111111100100111",
56148 => "1111111100100111",
56149 => "1111111100100111",
56150 => "1111111100100111",
56151 => "1111111100100111",
56152 => "1111111100100111",
56153 => "1111111100100111",
56154 => "1111111100100111",
56155 => "1111111100100111",
56156 => "1111111100100111",
56157 => "1111111100100111",
56158 => "1111111100100111",
56159 => "1111111100100111",
56160 => "1111111100100111",
56161 => "1111111100100111",
56162 => "1111111100100111",
56163 => "1111111100101000",
56164 => "1111111100101000",
56165 => "1111111100101000",
56166 => "1111111100101000",
56167 => "1111111100101000",
56168 => "1111111100101000",
56169 => "1111111100101000",
56170 => "1111111100101000",
56171 => "1111111100101000",
56172 => "1111111100101000",
56173 => "1111111100101000",
56174 => "1111111100101000",
56175 => "1111111100101000",
56176 => "1111111100101000",
56177 => "1111111100101000",
56178 => "1111111100101000",
56179 => "1111111100101000",
56180 => "1111111100101000",
56181 => "1111111100101000",
56182 => "1111111100101001",
56183 => "1111111100101001",
56184 => "1111111100101001",
56185 => "1111111100101001",
56186 => "1111111100101001",
56187 => "1111111100101001",
56188 => "1111111100101001",
56189 => "1111111100101001",
56190 => "1111111100101001",
56191 => "1111111100101001",
56192 => "1111111100101001",
56193 => "1111111100101001",
56194 => "1111111100101001",
56195 => "1111111100101001",
56196 => "1111111100101001",
56197 => "1111111100101001",
56198 => "1111111100101001",
56199 => "1111111100101001",
56200 => "1111111100101001",
56201 => "1111111100101010",
56202 => "1111111100101010",
56203 => "1111111100101010",
56204 => "1111111100101010",
56205 => "1111111100101010",
56206 => "1111111100101010",
56207 => "1111111100101010",
56208 => "1111111100101010",
56209 => "1111111100101010",
56210 => "1111111100101010",
56211 => "1111111100101010",
56212 => "1111111100101010",
56213 => "1111111100101010",
56214 => "1111111100101010",
56215 => "1111111100101010",
56216 => "1111111100101010",
56217 => "1111111100101010",
56218 => "1111111100101010",
56219 => "1111111100101010",
56220 => "1111111100101010",
56221 => "1111111100101011",
56222 => "1111111100101011",
56223 => "1111111100101011",
56224 => "1111111100101011",
56225 => "1111111100101011",
56226 => "1111111100101011",
56227 => "1111111100101011",
56228 => "1111111100101011",
56229 => "1111111100101011",
56230 => "1111111100101011",
56231 => "1111111100101011",
56232 => "1111111100101011",
56233 => "1111111100101011",
56234 => "1111111100101011",
56235 => "1111111100101011",
56236 => "1111111100101011",
56237 => "1111111100101011",
56238 => "1111111100101011",
56239 => "1111111100101011",
56240 => "1111111100101100",
56241 => "1111111100101100",
56242 => "1111111100101100",
56243 => "1111111100101100",
56244 => "1111111100101100",
56245 => "1111111100101100",
56246 => "1111111100101100",
56247 => "1111111100101100",
56248 => "1111111100101100",
56249 => "1111111100101100",
56250 => "1111111100101100",
56251 => "1111111100101100",
56252 => "1111111100101100",
56253 => "1111111100101100",
56254 => "1111111100101100",
56255 => "1111111100101100",
56256 => "1111111100101100",
56257 => "1111111100101100",
56258 => "1111111100101100",
56259 => "1111111100101101",
56260 => "1111111100101101",
56261 => "1111111100101101",
56262 => "1111111100101101",
56263 => "1111111100101101",
56264 => "1111111100101101",
56265 => "1111111100101101",
56266 => "1111111100101101",
56267 => "1111111100101101",
56268 => "1111111100101101",
56269 => "1111111100101101",
56270 => "1111111100101101",
56271 => "1111111100101101",
56272 => "1111111100101101",
56273 => "1111111100101101",
56274 => "1111111100101101",
56275 => "1111111100101101",
56276 => "1111111100101101",
56277 => "1111111100101101",
56278 => "1111111100101101",
56279 => "1111111100101110",
56280 => "1111111100101110",
56281 => "1111111100101110",
56282 => "1111111100101110",
56283 => "1111111100101110",
56284 => "1111111100101110",
56285 => "1111111100101110",
56286 => "1111111100101110",
56287 => "1111111100101110",
56288 => "1111111100101110",
56289 => "1111111100101110",
56290 => "1111111100101110",
56291 => "1111111100101110",
56292 => "1111111100101110",
56293 => "1111111100101110",
56294 => "1111111100101110",
56295 => "1111111100101110",
56296 => "1111111100101110",
56297 => "1111111100101110",
56298 => "1111111100101111",
56299 => "1111111100101111",
56300 => "1111111100101111",
56301 => "1111111100101111",
56302 => "1111111100101111",
56303 => "1111111100101111",
56304 => "1111111100101111",
56305 => "1111111100101111",
56306 => "1111111100101111",
56307 => "1111111100101111",
56308 => "1111111100101111",
56309 => "1111111100101111",
56310 => "1111111100101111",
56311 => "1111111100101111",
56312 => "1111111100101111",
56313 => "1111111100101111",
56314 => "1111111100101111",
56315 => "1111111100101111",
56316 => "1111111100101111",
56317 => "1111111100101111",
56318 => "1111111100110000",
56319 => "1111111100110000",
56320 => "1111111100110000",
56321 => "1111111100110000",
56322 => "1111111100110000",
56323 => "1111111100110000",
56324 => "1111111100110000",
56325 => "1111111100110000",
56326 => "1111111100110000",
56327 => "1111111100110000",
56328 => "1111111100110000",
56329 => "1111111100110000",
56330 => "1111111100110000",
56331 => "1111111100110000",
56332 => "1111111100110000",
56333 => "1111111100110000",
56334 => "1111111100110000",
56335 => "1111111100110000",
56336 => "1111111100110000",
56337 => "1111111100110000",
56338 => "1111111100110001",
56339 => "1111111100110001",
56340 => "1111111100110001",
56341 => "1111111100110001",
56342 => "1111111100110001",
56343 => "1111111100110001",
56344 => "1111111100110001",
56345 => "1111111100110001",
56346 => "1111111100110001",
56347 => "1111111100110001",
56348 => "1111111100110001",
56349 => "1111111100110001",
56350 => "1111111100110001",
56351 => "1111111100110001",
56352 => "1111111100110001",
56353 => "1111111100110001",
56354 => "1111111100110001",
56355 => "1111111100110001",
56356 => "1111111100110001",
56357 => "1111111100110001",
56358 => "1111111100110010",
56359 => "1111111100110010",
56360 => "1111111100110010",
56361 => "1111111100110010",
56362 => "1111111100110010",
56363 => "1111111100110010",
56364 => "1111111100110010",
56365 => "1111111100110010",
56366 => "1111111100110010",
56367 => "1111111100110010",
56368 => "1111111100110010",
56369 => "1111111100110010",
56370 => "1111111100110010",
56371 => "1111111100110010",
56372 => "1111111100110010",
56373 => "1111111100110010",
56374 => "1111111100110010",
56375 => "1111111100110010",
56376 => "1111111100110010",
56377 => "1111111100110010",
56378 => "1111111100110011",
56379 => "1111111100110011",
56380 => "1111111100110011",
56381 => "1111111100110011",
56382 => "1111111100110011",
56383 => "1111111100110011",
56384 => "1111111100110011",
56385 => "1111111100110011",
56386 => "1111111100110011",
56387 => "1111111100110011",
56388 => "1111111100110011",
56389 => "1111111100110011",
56390 => "1111111100110011",
56391 => "1111111100110011",
56392 => "1111111100110011",
56393 => "1111111100110011",
56394 => "1111111100110011",
56395 => "1111111100110011",
56396 => "1111111100110011",
56397 => "1111111100110011",
56398 => "1111111100110100",
56399 => "1111111100110100",
56400 => "1111111100110100",
56401 => "1111111100110100",
56402 => "1111111100110100",
56403 => "1111111100110100",
56404 => "1111111100110100",
56405 => "1111111100110100",
56406 => "1111111100110100",
56407 => "1111111100110100",
56408 => "1111111100110100",
56409 => "1111111100110100",
56410 => "1111111100110100",
56411 => "1111111100110100",
56412 => "1111111100110100",
56413 => "1111111100110100",
56414 => "1111111100110100",
56415 => "1111111100110100",
56416 => "1111111100110100",
56417 => "1111111100110100",
56418 => "1111111100110101",
56419 => "1111111100110101",
56420 => "1111111100110101",
56421 => "1111111100110101",
56422 => "1111111100110101",
56423 => "1111111100110101",
56424 => "1111111100110101",
56425 => "1111111100110101",
56426 => "1111111100110101",
56427 => "1111111100110101",
56428 => "1111111100110101",
56429 => "1111111100110101",
56430 => "1111111100110101",
56431 => "1111111100110101",
56432 => "1111111100110101",
56433 => "1111111100110101",
56434 => "1111111100110101",
56435 => "1111111100110101",
56436 => "1111111100110101",
56437 => "1111111100110101",
56438 => "1111111100110110",
56439 => "1111111100110110",
56440 => "1111111100110110",
56441 => "1111111100110110",
56442 => "1111111100110110",
56443 => "1111111100110110",
56444 => "1111111100110110",
56445 => "1111111100110110",
56446 => "1111111100110110",
56447 => "1111111100110110",
56448 => "1111111100110110",
56449 => "1111111100110110",
56450 => "1111111100110110",
56451 => "1111111100110110",
56452 => "1111111100110110",
56453 => "1111111100110110",
56454 => "1111111100110110",
56455 => "1111111100110110",
56456 => "1111111100110110",
56457 => "1111111100110110",
56458 => "1111111100110110",
56459 => "1111111100110111",
56460 => "1111111100110111",
56461 => "1111111100110111",
56462 => "1111111100110111",
56463 => "1111111100110111",
56464 => "1111111100110111",
56465 => "1111111100110111",
56466 => "1111111100110111",
56467 => "1111111100110111",
56468 => "1111111100110111",
56469 => "1111111100110111",
56470 => "1111111100110111",
56471 => "1111111100110111",
56472 => "1111111100110111",
56473 => "1111111100110111",
56474 => "1111111100110111",
56475 => "1111111100110111",
56476 => "1111111100110111",
56477 => "1111111100110111",
56478 => "1111111100110111",
56479 => "1111111100111000",
56480 => "1111111100111000",
56481 => "1111111100111000",
56482 => "1111111100111000",
56483 => "1111111100111000",
56484 => "1111111100111000",
56485 => "1111111100111000",
56486 => "1111111100111000",
56487 => "1111111100111000",
56488 => "1111111100111000",
56489 => "1111111100111000",
56490 => "1111111100111000",
56491 => "1111111100111000",
56492 => "1111111100111000",
56493 => "1111111100111000",
56494 => "1111111100111000",
56495 => "1111111100111000",
56496 => "1111111100111000",
56497 => "1111111100111000",
56498 => "1111111100111000",
56499 => "1111111100111000",
56500 => "1111111100111001",
56501 => "1111111100111001",
56502 => "1111111100111001",
56503 => "1111111100111001",
56504 => "1111111100111001",
56505 => "1111111100111001",
56506 => "1111111100111001",
56507 => "1111111100111001",
56508 => "1111111100111001",
56509 => "1111111100111001",
56510 => "1111111100111001",
56511 => "1111111100111001",
56512 => "1111111100111001",
56513 => "1111111100111001",
56514 => "1111111100111001",
56515 => "1111111100111001",
56516 => "1111111100111001",
56517 => "1111111100111001",
56518 => "1111111100111001",
56519 => "1111111100111001",
56520 => "1111111100111001",
56521 => "1111111100111010",
56522 => "1111111100111010",
56523 => "1111111100111010",
56524 => "1111111100111010",
56525 => "1111111100111010",
56526 => "1111111100111010",
56527 => "1111111100111010",
56528 => "1111111100111010",
56529 => "1111111100111010",
56530 => "1111111100111010",
56531 => "1111111100111010",
56532 => "1111111100111010",
56533 => "1111111100111010",
56534 => "1111111100111010",
56535 => "1111111100111010",
56536 => "1111111100111010",
56537 => "1111111100111010",
56538 => "1111111100111010",
56539 => "1111111100111010",
56540 => "1111111100111010",
56541 => "1111111100111011",
56542 => "1111111100111011",
56543 => "1111111100111011",
56544 => "1111111100111011",
56545 => "1111111100111011",
56546 => "1111111100111011",
56547 => "1111111100111011",
56548 => "1111111100111011",
56549 => "1111111100111011",
56550 => "1111111100111011",
56551 => "1111111100111011",
56552 => "1111111100111011",
56553 => "1111111100111011",
56554 => "1111111100111011",
56555 => "1111111100111011",
56556 => "1111111100111011",
56557 => "1111111100111011",
56558 => "1111111100111011",
56559 => "1111111100111011",
56560 => "1111111100111011",
56561 => "1111111100111011",
56562 => "1111111100111100",
56563 => "1111111100111100",
56564 => "1111111100111100",
56565 => "1111111100111100",
56566 => "1111111100111100",
56567 => "1111111100111100",
56568 => "1111111100111100",
56569 => "1111111100111100",
56570 => "1111111100111100",
56571 => "1111111100111100",
56572 => "1111111100111100",
56573 => "1111111100111100",
56574 => "1111111100111100",
56575 => "1111111100111100",
56576 => "1111111100111100",
56577 => "1111111100111100",
56578 => "1111111100111100",
56579 => "1111111100111100",
56580 => "1111111100111100",
56581 => "1111111100111100",
56582 => "1111111100111100",
56583 => "1111111100111101",
56584 => "1111111100111101",
56585 => "1111111100111101",
56586 => "1111111100111101",
56587 => "1111111100111101",
56588 => "1111111100111101",
56589 => "1111111100111101",
56590 => "1111111100111101",
56591 => "1111111100111101",
56592 => "1111111100111101",
56593 => "1111111100111101",
56594 => "1111111100111101",
56595 => "1111111100111101",
56596 => "1111111100111101",
56597 => "1111111100111101",
56598 => "1111111100111101",
56599 => "1111111100111101",
56600 => "1111111100111101",
56601 => "1111111100111101",
56602 => "1111111100111101",
56603 => "1111111100111101",
56604 => "1111111100111110",
56605 => "1111111100111110",
56606 => "1111111100111110",
56607 => "1111111100111110",
56608 => "1111111100111110",
56609 => "1111111100111110",
56610 => "1111111100111110",
56611 => "1111111100111110",
56612 => "1111111100111110",
56613 => "1111111100111110",
56614 => "1111111100111110",
56615 => "1111111100111110",
56616 => "1111111100111110",
56617 => "1111111100111110",
56618 => "1111111100111110",
56619 => "1111111100111110",
56620 => "1111111100111110",
56621 => "1111111100111110",
56622 => "1111111100111110",
56623 => "1111111100111110",
56624 => "1111111100111110",
56625 => "1111111100111110",
56626 => "1111111100111111",
56627 => "1111111100111111",
56628 => "1111111100111111",
56629 => "1111111100111111",
56630 => "1111111100111111",
56631 => "1111111100111111",
56632 => "1111111100111111",
56633 => "1111111100111111",
56634 => "1111111100111111",
56635 => "1111111100111111",
56636 => "1111111100111111",
56637 => "1111111100111111",
56638 => "1111111100111111",
56639 => "1111111100111111",
56640 => "1111111100111111",
56641 => "1111111100111111",
56642 => "1111111100111111",
56643 => "1111111100111111",
56644 => "1111111100111111",
56645 => "1111111100111111",
56646 => "1111111100111111",
56647 => "1111111101000000",
56648 => "1111111101000000",
56649 => "1111111101000000",
56650 => "1111111101000000",
56651 => "1111111101000000",
56652 => "1111111101000000",
56653 => "1111111101000000",
56654 => "1111111101000000",
56655 => "1111111101000000",
56656 => "1111111101000000",
56657 => "1111111101000000",
56658 => "1111111101000000",
56659 => "1111111101000000",
56660 => "1111111101000000",
56661 => "1111111101000000",
56662 => "1111111101000000",
56663 => "1111111101000000",
56664 => "1111111101000000",
56665 => "1111111101000000",
56666 => "1111111101000000",
56667 => "1111111101000000",
56668 => "1111111101000001",
56669 => "1111111101000001",
56670 => "1111111101000001",
56671 => "1111111101000001",
56672 => "1111111101000001",
56673 => "1111111101000001",
56674 => "1111111101000001",
56675 => "1111111101000001",
56676 => "1111111101000001",
56677 => "1111111101000001",
56678 => "1111111101000001",
56679 => "1111111101000001",
56680 => "1111111101000001",
56681 => "1111111101000001",
56682 => "1111111101000001",
56683 => "1111111101000001",
56684 => "1111111101000001",
56685 => "1111111101000001",
56686 => "1111111101000001",
56687 => "1111111101000001",
56688 => "1111111101000001",
56689 => "1111111101000001",
56690 => "1111111101000010",
56691 => "1111111101000010",
56692 => "1111111101000010",
56693 => "1111111101000010",
56694 => "1111111101000010",
56695 => "1111111101000010",
56696 => "1111111101000010",
56697 => "1111111101000010",
56698 => "1111111101000010",
56699 => "1111111101000010",
56700 => "1111111101000010",
56701 => "1111111101000010",
56702 => "1111111101000010",
56703 => "1111111101000010",
56704 => "1111111101000010",
56705 => "1111111101000010",
56706 => "1111111101000010",
56707 => "1111111101000010",
56708 => "1111111101000010",
56709 => "1111111101000010",
56710 => "1111111101000010",
56711 => "1111111101000010",
56712 => "1111111101000011",
56713 => "1111111101000011",
56714 => "1111111101000011",
56715 => "1111111101000011",
56716 => "1111111101000011",
56717 => "1111111101000011",
56718 => "1111111101000011",
56719 => "1111111101000011",
56720 => "1111111101000011",
56721 => "1111111101000011",
56722 => "1111111101000011",
56723 => "1111111101000011",
56724 => "1111111101000011",
56725 => "1111111101000011",
56726 => "1111111101000011",
56727 => "1111111101000011",
56728 => "1111111101000011",
56729 => "1111111101000011",
56730 => "1111111101000011",
56731 => "1111111101000011",
56732 => "1111111101000011",
56733 => "1111111101000100",
56734 => "1111111101000100",
56735 => "1111111101000100",
56736 => "1111111101000100",
56737 => "1111111101000100",
56738 => "1111111101000100",
56739 => "1111111101000100",
56740 => "1111111101000100",
56741 => "1111111101000100",
56742 => "1111111101000100",
56743 => "1111111101000100",
56744 => "1111111101000100",
56745 => "1111111101000100",
56746 => "1111111101000100",
56747 => "1111111101000100",
56748 => "1111111101000100",
56749 => "1111111101000100",
56750 => "1111111101000100",
56751 => "1111111101000100",
56752 => "1111111101000100",
56753 => "1111111101000100",
56754 => "1111111101000100",
56755 => "1111111101000101",
56756 => "1111111101000101",
56757 => "1111111101000101",
56758 => "1111111101000101",
56759 => "1111111101000101",
56760 => "1111111101000101",
56761 => "1111111101000101",
56762 => "1111111101000101",
56763 => "1111111101000101",
56764 => "1111111101000101",
56765 => "1111111101000101",
56766 => "1111111101000101",
56767 => "1111111101000101",
56768 => "1111111101000101",
56769 => "1111111101000101",
56770 => "1111111101000101",
56771 => "1111111101000101",
56772 => "1111111101000101",
56773 => "1111111101000101",
56774 => "1111111101000101",
56775 => "1111111101000101",
56776 => "1111111101000101",
56777 => "1111111101000110",
56778 => "1111111101000110",
56779 => "1111111101000110",
56780 => "1111111101000110",
56781 => "1111111101000110",
56782 => "1111111101000110",
56783 => "1111111101000110",
56784 => "1111111101000110",
56785 => "1111111101000110",
56786 => "1111111101000110",
56787 => "1111111101000110",
56788 => "1111111101000110",
56789 => "1111111101000110",
56790 => "1111111101000110",
56791 => "1111111101000110",
56792 => "1111111101000110",
56793 => "1111111101000110",
56794 => "1111111101000110",
56795 => "1111111101000110",
56796 => "1111111101000110",
56797 => "1111111101000110",
56798 => "1111111101000110",
56799 => "1111111101000110",
56800 => "1111111101000111",
56801 => "1111111101000111",
56802 => "1111111101000111",
56803 => "1111111101000111",
56804 => "1111111101000111",
56805 => "1111111101000111",
56806 => "1111111101000111",
56807 => "1111111101000111",
56808 => "1111111101000111",
56809 => "1111111101000111",
56810 => "1111111101000111",
56811 => "1111111101000111",
56812 => "1111111101000111",
56813 => "1111111101000111",
56814 => "1111111101000111",
56815 => "1111111101000111",
56816 => "1111111101000111",
56817 => "1111111101000111",
56818 => "1111111101000111",
56819 => "1111111101000111",
56820 => "1111111101000111",
56821 => "1111111101000111",
56822 => "1111111101001000",
56823 => "1111111101001000",
56824 => "1111111101001000",
56825 => "1111111101001000",
56826 => "1111111101001000",
56827 => "1111111101001000",
56828 => "1111111101001000",
56829 => "1111111101001000",
56830 => "1111111101001000",
56831 => "1111111101001000",
56832 => "1111111101001000",
56833 => "1111111101001000",
56834 => "1111111101001000",
56835 => "1111111101001000",
56836 => "1111111101001000",
56837 => "1111111101001000",
56838 => "1111111101001000",
56839 => "1111111101001000",
56840 => "1111111101001000",
56841 => "1111111101001000",
56842 => "1111111101001000",
56843 => "1111111101001000",
56844 => "1111111101001001",
56845 => "1111111101001001",
56846 => "1111111101001001",
56847 => "1111111101001001",
56848 => "1111111101001001",
56849 => "1111111101001001",
56850 => "1111111101001001",
56851 => "1111111101001001",
56852 => "1111111101001001",
56853 => "1111111101001001",
56854 => "1111111101001001",
56855 => "1111111101001001",
56856 => "1111111101001001",
56857 => "1111111101001001",
56858 => "1111111101001001",
56859 => "1111111101001001",
56860 => "1111111101001001",
56861 => "1111111101001001",
56862 => "1111111101001001",
56863 => "1111111101001001",
56864 => "1111111101001001",
56865 => "1111111101001001",
56866 => "1111111101001001",
56867 => "1111111101001010",
56868 => "1111111101001010",
56869 => "1111111101001010",
56870 => "1111111101001010",
56871 => "1111111101001010",
56872 => "1111111101001010",
56873 => "1111111101001010",
56874 => "1111111101001010",
56875 => "1111111101001010",
56876 => "1111111101001010",
56877 => "1111111101001010",
56878 => "1111111101001010",
56879 => "1111111101001010",
56880 => "1111111101001010",
56881 => "1111111101001010",
56882 => "1111111101001010",
56883 => "1111111101001010",
56884 => "1111111101001010",
56885 => "1111111101001010",
56886 => "1111111101001010",
56887 => "1111111101001010",
56888 => "1111111101001010",
56889 => "1111111101001011",
56890 => "1111111101001011",
56891 => "1111111101001011",
56892 => "1111111101001011",
56893 => "1111111101001011",
56894 => "1111111101001011",
56895 => "1111111101001011",
56896 => "1111111101001011",
56897 => "1111111101001011",
56898 => "1111111101001011",
56899 => "1111111101001011",
56900 => "1111111101001011",
56901 => "1111111101001011",
56902 => "1111111101001011",
56903 => "1111111101001011",
56904 => "1111111101001011",
56905 => "1111111101001011",
56906 => "1111111101001011",
56907 => "1111111101001011",
56908 => "1111111101001011",
56909 => "1111111101001011",
56910 => "1111111101001011",
56911 => "1111111101001011",
56912 => "1111111101001100",
56913 => "1111111101001100",
56914 => "1111111101001100",
56915 => "1111111101001100",
56916 => "1111111101001100",
56917 => "1111111101001100",
56918 => "1111111101001100",
56919 => "1111111101001100",
56920 => "1111111101001100",
56921 => "1111111101001100",
56922 => "1111111101001100",
56923 => "1111111101001100",
56924 => "1111111101001100",
56925 => "1111111101001100",
56926 => "1111111101001100",
56927 => "1111111101001100",
56928 => "1111111101001100",
56929 => "1111111101001100",
56930 => "1111111101001100",
56931 => "1111111101001100",
56932 => "1111111101001100",
56933 => "1111111101001100",
56934 => "1111111101001100",
56935 => "1111111101001101",
56936 => "1111111101001101",
56937 => "1111111101001101",
56938 => "1111111101001101",
56939 => "1111111101001101",
56940 => "1111111101001101",
56941 => "1111111101001101",
56942 => "1111111101001101",
56943 => "1111111101001101",
56944 => "1111111101001101",
56945 => "1111111101001101",
56946 => "1111111101001101",
56947 => "1111111101001101",
56948 => "1111111101001101",
56949 => "1111111101001101",
56950 => "1111111101001101",
56951 => "1111111101001101",
56952 => "1111111101001101",
56953 => "1111111101001101",
56954 => "1111111101001101",
56955 => "1111111101001101",
56956 => "1111111101001101",
56957 => "1111111101001101",
56958 => "1111111101001110",
56959 => "1111111101001110",
56960 => "1111111101001110",
56961 => "1111111101001110",
56962 => "1111111101001110",
56963 => "1111111101001110",
56964 => "1111111101001110",
56965 => "1111111101001110",
56966 => "1111111101001110",
56967 => "1111111101001110",
56968 => "1111111101001110",
56969 => "1111111101001110",
56970 => "1111111101001110",
56971 => "1111111101001110",
56972 => "1111111101001110",
56973 => "1111111101001110",
56974 => "1111111101001110",
56975 => "1111111101001110",
56976 => "1111111101001110",
56977 => "1111111101001110",
56978 => "1111111101001110",
56979 => "1111111101001110",
56980 => "1111111101001110",
56981 => "1111111101001111",
56982 => "1111111101001111",
56983 => "1111111101001111",
56984 => "1111111101001111",
56985 => "1111111101001111",
56986 => "1111111101001111",
56987 => "1111111101001111",
56988 => "1111111101001111",
56989 => "1111111101001111",
56990 => "1111111101001111",
56991 => "1111111101001111",
56992 => "1111111101001111",
56993 => "1111111101001111",
56994 => "1111111101001111",
56995 => "1111111101001111",
56996 => "1111111101001111",
56997 => "1111111101001111",
56998 => "1111111101001111",
56999 => "1111111101001111",
57000 => "1111111101001111",
57001 => "1111111101001111",
57002 => "1111111101001111",
57003 => "1111111101001111",
57004 => "1111111101010000",
57005 => "1111111101010000",
57006 => "1111111101010000",
57007 => "1111111101010000",
57008 => "1111111101010000",
57009 => "1111111101010000",
57010 => "1111111101010000",
57011 => "1111111101010000",
57012 => "1111111101010000",
57013 => "1111111101010000",
57014 => "1111111101010000",
57015 => "1111111101010000",
57016 => "1111111101010000",
57017 => "1111111101010000",
57018 => "1111111101010000",
57019 => "1111111101010000",
57020 => "1111111101010000",
57021 => "1111111101010000",
57022 => "1111111101010000",
57023 => "1111111101010000",
57024 => "1111111101010000",
57025 => "1111111101010000",
57026 => "1111111101010000",
57027 => "1111111101010000",
57028 => "1111111101010001",
57029 => "1111111101010001",
57030 => "1111111101010001",
57031 => "1111111101010001",
57032 => "1111111101010001",
57033 => "1111111101010001",
57034 => "1111111101010001",
57035 => "1111111101010001",
57036 => "1111111101010001",
57037 => "1111111101010001",
57038 => "1111111101010001",
57039 => "1111111101010001",
57040 => "1111111101010001",
57041 => "1111111101010001",
57042 => "1111111101010001",
57043 => "1111111101010001",
57044 => "1111111101010001",
57045 => "1111111101010001",
57046 => "1111111101010001",
57047 => "1111111101010001",
57048 => "1111111101010001",
57049 => "1111111101010001",
57050 => "1111111101010001",
57051 => "1111111101010010",
57052 => "1111111101010010",
57053 => "1111111101010010",
57054 => "1111111101010010",
57055 => "1111111101010010",
57056 => "1111111101010010",
57057 => "1111111101010010",
57058 => "1111111101010010",
57059 => "1111111101010010",
57060 => "1111111101010010",
57061 => "1111111101010010",
57062 => "1111111101010010",
57063 => "1111111101010010",
57064 => "1111111101010010",
57065 => "1111111101010010",
57066 => "1111111101010010",
57067 => "1111111101010010",
57068 => "1111111101010010",
57069 => "1111111101010010",
57070 => "1111111101010010",
57071 => "1111111101010010",
57072 => "1111111101010010",
57073 => "1111111101010010",
57074 => "1111111101010010",
57075 => "1111111101010011",
57076 => "1111111101010011",
57077 => "1111111101010011",
57078 => "1111111101010011",
57079 => "1111111101010011",
57080 => "1111111101010011",
57081 => "1111111101010011",
57082 => "1111111101010011",
57083 => "1111111101010011",
57084 => "1111111101010011",
57085 => "1111111101010011",
57086 => "1111111101010011",
57087 => "1111111101010011",
57088 => "1111111101010011",
57089 => "1111111101010011",
57090 => "1111111101010011",
57091 => "1111111101010011",
57092 => "1111111101010011",
57093 => "1111111101010011",
57094 => "1111111101010011",
57095 => "1111111101010011",
57096 => "1111111101010011",
57097 => "1111111101010011",
57098 => "1111111101010011",
57099 => "1111111101010100",
57100 => "1111111101010100",
57101 => "1111111101010100",
57102 => "1111111101010100",
57103 => "1111111101010100",
57104 => "1111111101010100",
57105 => "1111111101010100",
57106 => "1111111101010100",
57107 => "1111111101010100",
57108 => "1111111101010100",
57109 => "1111111101010100",
57110 => "1111111101010100",
57111 => "1111111101010100",
57112 => "1111111101010100",
57113 => "1111111101010100",
57114 => "1111111101010100",
57115 => "1111111101010100",
57116 => "1111111101010100",
57117 => "1111111101010100",
57118 => "1111111101010100",
57119 => "1111111101010100",
57120 => "1111111101010100",
57121 => "1111111101010100",
57122 => "1111111101010100",
57123 => "1111111101010101",
57124 => "1111111101010101",
57125 => "1111111101010101",
57126 => "1111111101010101",
57127 => "1111111101010101",
57128 => "1111111101010101",
57129 => "1111111101010101",
57130 => "1111111101010101",
57131 => "1111111101010101",
57132 => "1111111101010101",
57133 => "1111111101010101",
57134 => "1111111101010101",
57135 => "1111111101010101",
57136 => "1111111101010101",
57137 => "1111111101010101",
57138 => "1111111101010101",
57139 => "1111111101010101",
57140 => "1111111101010101",
57141 => "1111111101010101",
57142 => "1111111101010101",
57143 => "1111111101010101",
57144 => "1111111101010101",
57145 => "1111111101010101",
57146 => "1111111101010101",
57147 => "1111111101010110",
57148 => "1111111101010110",
57149 => "1111111101010110",
57150 => "1111111101010110",
57151 => "1111111101010110",
57152 => "1111111101010110",
57153 => "1111111101010110",
57154 => "1111111101010110",
57155 => "1111111101010110",
57156 => "1111111101010110",
57157 => "1111111101010110",
57158 => "1111111101010110",
57159 => "1111111101010110",
57160 => "1111111101010110",
57161 => "1111111101010110",
57162 => "1111111101010110",
57163 => "1111111101010110",
57164 => "1111111101010110",
57165 => "1111111101010110",
57166 => "1111111101010110",
57167 => "1111111101010110",
57168 => "1111111101010110",
57169 => "1111111101010110",
57170 => "1111111101010110",
57171 => "1111111101010111",
57172 => "1111111101010111",
57173 => "1111111101010111",
57174 => "1111111101010111",
57175 => "1111111101010111",
57176 => "1111111101010111",
57177 => "1111111101010111",
57178 => "1111111101010111",
57179 => "1111111101010111",
57180 => "1111111101010111",
57181 => "1111111101010111",
57182 => "1111111101010111",
57183 => "1111111101010111",
57184 => "1111111101010111",
57185 => "1111111101010111",
57186 => "1111111101010111",
57187 => "1111111101010111",
57188 => "1111111101010111",
57189 => "1111111101010111",
57190 => "1111111101010111",
57191 => "1111111101010111",
57192 => "1111111101010111",
57193 => "1111111101010111",
57194 => "1111111101010111",
57195 => "1111111101011000",
57196 => "1111111101011000",
57197 => "1111111101011000",
57198 => "1111111101011000",
57199 => "1111111101011000",
57200 => "1111111101011000",
57201 => "1111111101011000",
57202 => "1111111101011000",
57203 => "1111111101011000",
57204 => "1111111101011000",
57205 => "1111111101011000",
57206 => "1111111101011000",
57207 => "1111111101011000",
57208 => "1111111101011000",
57209 => "1111111101011000",
57210 => "1111111101011000",
57211 => "1111111101011000",
57212 => "1111111101011000",
57213 => "1111111101011000",
57214 => "1111111101011000",
57215 => "1111111101011000",
57216 => "1111111101011000",
57217 => "1111111101011000",
57218 => "1111111101011000",
57219 => "1111111101011000",
57220 => "1111111101011001",
57221 => "1111111101011001",
57222 => "1111111101011001",
57223 => "1111111101011001",
57224 => "1111111101011001",
57225 => "1111111101011001",
57226 => "1111111101011001",
57227 => "1111111101011001",
57228 => "1111111101011001",
57229 => "1111111101011001",
57230 => "1111111101011001",
57231 => "1111111101011001",
57232 => "1111111101011001",
57233 => "1111111101011001",
57234 => "1111111101011001",
57235 => "1111111101011001",
57236 => "1111111101011001",
57237 => "1111111101011001",
57238 => "1111111101011001",
57239 => "1111111101011001",
57240 => "1111111101011001",
57241 => "1111111101011001",
57242 => "1111111101011001",
57243 => "1111111101011001",
57244 => "1111111101011001",
57245 => "1111111101011010",
57246 => "1111111101011010",
57247 => "1111111101011010",
57248 => "1111111101011010",
57249 => "1111111101011010",
57250 => "1111111101011010",
57251 => "1111111101011010",
57252 => "1111111101011010",
57253 => "1111111101011010",
57254 => "1111111101011010",
57255 => "1111111101011010",
57256 => "1111111101011010",
57257 => "1111111101011010",
57258 => "1111111101011010",
57259 => "1111111101011010",
57260 => "1111111101011010",
57261 => "1111111101011010",
57262 => "1111111101011010",
57263 => "1111111101011010",
57264 => "1111111101011010",
57265 => "1111111101011010",
57266 => "1111111101011010",
57267 => "1111111101011010",
57268 => "1111111101011010",
57269 => "1111111101011011",
57270 => "1111111101011011",
57271 => "1111111101011011",
57272 => "1111111101011011",
57273 => "1111111101011011",
57274 => "1111111101011011",
57275 => "1111111101011011",
57276 => "1111111101011011",
57277 => "1111111101011011",
57278 => "1111111101011011",
57279 => "1111111101011011",
57280 => "1111111101011011",
57281 => "1111111101011011",
57282 => "1111111101011011",
57283 => "1111111101011011",
57284 => "1111111101011011",
57285 => "1111111101011011",
57286 => "1111111101011011",
57287 => "1111111101011011",
57288 => "1111111101011011",
57289 => "1111111101011011",
57290 => "1111111101011011",
57291 => "1111111101011011",
57292 => "1111111101011011",
57293 => "1111111101011011",
57294 => "1111111101011100",
57295 => "1111111101011100",
57296 => "1111111101011100",
57297 => "1111111101011100",
57298 => "1111111101011100",
57299 => "1111111101011100",
57300 => "1111111101011100",
57301 => "1111111101011100",
57302 => "1111111101011100",
57303 => "1111111101011100",
57304 => "1111111101011100",
57305 => "1111111101011100",
57306 => "1111111101011100",
57307 => "1111111101011100",
57308 => "1111111101011100",
57309 => "1111111101011100",
57310 => "1111111101011100",
57311 => "1111111101011100",
57312 => "1111111101011100",
57313 => "1111111101011100",
57314 => "1111111101011100",
57315 => "1111111101011100",
57316 => "1111111101011100",
57317 => "1111111101011100",
57318 => "1111111101011100",
57319 => "1111111101011100",
57320 => "1111111101011101",
57321 => "1111111101011101",
57322 => "1111111101011101",
57323 => "1111111101011101",
57324 => "1111111101011101",
57325 => "1111111101011101",
57326 => "1111111101011101",
57327 => "1111111101011101",
57328 => "1111111101011101",
57329 => "1111111101011101",
57330 => "1111111101011101",
57331 => "1111111101011101",
57332 => "1111111101011101",
57333 => "1111111101011101",
57334 => "1111111101011101",
57335 => "1111111101011101",
57336 => "1111111101011101",
57337 => "1111111101011101",
57338 => "1111111101011101",
57339 => "1111111101011101",
57340 => "1111111101011101",
57341 => "1111111101011101",
57342 => "1111111101011101",
57343 => "1111111101011101",
57344 => "1111111101011101",
57345 => "1111111101011110",
57346 => "1111111101011110",
57347 => "1111111101011110",
57348 => "1111111101011110",
57349 => "1111111101011110",
57350 => "1111111101011110",
57351 => "1111111101011110",
57352 => "1111111101011110",
57353 => "1111111101011110",
57354 => "1111111101011110",
57355 => "1111111101011110",
57356 => "1111111101011110",
57357 => "1111111101011110",
57358 => "1111111101011110",
57359 => "1111111101011110",
57360 => "1111111101011110",
57361 => "1111111101011110",
57362 => "1111111101011110",
57363 => "1111111101011110",
57364 => "1111111101011110",
57365 => "1111111101011110",
57366 => "1111111101011110",
57367 => "1111111101011110",
57368 => "1111111101011110",
57369 => "1111111101011110",
57370 => "1111111101011111",
57371 => "1111111101011111",
57372 => "1111111101011111",
57373 => "1111111101011111",
57374 => "1111111101011111",
57375 => "1111111101011111",
57376 => "1111111101011111",
57377 => "1111111101011111",
57378 => "1111111101011111",
57379 => "1111111101011111",
57380 => "1111111101011111",
57381 => "1111111101011111",
57382 => "1111111101011111",
57383 => "1111111101011111",
57384 => "1111111101011111",
57385 => "1111111101011111",
57386 => "1111111101011111",
57387 => "1111111101011111",
57388 => "1111111101011111",
57389 => "1111111101011111",
57390 => "1111111101011111",
57391 => "1111111101011111",
57392 => "1111111101011111",
57393 => "1111111101011111",
57394 => "1111111101011111",
57395 => "1111111101011111",
57396 => "1111111101100000",
57397 => "1111111101100000",
57398 => "1111111101100000",
57399 => "1111111101100000",
57400 => "1111111101100000",
57401 => "1111111101100000",
57402 => "1111111101100000",
57403 => "1111111101100000",
57404 => "1111111101100000",
57405 => "1111111101100000",
57406 => "1111111101100000",
57407 => "1111111101100000",
57408 => "1111111101100000",
57409 => "1111111101100000",
57410 => "1111111101100000",
57411 => "1111111101100000",
57412 => "1111111101100000",
57413 => "1111111101100000",
57414 => "1111111101100000",
57415 => "1111111101100000",
57416 => "1111111101100000",
57417 => "1111111101100000",
57418 => "1111111101100000",
57419 => "1111111101100000",
57420 => "1111111101100000",
57421 => "1111111101100000",
57422 => "1111111101100001",
57423 => "1111111101100001",
57424 => "1111111101100001",
57425 => "1111111101100001",
57426 => "1111111101100001",
57427 => "1111111101100001",
57428 => "1111111101100001",
57429 => "1111111101100001",
57430 => "1111111101100001",
57431 => "1111111101100001",
57432 => "1111111101100001",
57433 => "1111111101100001",
57434 => "1111111101100001",
57435 => "1111111101100001",
57436 => "1111111101100001",
57437 => "1111111101100001",
57438 => "1111111101100001",
57439 => "1111111101100001",
57440 => "1111111101100001",
57441 => "1111111101100001",
57442 => "1111111101100001",
57443 => "1111111101100001",
57444 => "1111111101100001",
57445 => "1111111101100001",
57446 => "1111111101100001",
57447 => "1111111101100010",
57448 => "1111111101100010",
57449 => "1111111101100010",
57450 => "1111111101100010",
57451 => "1111111101100010",
57452 => "1111111101100010",
57453 => "1111111101100010",
57454 => "1111111101100010",
57455 => "1111111101100010",
57456 => "1111111101100010",
57457 => "1111111101100010",
57458 => "1111111101100010",
57459 => "1111111101100010",
57460 => "1111111101100010",
57461 => "1111111101100010",
57462 => "1111111101100010",
57463 => "1111111101100010",
57464 => "1111111101100010",
57465 => "1111111101100010",
57466 => "1111111101100010",
57467 => "1111111101100010",
57468 => "1111111101100010",
57469 => "1111111101100010",
57470 => "1111111101100010",
57471 => "1111111101100010",
57472 => "1111111101100010",
57473 => "1111111101100010",
57474 => "1111111101100011",
57475 => "1111111101100011",
57476 => "1111111101100011",
57477 => "1111111101100011",
57478 => "1111111101100011",
57479 => "1111111101100011",
57480 => "1111111101100011",
57481 => "1111111101100011",
57482 => "1111111101100011",
57483 => "1111111101100011",
57484 => "1111111101100011",
57485 => "1111111101100011",
57486 => "1111111101100011",
57487 => "1111111101100011",
57488 => "1111111101100011",
57489 => "1111111101100011",
57490 => "1111111101100011",
57491 => "1111111101100011",
57492 => "1111111101100011",
57493 => "1111111101100011",
57494 => "1111111101100011",
57495 => "1111111101100011",
57496 => "1111111101100011",
57497 => "1111111101100011",
57498 => "1111111101100011",
57499 => "1111111101100011",
57500 => "1111111101100100",
57501 => "1111111101100100",
57502 => "1111111101100100",
57503 => "1111111101100100",
57504 => "1111111101100100",
57505 => "1111111101100100",
57506 => "1111111101100100",
57507 => "1111111101100100",
57508 => "1111111101100100",
57509 => "1111111101100100",
57510 => "1111111101100100",
57511 => "1111111101100100",
57512 => "1111111101100100",
57513 => "1111111101100100",
57514 => "1111111101100100",
57515 => "1111111101100100",
57516 => "1111111101100100",
57517 => "1111111101100100",
57518 => "1111111101100100",
57519 => "1111111101100100",
57520 => "1111111101100100",
57521 => "1111111101100100",
57522 => "1111111101100100",
57523 => "1111111101100100",
57524 => "1111111101100100",
57525 => "1111111101100100",
57526 => "1111111101100101",
57527 => "1111111101100101",
57528 => "1111111101100101",
57529 => "1111111101100101",
57530 => "1111111101100101",
57531 => "1111111101100101",
57532 => "1111111101100101",
57533 => "1111111101100101",
57534 => "1111111101100101",
57535 => "1111111101100101",
57536 => "1111111101100101",
57537 => "1111111101100101",
57538 => "1111111101100101",
57539 => "1111111101100101",
57540 => "1111111101100101",
57541 => "1111111101100101",
57542 => "1111111101100101",
57543 => "1111111101100101",
57544 => "1111111101100101",
57545 => "1111111101100101",
57546 => "1111111101100101",
57547 => "1111111101100101",
57548 => "1111111101100101",
57549 => "1111111101100101",
57550 => "1111111101100101",
57551 => "1111111101100101",
57552 => "1111111101100101",
57553 => "1111111101100110",
57554 => "1111111101100110",
57555 => "1111111101100110",
57556 => "1111111101100110",
57557 => "1111111101100110",
57558 => "1111111101100110",
57559 => "1111111101100110",
57560 => "1111111101100110",
57561 => "1111111101100110",
57562 => "1111111101100110",
57563 => "1111111101100110",
57564 => "1111111101100110",
57565 => "1111111101100110",
57566 => "1111111101100110",
57567 => "1111111101100110",
57568 => "1111111101100110",
57569 => "1111111101100110",
57570 => "1111111101100110",
57571 => "1111111101100110",
57572 => "1111111101100110",
57573 => "1111111101100110",
57574 => "1111111101100110",
57575 => "1111111101100110",
57576 => "1111111101100110",
57577 => "1111111101100110",
57578 => "1111111101100110",
57579 => "1111111101100111",
57580 => "1111111101100111",
57581 => "1111111101100111",
57582 => "1111111101100111",
57583 => "1111111101100111",
57584 => "1111111101100111",
57585 => "1111111101100111",
57586 => "1111111101100111",
57587 => "1111111101100111",
57588 => "1111111101100111",
57589 => "1111111101100111",
57590 => "1111111101100111",
57591 => "1111111101100111",
57592 => "1111111101100111",
57593 => "1111111101100111",
57594 => "1111111101100111",
57595 => "1111111101100111",
57596 => "1111111101100111",
57597 => "1111111101100111",
57598 => "1111111101100111",
57599 => "1111111101100111",
57600 => "1111111101100111",
57601 => "1111111101100111",
57602 => "1111111101100111",
57603 => "1111111101100111",
57604 => "1111111101100111",
57605 => "1111111101100111",
57606 => "1111111101101000",
57607 => "1111111101101000",
57608 => "1111111101101000",
57609 => "1111111101101000",
57610 => "1111111101101000",
57611 => "1111111101101000",
57612 => "1111111101101000",
57613 => "1111111101101000",
57614 => "1111111101101000",
57615 => "1111111101101000",
57616 => "1111111101101000",
57617 => "1111111101101000",
57618 => "1111111101101000",
57619 => "1111111101101000",
57620 => "1111111101101000",
57621 => "1111111101101000",
57622 => "1111111101101000",
57623 => "1111111101101000",
57624 => "1111111101101000",
57625 => "1111111101101000",
57626 => "1111111101101000",
57627 => "1111111101101000",
57628 => "1111111101101000",
57629 => "1111111101101000",
57630 => "1111111101101000",
57631 => "1111111101101000",
57632 => "1111111101101000",
57633 => "1111111101101001",
57634 => "1111111101101001",
57635 => "1111111101101001",
57636 => "1111111101101001",
57637 => "1111111101101001",
57638 => "1111111101101001",
57639 => "1111111101101001",
57640 => "1111111101101001",
57641 => "1111111101101001",
57642 => "1111111101101001",
57643 => "1111111101101001",
57644 => "1111111101101001",
57645 => "1111111101101001",
57646 => "1111111101101001",
57647 => "1111111101101001",
57648 => "1111111101101001",
57649 => "1111111101101001",
57650 => "1111111101101001",
57651 => "1111111101101001",
57652 => "1111111101101001",
57653 => "1111111101101001",
57654 => "1111111101101001",
57655 => "1111111101101001",
57656 => "1111111101101001",
57657 => "1111111101101001",
57658 => "1111111101101001",
57659 => "1111111101101001",
57660 => "1111111101101001",
57661 => "1111111101101010",
57662 => "1111111101101010",
57663 => "1111111101101010",
57664 => "1111111101101010",
57665 => "1111111101101010",
57666 => "1111111101101010",
57667 => "1111111101101010",
57668 => "1111111101101010",
57669 => "1111111101101010",
57670 => "1111111101101010",
57671 => "1111111101101010",
57672 => "1111111101101010",
57673 => "1111111101101010",
57674 => "1111111101101010",
57675 => "1111111101101010",
57676 => "1111111101101010",
57677 => "1111111101101010",
57678 => "1111111101101010",
57679 => "1111111101101010",
57680 => "1111111101101010",
57681 => "1111111101101010",
57682 => "1111111101101010",
57683 => "1111111101101010",
57684 => "1111111101101010",
57685 => "1111111101101010",
57686 => "1111111101101010",
57687 => "1111111101101010",
57688 => "1111111101101011",
57689 => "1111111101101011",
57690 => "1111111101101011",
57691 => "1111111101101011",
57692 => "1111111101101011",
57693 => "1111111101101011",
57694 => "1111111101101011",
57695 => "1111111101101011",
57696 => "1111111101101011",
57697 => "1111111101101011",
57698 => "1111111101101011",
57699 => "1111111101101011",
57700 => "1111111101101011",
57701 => "1111111101101011",
57702 => "1111111101101011",
57703 => "1111111101101011",
57704 => "1111111101101011",
57705 => "1111111101101011",
57706 => "1111111101101011",
57707 => "1111111101101011",
57708 => "1111111101101011",
57709 => "1111111101101011",
57710 => "1111111101101011",
57711 => "1111111101101011",
57712 => "1111111101101011",
57713 => "1111111101101011",
57714 => "1111111101101011",
57715 => "1111111101101011",
57716 => "1111111101101100",
57717 => "1111111101101100",
57718 => "1111111101101100",
57719 => "1111111101101100",
57720 => "1111111101101100",
57721 => "1111111101101100",
57722 => "1111111101101100",
57723 => "1111111101101100",
57724 => "1111111101101100",
57725 => "1111111101101100",
57726 => "1111111101101100",
57727 => "1111111101101100",
57728 => "1111111101101100",
57729 => "1111111101101100",
57730 => "1111111101101100",
57731 => "1111111101101100",
57732 => "1111111101101100",
57733 => "1111111101101100",
57734 => "1111111101101100",
57735 => "1111111101101100",
57736 => "1111111101101100",
57737 => "1111111101101100",
57738 => "1111111101101100",
57739 => "1111111101101100",
57740 => "1111111101101100",
57741 => "1111111101101100",
57742 => "1111111101101100",
57743 => "1111111101101100",
57744 => "1111111101101101",
57745 => "1111111101101101",
57746 => "1111111101101101",
57747 => "1111111101101101",
57748 => "1111111101101101",
57749 => "1111111101101101",
57750 => "1111111101101101",
57751 => "1111111101101101",
57752 => "1111111101101101",
57753 => "1111111101101101",
57754 => "1111111101101101",
57755 => "1111111101101101",
57756 => "1111111101101101",
57757 => "1111111101101101",
57758 => "1111111101101101",
57759 => "1111111101101101",
57760 => "1111111101101101",
57761 => "1111111101101101",
57762 => "1111111101101101",
57763 => "1111111101101101",
57764 => "1111111101101101",
57765 => "1111111101101101",
57766 => "1111111101101101",
57767 => "1111111101101101",
57768 => "1111111101101101",
57769 => "1111111101101101",
57770 => "1111111101101101",
57771 => "1111111101101101",
57772 => "1111111101101110",
57773 => "1111111101101110",
57774 => "1111111101101110",
57775 => "1111111101101110",
57776 => "1111111101101110",
57777 => "1111111101101110",
57778 => "1111111101101110",
57779 => "1111111101101110",
57780 => "1111111101101110",
57781 => "1111111101101110",
57782 => "1111111101101110",
57783 => "1111111101101110",
57784 => "1111111101101110",
57785 => "1111111101101110",
57786 => "1111111101101110",
57787 => "1111111101101110",
57788 => "1111111101101110",
57789 => "1111111101101110",
57790 => "1111111101101110",
57791 => "1111111101101110",
57792 => "1111111101101110",
57793 => "1111111101101110",
57794 => "1111111101101110",
57795 => "1111111101101110",
57796 => "1111111101101110",
57797 => "1111111101101110",
57798 => "1111111101101110",
57799 => "1111111101101110",
57800 => "1111111101101111",
57801 => "1111111101101111",
57802 => "1111111101101111",
57803 => "1111111101101111",
57804 => "1111111101101111",
57805 => "1111111101101111",
57806 => "1111111101101111",
57807 => "1111111101101111",
57808 => "1111111101101111",
57809 => "1111111101101111",
57810 => "1111111101101111",
57811 => "1111111101101111",
57812 => "1111111101101111",
57813 => "1111111101101111",
57814 => "1111111101101111",
57815 => "1111111101101111",
57816 => "1111111101101111",
57817 => "1111111101101111",
57818 => "1111111101101111",
57819 => "1111111101101111",
57820 => "1111111101101111",
57821 => "1111111101101111",
57822 => "1111111101101111",
57823 => "1111111101101111",
57824 => "1111111101101111",
57825 => "1111111101101111",
57826 => "1111111101101111",
57827 => "1111111101101111",
57828 => "1111111101110000",
57829 => "1111111101110000",
57830 => "1111111101110000",
57831 => "1111111101110000",
57832 => "1111111101110000",
57833 => "1111111101110000",
57834 => "1111111101110000",
57835 => "1111111101110000",
57836 => "1111111101110000",
57837 => "1111111101110000",
57838 => "1111111101110000",
57839 => "1111111101110000",
57840 => "1111111101110000",
57841 => "1111111101110000",
57842 => "1111111101110000",
57843 => "1111111101110000",
57844 => "1111111101110000",
57845 => "1111111101110000",
57846 => "1111111101110000",
57847 => "1111111101110000",
57848 => "1111111101110000",
57849 => "1111111101110000",
57850 => "1111111101110000",
57851 => "1111111101110000",
57852 => "1111111101110000",
57853 => "1111111101110000",
57854 => "1111111101110000",
57855 => "1111111101110000",
57856 => "1111111101110000",
57857 => "1111111101110001",
57858 => "1111111101110001",
57859 => "1111111101110001",
57860 => "1111111101110001",
57861 => "1111111101110001",
57862 => "1111111101110001",
57863 => "1111111101110001",
57864 => "1111111101110001",
57865 => "1111111101110001",
57866 => "1111111101110001",
57867 => "1111111101110001",
57868 => "1111111101110001",
57869 => "1111111101110001",
57870 => "1111111101110001",
57871 => "1111111101110001",
57872 => "1111111101110001",
57873 => "1111111101110001",
57874 => "1111111101110001",
57875 => "1111111101110001",
57876 => "1111111101110001",
57877 => "1111111101110001",
57878 => "1111111101110001",
57879 => "1111111101110001",
57880 => "1111111101110001",
57881 => "1111111101110001",
57882 => "1111111101110001",
57883 => "1111111101110001",
57884 => "1111111101110001",
57885 => "1111111101110001",
57886 => "1111111101110010",
57887 => "1111111101110010",
57888 => "1111111101110010",
57889 => "1111111101110010",
57890 => "1111111101110010",
57891 => "1111111101110010",
57892 => "1111111101110010",
57893 => "1111111101110010",
57894 => "1111111101110010",
57895 => "1111111101110010",
57896 => "1111111101110010",
57897 => "1111111101110010",
57898 => "1111111101110010",
57899 => "1111111101110010",
57900 => "1111111101110010",
57901 => "1111111101110010",
57902 => "1111111101110010",
57903 => "1111111101110010",
57904 => "1111111101110010",
57905 => "1111111101110010",
57906 => "1111111101110010",
57907 => "1111111101110010",
57908 => "1111111101110010",
57909 => "1111111101110010",
57910 => "1111111101110010",
57911 => "1111111101110010",
57912 => "1111111101110010",
57913 => "1111111101110010",
57914 => "1111111101110010",
57915 => "1111111101110011",
57916 => "1111111101110011",
57917 => "1111111101110011",
57918 => "1111111101110011",
57919 => "1111111101110011",
57920 => "1111111101110011",
57921 => "1111111101110011",
57922 => "1111111101110011",
57923 => "1111111101110011",
57924 => "1111111101110011",
57925 => "1111111101110011",
57926 => "1111111101110011",
57927 => "1111111101110011",
57928 => "1111111101110011",
57929 => "1111111101110011",
57930 => "1111111101110011",
57931 => "1111111101110011",
57932 => "1111111101110011",
57933 => "1111111101110011",
57934 => "1111111101110011",
57935 => "1111111101110011",
57936 => "1111111101110011",
57937 => "1111111101110011",
57938 => "1111111101110011",
57939 => "1111111101110011",
57940 => "1111111101110011",
57941 => "1111111101110011",
57942 => "1111111101110011",
57943 => "1111111101110011",
57944 => "1111111101110100",
57945 => "1111111101110100",
57946 => "1111111101110100",
57947 => "1111111101110100",
57948 => "1111111101110100",
57949 => "1111111101110100",
57950 => "1111111101110100",
57951 => "1111111101110100",
57952 => "1111111101110100",
57953 => "1111111101110100",
57954 => "1111111101110100",
57955 => "1111111101110100",
57956 => "1111111101110100",
57957 => "1111111101110100",
57958 => "1111111101110100",
57959 => "1111111101110100",
57960 => "1111111101110100",
57961 => "1111111101110100",
57962 => "1111111101110100",
57963 => "1111111101110100",
57964 => "1111111101110100",
57965 => "1111111101110100",
57966 => "1111111101110100",
57967 => "1111111101110100",
57968 => "1111111101110100",
57969 => "1111111101110100",
57970 => "1111111101110100",
57971 => "1111111101110100",
57972 => "1111111101110100",
57973 => "1111111101110101",
57974 => "1111111101110101",
57975 => "1111111101110101",
57976 => "1111111101110101",
57977 => "1111111101110101",
57978 => "1111111101110101",
57979 => "1111111101110101",
57980 => "1111111101110101",
57981 => "1111111101110101",
57982 => "1111111101110101",
57983 => "1111111101110101",
57984 => "1111111101110101",
57985 => "1111111101110101",
57986 => "1111111101110101",
57987 => "1111111101110101",
57988 => "1111111101110101",
57989 => "1111111101110101",
57990 => "1111111101110101",
57991 => "1111111101110101",
57992 => "1111111101110101",
57993 => "1111111101110101",
57994 => "1111111101110101",
57995 => "1111111101110101",
57996 => "1111111101110101",
57997 => "1111111101110101",
57998 => "1111111101110101",
57999 => "1111111101110101",
58000 => "1111111101110101",
58001 => "1111111101110101",
58002 => "1111111101110101",
58003 => "1111111101110110",
58004 => "1111111101110110",
58005 => "1111111101110110",
58006 => "1111111101110110",
58007 => "1111111101110110",
58008 => "1111111101110110",
58009 => "1111111101110110",
58010 => "1111111101110110",
58011 => "1111111101110110",
58012 => "1111111101110110",
58013 => "1111111101110110",
58014 => "1111111101110110",
58015 => "1111111101110110",
58016 => "1111111101110110",
58017 => "1111111101110110",
58018 => "1111111101110110",
58019 => "1111111101110110",
58020 => "1111111101110110",
58021 => "1111111101110110",
58022 => "1111111101110110",
58023 => "1111111101110110",
58024 => "1111111101110110",
58025 => "1111111101110110",
58026 => "1111111101110110",
58027 => "1111111101110110",
58028 => "1111111101110110",
58029 => "1111111101110110",
58030 => "1111111101110110",
58031 => "1111111101110110",
58032 => "1111111101110110",
58033 => "1111111101110111",
58034 => "1111111101110111",
58035 => "1111111101110111",
58036 => "1111111101110111",
58037 => "1111111101110111",
58038 => "1111111101110111",
58039 => "1111111101110111",
58040 => "1111111101110111",
58041 => "1111111101110111",
58042 => "1111111101110111",
58043 => "1111111101110111",
58044 => "1111111101110111",
58045 => "1111111101110111",
58046 => "1111111101110111",
58047 => "1111111101110111",
58048 => "1111111101110111",
58049 => "1111111101110111",
58050 => "1111111101110111",
58051 => "1111111101110111",
58052 => "1111111101110111",
58053 => "1111111101110111",
58054 => "1111111101110111",
58055 => "1111111101110111",
58056 => "1111111101110111",
58057 => "1111111101110111",
58058 => "1111111101110111",
58059 => "1111111101110111",
58060 => "1111111101110111",
58061 => "1111111101110111",
58062 => "1111111101110111",
58063 => "1111111101111000",
58064 => "1111111101111000",
58065 => "1111111101111000",
58066 => "1111111101111000",
58067 => "1111111101111000",
58068 => "1111111101111000",
58069 => "1111111101111000",
58070 => "1111111101111000",
58071 => "1111111101111000",
58072 => "1111111101111000",
58073 => "1111111101111000",
58074 => "1111111101111000",
58075 => "1111111101111000",
58076 => "1111111101111000",
58077 => "1111111101111000",
58078 => "1111111101111000",
58079 => "1111111101111000",
58080 => "1111111101111000",
58081 => "1111111101111000",
58082 => "1111111101111000",
58083 => "1111111101111000",
58084 => "1111111101111000",
58085 => "1111111101111000",
58086 => "1111111101111000",
58087 => "1111111101111000",
58088 => "1111111101111000",
58089 => "1111111101111000",
58090 => "1111111101111000",
58091 => "1111111101111000",
58092 => "1111111101111000",
58093 => "1111111101111001",
58094 => "1111111101111001",
58095 => "1111111101111001",
58096 => "1111111101111001",
58097 => "1111111101111001",
58098 => "1111111101111001",
58099 => "1111111101111001",
58100 => "1111111101111001",
58101 => "1111111101111001",
58102 => "1111111101111001",
58103 => "1111111101111001",
58104 => "1111111101111001",
58105 => "1111111101111001",
58106 => "1111111101111001",
58107 => "1111111101111001",
58108 => "1111111101111001",
58109 => "1111111101111001",
58110 => "1111111101111001",
58111 => "1111111101111001",
58112 => "1111111101111001",
58113 => "1111111101111001",
58114 => "1111111101111001",
58115 => "1111111101111001",
58116 => "1111111101111001",
58117 => "1111111101111001",
58118 => "1111111101111001",
58119 => "1111111101111001",
58120 => "1111111101111001",
58121 => "1111111101111001",
58122 => "1111111101111001",
58123 => "1111111101111001",
58124 => "1111111101111010",
58125 => "1111111101111010",
58126 => "1111111101111010",
58127 => "1111111101111010",
58128 => "1111111101111010",
58129 => "1111111101111010",
58130 => "1111111101111010",
58131 => "1111111101111010",
58132 => "1111111101111010",
58133 => "1111111101111010",
58134 => "1111111101111010",
58135 => "1111111101111010",
58136 => "1111111101111010",
58137 => "1111111101111010",
58138 => "1111111101111010",
58139 => "1111111101111010",
58140 => "1111111101111010",
58141 => "1111111101111010",
58142 => "1111111101111010",
58143 => "1111111101111010",
58144 => "1111111101111010",
58145 => "1111111101111010",
58146 => "1111111101111010",
58147 => "1111111101111010",
58148 => "1111111101111010",
58149 => "1111111101111010",
58150 => "1111111101111010",
58151 => "1111111101111010",
58152 => "1111111101111010",
58153 => "1111111101111010",
58154 => "1111111101111010",
58155 => "1111111101111011",
58156 => "1111111101111011",
58157 => "1111111101111011",
58158 => "1111111101111011",
58159 => "1111111101111011",
58160 => "1111111101111011",
58161 => "1111111101111011",
58162 => "1111111101111011",
58163 => "1111111101111011",
58164 => "1111111101111011",
58165 => "1111111101111011",
58166 => "1111111101111011",
58167 => "1111111101111011",
58168 => "1111111101111011",
58169 => "1111111101111011",
58170 => "1111111101111011",
58171 => "1111111101111011",
58172 => "1111111101111011",
58173 => "1111111101111011",
58174 => "1111111101111011",
58175 => "1111111101111011",
58176 => "1111111101111011",
58177 => "1111111101111011",
58178 => "1111111101111011",
58179 => "1111111101111011",
58180 => "1111111101111011",
58181 => "1111111101111011",
58182 => "1111111101111011",
58183 => "1111111101111011",
58184 => "1111111101111011",
58185 => "1111111101111100",
58186 => "1111111101111100",
58187 => "1111111101111100",
58188 => "1111111101111100",
58189 => "1111111101111100",
58190 => "1111111101111100",
58191 => "1111111101111100",
58192 => "1111111101111100",
58193 => "1111111101111100",
58194 => "1111111101111100",
58195 => "1111111101111100",
58196 => "1111111101111100",
58197 => "1111111101111100",
58198 => "1111111101111100",
58199 => "1111111101111100",
58200 => "1111111101111100",
58201 => "1111111101111100",
58202 => "1111111101111100",
58203 => "1111111101111100",
58204 => "1111111101111100",
58205 => "1111111101111100",
58206 => "1111111101111100",
58207 => "1111111101111100",
58208 => "1111111101111100",
58209 => "1111111101111100",
58210 => "1111111101111100",
58211 => "1111111101111100",
58212 => "1111111101111100",
58213 => "1111111101111100",
58214 => "1111111101111100",
58215 => "1111111101111100",
58216 => "1111111101111100",
58217 => "1111111101111101",
58218 => "1111111101111101",
58219 => "1111111101111101",
58220 => "1111111101111101",
58221 => "1111111101111101",
58222 => "1111111101111101",
58223 => "1111111101111101",
58224 => "1111111101111101",
58225 => "1111111101111101",
58226 => "1111111101111101",
58227 => "1111111101111101",
58228 => "1111111101111101",
58229 => "1111111101111101",
58230 => "1111111101111101",
58231 => "1111111101111101",
58232 => "1111111101111101",
58233 => "1111111101111101",
58234 => "1111111101111101",
58235 => "1111111101111101",
58236 => "1111111101111101",
58237 => "1111111101111101",
58238 => "1111111101111101",
58239 => "1111111101111101",
58240 => "1111111101111101",
58241 => "1111111101111101",
58242 => "1111111101111101",
58243 => "1111111101111101",
58244 => "1111111101111101",
58245 => "1111111101111101",
58246 => "1111111101111101",
58247 => "1111111101111101",
58248 => "1111111101111110",
58249 => "1111111101111110",
58250 => "1111111101111110",
58251 => "1111111101111110",
58252 => "1111111101111110",
58253 => "1111111101111110",
58254 => "1111111101111110",
58255 => "1111111101111110",
58256 => "1111111101111110",
58257 => "1111111101111110",
58258 => "1111111101111110",
58259 => "1111111101111110",
58260 => "1111111101111110",
58261 => "1111111101111110",
58262 => "1111111101111110",
58263 => "1111111101111110",
58264 => "1111111101111110",
58265 => "1111111101111110",
58266 => "1111111101111110",
58267 => "1111111101111110",
58268 => "1111111101111110",
58269 => "1111111101111110",
58270 => "1111111101111110",
58271 => "1111111101111110",
58272 => "1111111101111110",
58273 => "1111111101111110",
58274 => "1111111101111110",
58275 => "1111111101111110",
58276 => "1111111101111110",
58277 => "1111111101111110",
58278 => "1111111101111110",
58279 => "1111111101111110",
58280 => "1111111101111111",
58281 => "1111111101111111",
58282 => "1111111101111111",
58283 => "1111111101111111",
58284 => "1111111101111111",
58285 => "1111111101111111",
58286 => "1111111101111111",
58287 => "1111111101111111",
58288 => "1111111101111111",
58289 => "1111111101111111",
58290 => "1111111101111111",
58291 => "1111111101111111",
58292 => "1111111101111111",
58293 => "1111111101111111",
58294 => "1111111101111111",
58295 => "1111111101111111",
58296 => "1111111101111111",
58297 => "1111111101111111",
58298 => "1111111101111111",
58299 => "1111111101111111",
58300 => "1111111101111111",
58301 => "1111111101111111",
58302 => "1111111101111111",
58303 => "1111111101111111",
58304 => "1111111101111111",
58305 => "1111111101111111",
58306 => "1111111101111111",
58307 => "1111111101111111",
58308 => "1111111101111111",
58309 => "1111111101111111",
58310 => "1111111101111111",
58311 => "1111111101111111",
58312 => "1111111110000000",
58313 => "1111111110000000",
58314 => "1111111110000000",
58315 => "1111111110000000",
58316 => "1111111110000000",
58317 => "1111111110000000",
58318 => "1111111110000000",
58319 => "1111111110000000",
58320 => "1111111110000000",
58321 => "1111111110000000",
58322 => "1111111110000000",
58323 => "1111111110000000",
58324 => "1111111110000000",
58325 => "1111111110000000",
58326 => "1111111110000000",
58327 => "1111111110000000",
58328 => "1111111110000000",
58329 => "1111111110000000",
58330 => "1111111110000000",
58331 => "1111111110000000",
58332 => "1111111110000000",
58333 => "1111111110000000",
58334 => "1111111110000000",
58335 => "1111111110000000",
58336 => "1111111110000000",
58337 => "1111111110000000",
58338 => "1111111110000000",
58339 => "1111111110000000",
58340 => "1111111110000000",
58341 => "1111111110000000",
58342 => "1111111110000000",
58343 => "1111111110000000",
58344 => "1111111110000001",
58345 => "1111111110000001",
58346 => "1111111110000001",
58347 => "1111111110000001",
58348 => "1111111110000001",
58349 => "1111111110000001",
58350 => "1111111110000001",
58351 => "1111111110000001",
58352 => "1111111110000001",
58353 => "1111111110000001",
58354 => "1111111110000001",
58355 => "1111111110000001",
58356 => "1111111110000001",
58357 => "1111111110000001",
58358 => "1111111110000001",
58359 => "1111111110000001",
58360 => "1111111110000001",
58361 => "1111111110000001",
58362 => "1111111110000001",
58363 => "1111111110000001",
58364 => "1111111110000001",
58365 => "1111111110000001",
58366 => "1111111110000001",
58367 => "1111111110000001",
58368 => "1111111110000001",
58369 => "1111111110000001",
58370 => "1111111110000001",
58371 => "1111111110000001",
58372 => "1111111110000001",
58373 => "1111111110000001",
58374 => "1111111110000001",
58375 => "1111111110000001",
58376 => "1111111110000010",
58377 => "1111111110000010",
58378 => "1111111110000010",
58379 => "1111111110000010",
58380 => "1111111110000010",
58381 => "1111111110000010",
58382 => "1111111110000010",
58383 => "1111111110000010",
58384 => "1111111110000010",
58385 => "1111111110000010",
58386 => "1111111110000010",
58387 => "1111111110000010",
58388 => "1111111110000010",
58389 => "1111111110000010",
58390 => "1111111110000010",
58391 => "1111111110000010",
58392 => "1111111110000010",
58393 => "1111111110000010",
58394 => "1111111110000010",
58395 => "1111111110000010",
58396 => "1111111110000010",
58397 => "1111111110000010",
58398 => "1111111110000010",
58399 => "1111111110000010",
58400 => "1111111110000010",
58401 => "1111111110000010",
58402 => "1111111110000010",
58403 => "1111111110000010",
58404 => "1111111110000010",
58405 => "1111111110000010",
58406 => "1111111110000010",
58407 => "1111111110000010",
58408 => "1111111110000010",
58409 => "1111111110000011",
58410 => "1111111110000011",
58411 => "1111111110000011",
58412 => "1111111110000011",
58413 => "1111111110000011",
58414 => "1111111110000011",
58415 => "1111111110000011",
58416 => "1111111110000011",
58417 => "1111111110000011",
58418 => "1111111110000011",
58419 => "1111111110000011",
58420 => "1111111110000011",
58421 => "1111111110000011",
58422 => "1111111110000011",
58423 => "1111111110000011",
58424 => "1111111110000011",
58425 => "1111111110000011",
58426 => "1111111110000011",
58427 => "1111111110000011",
58428 => "1111111110000011",
58429 => "1111111110000011",
58430 => "1111111110000011",
58431 => "1111111110000011",
58432 => "1111111110000011",
58433 => "1111111110000011",
58434 => "1111111110000011",
58435 => "1111111110000011",
58436 => "1111111110000011",
58437 => "1111111110000011",
58438 => "1111111110000011",
58439 => "1111111110000011",
58440 => "1111111110000011",
58441 => "1111111110000011",
58442 => "1111111110000100",
58443 => "1111111110000100",
58444 => "1111111110000100",
58445 => "1111111110000100",
58446 => "1111111110000100",
58447 => "1111111110000100",
58448 => "1111111110000100",
58449 => "1111111110000100",
58450 => "1111111110000100",
58451 => "1111111110000100",
58452 => "1111111110000100",
58453 => "1111111110000100",
58454 => "1111111110000100",
58455 => "1111111110000100",
58456 => "1111111110000100",
58457 => "1111111110000100",
58458 => "1111111110000100",
58459 => "1111111110000100",
58460 => "1111111110000100",
58461 => "1111111110000100",
58462 => "1111111110000100",
58463 => "1111111110000100",
58464 => "1111111110000100",
58465 => "1111111110000100",
58466 => "1111111110000100",
58467 => "1111111110000100",
58468 => "1111111110000100",
58469 => "1111111110000100",
58470 => "1111111110000100",
58471 => "1111111110000100",
58472 => "1111111110000100",
58473 => "1111111110000100",
58474 => "1111111110000100",
58475 => "1111111110000101",
58476 => "1111111110000101",
58477 => "1111111110000101",
58478 => "1111111110000101",
58479 => "1111111110000101",
58480 => "1111111110000101",
58481 => "1111111110000101",
58482 => "1111111110000101",
58483 => "1111111110000101",
58484 => "1111111110000101",
58485 => "1111111110000101",
58486 => "1111111110000101",
58487 => "1111111110000101",
58488 => "1111111110000101",
58489 => "1111111110000101",
58490 => "1111111110000101",
58491 => "1111111110000101",
58492 => "1111111110000101",
58493 => "1111111110000101",
58494 => "1111111110000101",
58495 => "1111111110000101",
58496 => "1111111110000101",
58497 => "1111111110000101",
58498 => "1111111110000101",
58499 => "1111111110000101",
58500 => "1111111110000101",
58501 => "1111111110000101",
58502 => "1111111110000101",
58503 => "1111111110000101",
58504 => "1111111110000101",
58505 => "1111111110000101",
58506 => "1111111110000101",
58507 => "1111111110000101",
58508 => "1111111110000101",
58509 => "1111111110000110",
58510 => "1111111110000110",
58511 => "1111111110000110",
58512 => "1111111110000110",
58513 => "1111111110000110",
58514 => "1111111110000110",
58515 => "1111111110000110",
58516 => "1111111110000110",
58517 => "1111111110000110",
58518 => "1111111110000110",
58519 => "1111111110000110",
58520 => "1111111110000110",
58521 => "1111111110000110",
58522 => "1111111110000110",
58523 => "1111111110000110",
58524 => "1111111110000110",
58525 => "1111111110000110",
58526 => "1111111110000110",
58527 => "1111111110000110",
58528 => "1111111110000110",
58529 => "1111111110000110",
58530 => "1111111110000110",
58531 => "1111111110000110",
58532 => "1111111110000110",
58533 => "1111111110000110",
58534 => "1111111110000110",
58535 => "1111111110000110",
58536 => "1111111110000110",
58537 => "1111111110000110",
58538 => "1111111110000110",
58539 => "1111111110000110",
58540 => "1111111110000110",
58541 => "1111111110000110",
58542 => "1111111110000110",
58543 => "1111111110000111",
58544 => "1111111110000111",
58545 => "1111111110000111",
58546 => "1111111110000111",
58547 => "1111111110000111",
58548 => "1111111110000111",
58549 => "1111111110000111",
58550 => "1111111110000111",
58551 => "1111111110000111",
58552 => "1111111110000111",
58553 => "1111111110000111",
58554 => "1111111110000111",
58555 => "1111111110000111",
58556 => "1111111110000111",
58557 => "1111111110000111",
58558 => "1111111110000111",
58559 => "1111111110000111",
58560 => "1111111110000111",
58561 => "1111111110000111",
58562 => "1111111110000111",
58563 => "1111111110000111",
58564 => "1111111110000111",
58565 => "1111111110000111",
58566 => "1111111110000111",
58567 => "1111111110000111",
58568 => "1111111110000111",
58569 => "1111111110000111",
58570 => "1111111110000111",
58571 => "1111111110000111",
58572 => "1111111110000111",
58573 => "1111111110000111",
58574 => "1111111110000111",
58575 => "1111111110000111",
58576 => "1111111110000111",
58577 => "1111111110001000",
58578 => "1111111110001000",
58579 => "1111111110001000",
58580 => "1111111110001000",
58581 => "1111111110001000",
58582 => "1111111110001000",
58583 => "1111111110001000",
58584 => "1111111110001000",
58585 => "1111111110001000",
58586 => "1111111110001000",
58587 => "1111111110001000",
58588 => "1111111110001000",
58589 => "1111111110001000",
58590 => "1111111110001000",
58591 => "1111111110001000",
58592 => "1111111110001000",
58593 => "1111111110001000",
58594 => "1111111110001000",
58595 => "1111111110001000",
58596 => "1111111110001000",
58597 => "1111111110001000",
58598 => "1111111110001000",
58599 => "1111111110001000",
58600 => "1111111110001000",
58601 => "1111111110001000",
58602 => "1111111110001000",
58603 => "1111111110001000",
58604 => "1111111110001000",
58605 => "1111111110001000",
58606 => "1111111110001000",
58607 => "1111111110001000",
58608 => "1111111110001000",
58609 => "1111111110001000",
58610 => "1111111110001000",
58611 => "1111111110001001",
58612 => "1111111110001001",
58613 => "1111111110001001",
58614 => "1111111110001001",
58615 => "1111111110001001",
58616 => "1111111110001001",
58617 => "1111111110001001",
58618 => "1111111110001001",
58619 => "1111111110001001",
58620 => "1111111110001001",
58621 => "1111111110001001",
58622 => "1111111110001001",
58623 => "1111111110001001",
58624 => "1111111110001001",
58625 => "1111111110001001",
58626 => "1111111110001001",
58627 => "1111111110001001",
58628 => "1111111110001001",
58629 => "1111111110001001",
58630 => "1111111110001001",
58631 => "1111111110001001",
58632 => "1111111110001001",
58633 => "1111111110001001",
58634 => "1111111110001001",
58635 => "1111111110001001",
58636 => "1111111110001001",
58637 => "1111111110001001",
58638 => "1111111110001001",
58639 => "1111111110001001",
58640 => "1111111110001001",
58641 => "1111111110001001",
58642 => "1111111110001001",
58643 => "1111111110001001",
58644 => "1111111110001001",
58645 => "1111111110001001",
58646 => "1111111110001010",
58647 => "1111111110001010",
58648 => "1111111110001010",
58649 => "1111111110001010",
58650 => "1111111110001010",
58651 => "1111111110001010",
58652 => "1111111110001010",
58653 => "1111111110001010",
58654 => "1111111110001010",
58655 => "1111111110001010",
58656 => "1111111110001010",
58657 => "1111111110001010",
58658 => "1111111110001010",
58659 => "1111111110001010",
58660 => "1111111110001010",
58661 => "1111111110001010",
58662 => "1111111110001010",
58663 => "1111111110001010",
58664 => "1111111110001010",
58665 => "1111111110001010",
58666 => "1111111110001010",
58667 => "1111111110001010",
58668 => "1111111110001010",
58669 => "1111111110001010",
58670 => "1111111110001010",
58671 => "1111111110001010",
58672 => "1111111110001010",
58673 => "1111111110001010",
58674 => "1111111110001010",
58675 => "1111111110001010",
58676 => "1111111110001010",
58677 => "1111111110001010",
58678 => "1111111110001010",
58679 => "1111111110001010",
58680 => "1111111110001010",
58681 => "1111111110001011",
58682 => "1111111110001011",
58683 => "1111111110001011",
58684 => "1111111110001011",
58685 => "1111111110001011",
58686 => "1111111110001011",
58687 => "1111111110001011",
58688 => "1111111110001011",
58689 => "1111111110001011",
58690 => "1111111110001011",
58691 => "1111111110001011",
58692 => "1111111110001011",
58693 => "1111111110001011",
58694 => "1111111110001011",
58695 => "1111111110001011",
58696 => "1111111110001011",
58697 => "1111111110001011",
58698 => "1111111110001011",
58699 => "1111111110001011",
58700 => "1111111110001011",
58701 => "1111111110001011",
58702 => "1111111110001011",
58703 => "1111111110001011",
58704 => "1111111110001011",
58705 => "1111111110001011",
58706 => "1111111110001011",
58707 => "1111111110001011",
58708 => "1111111110001011",
58709 => "1111111110001011",
58710 => "1111111110001011",
58711 => "1111111110001011",
58712 => "1111111110001011",
58713 => "1111111110001011",
58714 => "1111111110001011",
58715 => "1111111110001011",
58716 => "1111111110001100",
58717 => "1111111110001100",
58718 => "1111111110001100",
58719 => "1111111110001100",
58720 => "1111111110001100",
58721 => "1111111110001100",
58722 => "1111111110001100",
58723 => "1111111110001100",
58724 => "1111111110001100",
58725 => "1111111110001100",
58726 => "1111111110001100",
58727 => "1111111110001100",
58728 => "1111111110001100",
58729 => "1111111110001100",
58730 => "1111111110001100",
58731 => "1111111110001100",
58732 => "1111111110001100",
58733 => "1111111110001100",
58734 => "1111111110001100",
58735 => "1111111110001100",
58736 => "1111111110001100",
58737 => "1111111110001100",
58738 => "1111111110001100",
58739 => "1111111110001100",
58740 => "1111111110001100",
58741 => "1111111110001100",
58742 => "1111111110001100",
58743 => "1111111110001100",
58744 => "1111111110001100",
58745 => "1111111110001100",
58746 => "1111111110001100",
58747 => "1111111110001100",
58748 => "1111111110001100",
58749 => "1111111110001100",
58750 => "1111111110001100",
58751 => "1111111110001101",
58752 => "1111111110001101",
58753 => "1111111110001101",
58754 => "1111111110001101",
58755 => "1111111110001101",
58756 => "1111111110001101",
58757 => "1111111110001101",
58758 => "1111111110001101",
58759 => "1111111110001101",
58760 => "1111111110001101",
58761 => "1111111110001101",
58762 => "1111111110001101",
58763 => "1111111110001101",
58764 => "1111111110001101",
58765 => "1111111110001101",
58766 => "1111111110001101",
58767 => "1111111110001101",
58768 => "1111111110001101",
58769 => "1111111110001101",
58770 => "1111111110001101",
58771 => "1111111110001101",
58772 => "1111111110001101",
58773 => "1111111110001101",
58774 => "1111111110001101",
58775 => "1111111110001101",
58776 => "1111111110001101",
58777 => "1111111110001101",
58778 => "1111111110001101",
58779 => "1111111110001101",
58780 => "1111111110001101",
58781 => "1111111110001101",
58782 => "1111111110001101",
58783 => "1111111110001101",
58784 => "1111111110001101",
58785 => "1111111110001101",
58786 => "1111111110001101",
58787 => "1111111110001110",
58788 => "1111111110001110",
58789 => "1111111110001110",
58790 => "1111111110001110",
58791 => "1111111110001110",
58792 => "1111111110001110",
58793 => "1111111110001110",
58794 => "1111111110001110",
58795 => "1111111110001110",
58796 => "1111111110001110",
58797 => "1111111110001110",
58798 => "1111111110001110",
58799 => "1111111110001110",
58800 => "1111111110001110",
58801 => "1111111110001110",
58802 => "1111111110001110",
58803 => "1111111110001110",
58804 => "1111111110001110",
58805 => "1111111110001110",
58806 => "1111111110001110",
58807 => "1111111110001110",
58808 => "1111111110001110",
58809 => "1111111110001110",
58810 => "1111111110001110",
58811 => "1111111110001110",
58812 => "1111111110001110",
58813 => "1111111110001110",
58814 => "1111111110001110",
58815 => "1111111110001110",
58816 => "1111111110001110",
58817 => "1111111110001110",
58818 => "1111111110001110",
58819 => "1111111110001110",
58820 => "1111111110001110",
58821 => "1111111110001110",
58822 => "1111111110001110",
58823 => "1111111110001111",
58824 => "1111111110001111",
58825 => "1111111110001111",
58826 => "1111111110001111",
58827 => "1111111110001111",
58828 => "1111111110001111",
58829 => "1111111110001111",
58830 => "1111111110001111",
58831 => "1111111110001111",
58832 => "1111111110001111",
58833 => "1111111110001111",
58834 => "1111111110001111",
58835 => "1111111110001111",
58836 => "1111111110001111",
58837 => "1111111110001111",
58838 => "1111111110001111",
58839 => "1111111110001111",
58840 => "1111111110001111",
58841 => "1111111110001111",
58842 => "1111111110001111",
58843 => "1111111110001111",
58844 => "1111111110001111",
58845 => "1111111110001111",
58846 => "1111111110001111",
58847 => "1111111110001111",
58848 => "1111111110001111",
58849 => "1111111110001111",
58850 => "1111111110001111",
58851 => "1111111110001111",
58852 => "1111111110001111",
58853 => "1111111110001111",
58854 => "1111111110001111",
58855 => "1111111110001111",
58856 => "1111111110001111",
58857 => "1111111110001111",
58858 => "1111111110001111",
58859 => "1111111110001111",
58860 => "1111111110010000",
58861 => "1111111110010000",
58862 => "1111111110010000",
58863 => "1111111110010000",
58864 => "1111111110010000",
58865 => "1111111110010000",
58866 => "1111111110010000",
58867 => "1111111110010000",
58868 => "1111111110010000",
58869 => "1111111110010000",
58870 => "1111111110010000",
58871 => "1111111110010000",
58872 => "1111111110010000",
58873 => "1111111110010000",
58874 => "1111111110010000",
58875 => "1111111110010000",
58876 => "1111111110010000",
58877 => "1111111110010000",
58878 => "1111111110010000",
58879 => "1111111110010000",
58880 => "1111111110010000",
58881 => "1111111110010000",
58882 => "1111111110010000",
58883 => "1111111110010000",
58884 => "1111111110010000",
58885 => "1111111110010000",
58886 => "1111111110010000",
58887 => "1111111110010000",
58888 => "1111111110010000",
58889 => "1111111110010000",
58890 => "1111111110010000",
58891 => "1111111110010000",
58892 => "1111111110010000",
58893 => "1111111110010000",
58894 => "1111111110010000",
58895 => "1111111110010000",
58896 => "1111111110010000",
58897 => "1111111110010001",
58898 => "1111111110010001",
58899 => "1111111110010001",
58900 => "1111111110010001",
58901 => "1111111110010001",
58902 => "1111111110010001",
58903 => "1111111110010001",
58904 => "1111111110010001",
58905 => "1111111110010001",
58906 => "1111111110010001",
58907 => "1111111110010001",
58908 => "1111111110010001",
58909 => "1111111110010001",
58910 => "1111111110010001",
58911 => "1111111110010001",
58912 => "1111111110010001",
58913 => "1111111110010001",
58914 => "1111111110010001",
58915 => "1111111110010001",
58916 => "1111111110010001",
58917 => "1111111110010001",
58918 => "1111111110010001",
58919 => "1111111110010001",
58920 => "1111111110010001",
58921 => "1111111110010001",
58922 => "1111111110010001",
58923 => "1111111110010001",
58924 => "1111111110010001",
58925 => "1111111110010001",
58926 => "1111111110010001",
58927 => "1111111110010001",
58928 => "1111111110010001",
58929 => "1111111110010001",
58930 => "1111111110010001",
58931 => "1111111110010001",
58932 => "1111111110010001",
58933 => "1111111110010001",
58934 => "1111111110010010",
58935 => "1111111110010010",
58936 => "1111111110010010",
58937 => "1111111110010010",
58938 => "1111111110010010",
58939 => "1111111110010010",
58940 => "1111111110010010",
58941 => "1111111110010010",
58942 => "1111111110010010",
58943 => "1111111110010010",
58944 => "1111111110010010",
58945 => "1111111110010010",
58946 => "1111111110010010",
58947 => "1111111110010010",
58948 => "1111111110010010",
58949 => "1111111110010010",
58950 => "1111111110010010",
58951 => "1111111110010010",
58952 => "1111111110010010",
58953 => "1111111110010010",
58954 => "1111111110010010",
58955 => "1111111110010010",
58956 => "1111111110010010",
58957 => "1111111110010010",
58958 => "1111111110010010",
58959 => "1111111110010010",
58960 => "1111111110010010",
58961 => "1111111110010010",
58962 => "1111111110010010",
58963 => "1111111110010010",
58964 => "1111111110010010",
58965 => "1111111110010010",
58966 => "1111111110010010",
58967 => "1111111110010010",
58968 => "1111111110010010",
58969 => "1111111110010010",
58970 => "1111111110010010",
58971 => "1111111110010011",
58972 => "1111111110010011",
58973 => "1111111110010011",
58974 => "1111111110010011",
58975 => "1111111110010011",
58976 => "1111111110010011",
58977 => "1111111110010011",
58978 => "1111111110010011",
58979 => "1111111110010011",
58980 => "1111111110010011",
58981 => "1111111110010011",
58982 => "1111111110010011",
58983 => "1111111110010011",
58984 => "1111111110010011",
58985 => "1111111110010011",
58986 => "1111111110010011",
58987 => "1111111110010011",
58988 => "1111111110010011",
58989 => "1111111110010011",
58990 => "1111111110010011",
58991 => "1111111110010011",
58992 => "1111111110010011",
58993 => "1111111110010011",
58994 => "1111111110010011",
58995 => "1111111110010011",
58996 => "1111111110010011",
58997 => "1111111110010011",
58998 => "1111111110010011",
58999 => "1111111110010011",
59000 => "1111111110010011",
59001 => "1111111110010011",
59002 => "1111111110010011",
59003 => "1111111110010011",
59004 => "1111111110010011",
59005 => "1111111110010011",
59006 => "1111111110010011",
59007 => "1111111110010011",
59008 => "1111111110010011",
59009 => "1111111110010100",
59010 => "1111111110010100",
59011 => "1111111110010100",
59012 => "1111111110010100",
59013 => "1111111110010100",
59014 => "1111111110010100",
59015 => "1111111110010100",
59016 => "1111111110010100",
59017 => "1111111110010100",
59018 => "1111111110010100",
59019 => "1111111110010100",
59020 => "1111111110010100",
59021 => "1111111110010100",
59022 => "1111111110010100",
59023 => "1111111110010100",
59024 => "1111111110010100",
59025 => "1111111110010100",
59026 => "1111111110010100",
59027 => "1111111110010100",
59028 => "1111111110010100",
59029 => "1111111110010100",
59030 => "1111111110010100",
59031 => "1111111110010100",
59032 => "1111111110010100",
59033 => "1111111110010100",
59034 => "1111111110010100",
59035 => "1111111110010100",
59036 => "1111111110010100",
59037 => "1111111110010100",
59038 => "1111111110010100",
59039 => "1111111110010100",
59040 => "1111111110010100",
59041 => "1111111110010100",
59042 => "1111111110010100",
59043 => "1111111110010100",
59044 => "1111111110010100",
59045 => "1111111110010100",
59046 => "1111111110010100",
59047 => "1111111110010101",
59048 => "1111111110010101",
59049 => "1111111110010101",
59050 => "1111111110010101",
59051 => "1111111110010101",
59052 => "1111111110010101",
59053 => "1111111110010101",
59054 => "1111111110010101",
59055 => "1111111110010101",
59056 => "1111111110010101",
59057 => "1111111110010101",
59058 => "1111111110010101",
59059 => "1111111110010101",
59060 => "1111111110010101",
59061 => "1111111110010101",
59062 => "1111111110010101",
59063 => "1111111110010101",
59064 => "1111111110010101",
59065 => "1111111110010101",
59066 => "1111111110010101",
59067 => "1111111110010101",
59068 => "1111111110010101",
59069 => "1111111110010101",
59070 => "1111111110010101",
59071 => "1111111110010101",
59072 => "1111111110010101",
59073 => "1111111110010101",
59074 => "1111111110010101",
59075 => "1111111110010101",
59076 => "1111111110010101",
59077 => "1111111110010101",
59078 => "1111111110010101",
59079 => "1111111110010101",
59080 => "1111111110010101",
59081 => "1111111110010101",
59082 => "1111111110010101",
59083 => "1111111110010101",
59084 => "1111111110010101",
59085 => "1111111110010101",
59086 => "1111111110010110",
59087 => "1111111110010110",
59088 => "1111111110010110",
59089 => "1111111110010110",
59090 => "1111111110010110",
59091 => "1111111110010110",
59092 => "1111111110010110",
59093 => "1111111110010110",
59094 => "1111111110010110",
59095 => "1111111110010110",
59096 => "1111111110010110",
59097 => "1111111110010110",
59098 => "1111111110010110",
59099 => "1111111110010110",
59100 => "1111111110010110",
59101 => "1111111110010110",
59102 => "1111111110010110",
59103 => "1111111110010110",
59104 => "1111111110010110",
59105 => "1111111110010110",
59106 => "1111111110010110",
59107 => "1111111110010110",
59108 => "1111111110010110",
59109 => "1111111110010110",
59110 => "1111111110010110",
59111 => "1111111110010110",
59112 => "1111111110010110",
59113 => "1111111110010110",
59114 => "1111111110010110",
59115 => "1111111110010110",
59116 => "1111111110010110",
59117 => "1111111110010110",
59118 => "1111111110010110",
59119 => "1111111110010110",
59120 => "1111111110010110",
59121 => "1111111110010110",
59122 => "1111111110010110",
59123 => "1111111110010110",
59124 => "1111111110010110",
59125 => "1111111110010111",
59126 => "1111111110010111",
59127 => "1111111110010111",
59128 => "1111111110010111",
59129 => "1111111110010111",
59130 => "1111111110010111",
59131 => "1111111110010111",
59132 => "1111111110010111",
59133 => "1111111110010111",
59134 => "1111111110010111",
59135 => "1111111110010111",
59136 => "1111111110010111",
59137 => "1111111110010111",
59138 => "1111111110010111",
59139 => "1111111110010111",
59140 => "1111111110010111",
59141 => "1111111110010111",
59142 => "1111111110010111",
59143 => "1111111110010111",
59144 => "1111111110010111",
59145 => "1111111110010111",
59146 => "1111111110010111",
59147 => "1111111110010111",
59148 => "1111111110010111",
59149 => "1111111110010111",
59150 => "1111111110010111",
59151 => "1111111110010111",
59152 => "1111111110010111",
59153 => "1111111110010111",
59154 => "1111111110010111",
59155 => "1111111110010111",
59156 => "1111111110010111",
59157 => "1111111110010111",
59158 => "1111111110010111",
59159 => "1111111110010111",
59160 => "1111111110010111",
59161 => "1111111110010111",
59162 => "1111111110010111",
59163 => "1111111110010111",
59164 => "1111111110011000",
59165 => "1111111110011000",
59166 => "1111111110011000",
59167 => "1111111110011000",
59168 => "1111111110011000",
59169 => "1111111110011000",
59170 => "1111111110011000",
59171 => "1111111110011000",
59172 => "1111111110011000",
59173 => "1111111110011000",
59174 => "1111111110011000",
59175 => "1111111110011000",
59176 => "1111111110011000",
59177 => "1111111110011000",
59178 => "1111111110011000",
59179 => "1111111110011000",
59180 => "1111111110011000",
59181 => "1111111110011000",
59182 => "1111111110011000",
59183 => "1111111110011000",
59184 => "1111111110011000",
59185 => "1111111110011000",
59186 => "1111111110011000",
59187 => "1111111110011000",
59188 => "1111111110011000",
59189 => "1111111110011000",
59190 => "1111111110011000",
59191 => "1111111110011000",
59192 => "1111111110011000",
59193 => "1111111110011000",
59194 => "1111111110011000",
59195 => "1111111110011000",
59196 => "1111111110011000",
59197 => "1111111110011000",
59198 => "1111111110011000",
59199 => "1111111110011000",
59200 => "1111111110011000",
59201 => "1111111110011000",
59202 => "1111111110011000",
59203 => "1111111110011001",
59204 => "1111111110011001",
59205 => "1111111110011001",
59206 => "1111111110011001",
59207 => "1111111110011001",
59208 => "1111111110011001",
59209 => "1111111110011001",
59210 => "1111111110011001",
59211 => "1111111110011001",
59212 => "1111111110011001",
59213 => "1111111110011001",
59214 => "1111111110011001",
59215 => "1111111110011001",
59216 => "1111111110011001",
59217 => "1111111110011001",
59218 => "1111111110011001",
59219 => "1111111110011001",
59220 => "1111111110011001",
59221 => "1111111110011001",
59222 => "1111111110011001",
59223 => "1111111110011001",
59224 => "1111111110011001",
59225 => "1111111110011001",
59226 => "1111111110011001",
59227 => "1111111110011001",
59228 => "1111111110011001",
59229 => "1111111110011001",
59230 => "1111111110011001",
59231 => "1111111110011001",
59232 => "1111111110011001",
59233 => "1111111110011001",
59234 => "1111111110011001",
59235 => "1111111110011001",
59236 => "1111111110011001",
59237 => "1111111110011001",
59238 => "1111111110011001",
59239 => "1111111110011001",
59240 => "1111111110011001",
59241 => "1111111110011001",
59242 => "1111111110011001",
59243 => "1111111110011010",
59244 => "1111111110011010",
59245 => "1111111110011010",
59246 => "1111111110011010",
59247 => "1111111110011010",
59248 => "1111111110011010",
59249 => "1111111110011010",
59250 => "1111111110011010",
59251 => "1111111110011010",
59252 => "1111111110011010",
59253 => "1111111110011010",
59254 => "1111111110011010",
59255 => "1111111110011010",
59256 => "1111111110011010",
59257 => "1111111110011010",
59258 => "1111111110011010",
59259 => "1111111110011010",
59260 => "1111111110011010",
59261 => "1111111110011010",
59262 => "1111111110011010",
59263 => "1111111110011010",
59264 => "1111111110011010",
59265 => "1111111110011010",
59266 => "1111111110011010",
59267 => "1111111110011010",
59268 => "1111111110011010",
59269 => "1111111110011010",
59270 => "1111111110011010",
59271 => "1111111110011010",
59272 => "1111111110011010",
59273 => "1111111110011010",
59274 => "1111111110011010",
59275 => "1111111110011010",
59276 => "1111111110011010",
59277 => "1111111110011010",
59278 => "1111111110011010",
59279 => "1111111110011010",
59280 => "1111111110011010",
59281 => "1111111110011010",
59282 => "1111111110011010",
59283 => "1111111110011010",
59284 => "1111111110011011",
59285 => "1111111110011011",
59286 => "1111111110011011",
59287 => "1111111110011011",
59288 => "1111111110011011",
59289 => "1111111110011011",
59290 => "1111111110011011",
59291 => "1111111110011011",
59292 => "1111111110011011",
59293 => "1111111110011011",
59294 => "1111111110011011",
59295 => "1111111110011011",
59296 => "1111111110011011",
59297 => "1111111110011011",
59298 => "1111111110011011",
59299 => "1111111110011011",
59300 => "1111111110011011",
59301 => "1111111110011011",
59302 => "1111111110011011",
59303 => "1111111110011011",
59304 => "1111111110011011",
59305 => "1111111110011011",
59306 => "1111111110011011",
59307 => "1111111110011011",
59308 => "1111111110011011",
59309 => "1111111110011011",
59310 => "1111111110011011",
59311 => "1111111110011011",
59312 => "1111111110011011",
59313 => "1111111110011011",
59314 => "1111111110011011",
59315 => "1111111110011011",
59316 => "1111111110011011",
59317 => "1111111110011011",
59318 => "1111111110011011",
59319 => "1111111110011011",
59320 => "1111111110011011",
59321 => "1111111110011011",
59322 => "1111111110011011",
59323 => "1111111110011011",
59324 => "1111111110011011",
59325 => "1111111110011100",
59326 => "1111111110011100",
59327 => "1111111110011100",
59328 => "1111111110011100",
59329 => "1111111110011100",
59330 => "1111111110011100",
59331 => "1111111110011100",
59332 => "1111111110011100",
59333 => "1111111110011100",
59334 => "1111111110011100",
59335 => "1111111110011100",
59336 => "1111111110011100",
59337 => "1111111110011100",
59338 => "1111111110011100",
59339 => "1111111110011100",
59340 => "1111111110011100",
59341 => "1111111110011100",
59342 => "1111111110011100",
59343 => "1111111110011100",
59344 => "1111111110011100",
59345 => "1111111110011100",
59346 => "1111111110011100",
59347 => "1111111110011100",
59348 => "1111111110011100",
59349 => "1111111110011100",
59350 => "1111111110011100",
59351 => "1111111110011100",
59352 => "1111111110011100",
59353 => "1111111110011100",
59354 => "1111111110011100",
59355 => "1111111110011100",
59356 => "1111111110011100",
59357 => "1111111110011100",
59358 => "1111111110011100",
59359 => "1111111110011100",
59360 => "1111111110011100",
59361 => "1111111110011100",
59362 => "1111111110011100",
59363 => "1111111110011100",
59364 => "1111111110011100",
59365 => "1111111110011100",
59366 => "1111111110011101",
59367 => "1111111110011101",
59368 => "1111111110011101",
59369 => "1111111110011101",
59370 => "1111111110011101",
59371 => "1111111110011101",
59372 => "1111111110011101",
59373 => "1111111110011101",
59374 => "1111111110011101",
59375 => "1111111110011101",
59376 => "1111111110011101",
59377 => "1111111110011101",
59378 => "1111111110011101",
59379 => "1111111110011101",
59380 => "1111111110011101",
59381 => "1111111110011101",
59382 => "1111111110011101",
59383 => "1111111110011101",
59384 => "1111111110011101",
59385 => "1111111110011101",
59386 => "1111111110011101",
59387 => "1111111110011101",
59388 => "1111111110011101",
59389 => "1111111110011101",
59390 => "1111111110011101",
59391 => "1111111110011101",
59392 => "1111111110011101",
59393 => "1111111110011101",
59394 => "1111111110011101",
59395 => "1111111110011101",
59396 => "1111111110011101",
59397 => "1111111110011101",
59398 => "1111111110011101",
59399 => "1111111110011101",
59400 => "1111111110011101",
59401 => "1111111110011101",
59402 => "1111111110011101",
59403 => "1111111110011101",
59404 => "1111111110011101",
59405 => "1111111110011101",
59406 => "1111111110011101",
59407 => "1111111110011101",
59408 => "1111111110011110",
59409 => "1111111110011110",
59410 => "1111111110011110",
59411 => "1111111110011110",
59412 => "1111111110011110",
59413 => "1111111110011110",
59414 => "1111111110011110",
59415 => "1111111110011110",
59416 => "1111111110011110",
59417 => "1111111110011110",
59418 => "1111111110011110",
59419 => "1111111110011110",
59420 => "1111111110011110",
59421 => "1111111110011110",
59422 => "1111111110011110",
59423 => "1111111110011110",
59424 => "1111111110011110",
59425 => "1111111110011110",
59426 => "1111111110011110",
59427 => "1111111110011110",
59428 => "1111111110011110",
59429 => "1111111110011110",
59430 => "1111111110011110",
59431 => "1111111110011110",
59432 => "1111111110011110",
59433 => "1111111110011110",
59434 => "1111111110011110",
59435 => "1111111110011110",
59436 => "1111111110011110",
59437 => "1111111110011110",
59438 => "1111111110011110",
59439 => "1111111110011110",
59440 => "1111111110011110",
59441 => "1111111110011110",
59442 => "1111111110011110",
59443 => "1111111110011110",
59444 => "1111111110011110",
59445 => "1111111110011110",
59446 => "1111111110011110",
59447 => "1111111110011110",
59448 => "1111111110011110",
59449 => "1111111110011110",
59450 => "1111111110011111",
59451 => "1111111110011111",
59452 => "1111111110011111",
59453 => "1111111110011111",
59454 => "1111111110011111",
59455 => "1111111110011111",
59456 => "1111111110011111",
59457 => "1111111110011111",
59458 => "1111111110011111",
59459 => "1111111110011111",
59460 => "1111111110011111",
59461 => "1111111110011111",
59462 => "1111111110011111",
59463 => "1111111110011111",
59464 => "1111111110011111",
59465 => "1111111110011111",
59466 => "1111111110011111",
59467 => "1111111110011111",
59468 => "1111111110011111",
59469 => "1111111110011111",
59470 => "1111111110011111",
59471 => "1111111110011111",
59472 => "1111111110011111",
59473 => "1111111110011111",
59474 => "1111111110011111",
59475 => "1111111110011111",
59476 => "1111111110011111",
59477 => "1111111110011111",
59478 => "1111111110011111",
59479 => "1111111110011111",
59480 => "1111111110011111",
59481 => "1111111110011111",
59482 => "1111111110011111",
59483 => "1111111110011111",
59484 => "1111111110011111",
59485 => "1111111110011111",
59486 => "1111111110011111",
59487 => "1111111110011111",
59488 => "1111111110011111",
59489 => "1111111110011111",
59490 => "1111111110011111",
59491 => "1111111110011111",
59492 => "1111111110100000",
59493 => "1111111110100000",
59494 => "1111111110100000",
59495 => "1111111110100000",
59496 => "1111111110100000",
59497 => "1111111110100000",
59498 => "1111111110100000",
59499 => "1111111110100000",
59500 => "1111111110100000",
59501 => "1111111110100000",
59502 => "1111111110100000",
59503 => "1111111110100000",
59504 => "1111111110100000",
59505 => "1111111110100000",
59506 => "1111111110100000",
59507 => "1111111110100000",
59508 => "1111111110100000",
59509 => "1111111110100000",
59510 => "1111111110100000",
59511 => "1111111110100000",
59512 => "1111111110100000",
59513 => "1111111110100000",
59514 => "1111111110100000",
59515 => "1111111110100000",
59516 => "1111111110100000",
59517 => "1111111110100000",
59518 => "1111111110100000",
59519 => "1111111110100000",
59520 => "1111111110100000",
59521 => "1111111110100000",
59522 => "1111111110100000",
59523 => "1111111110100000",
59524 => "1111111110100000",
59525 => "1111111110100000",
59526 => "1111111110100000",
59527 => "1111111110100000",
59528 => "1111111110100000",
59529 => "1111111110100000",
59530 => "1111111110100000",
59531 => "1111111110100000",
59532 => "1111111110100000",
59533 => "1111111110100000",
59534 => "1111111110100000",
59535 => "1111111110100001",
59536 => "1111111110100001",
59537 => "1111111110100001",
59538 => "1111111110100001",
59539 => "1111111110100001",
59540 => "1111111110100001",
59541 => "1111111110100001",
59542 => "1111111110100001",
59543 => "1111111110100001",
59544 => "1111111110100001",
59545 => "1111111110100001",
59546 => "1111111110100001",
59547 => "1111111110100001",
59548 => "1111111110100001",
59549 => "1111111110100001",
59550 => "1111111110100001",
59551 => "1111111110100001",
59552 => "1111111110100001",
59553 => "1111111110100001",
59554 => "1111111110100001",
59555 => "1111111110100001",
59556 => "1111111110100001",
59557 => "1111111110100001",
59558 => "1111111110100001",
59559 => "1111111110100001",
59560 => "1111111110100001",
59561 => "1111111110100001",
59562 => "1111111110100001",
59563 => "1111111110100001",
59564 => "1111111110100001",
59565 => "1111111110100001",
59566 => "1111111110100001",
59567 => "1111111110100001",
59568 => "1111111110100001",
59569 => "1111111110100001",
59570 => "1111111110100001",
59571 => "1111111110100001",
59572 => "1111111110100001",
59573 => "1111111110100001",
59574 => "1111111110100001",
59575 => "1111111110100001",
59576 => "1111111110100001",
59577 => "1111111110100001",
59578 => "1111111110100010",
59579 => "1111111110100010",
59580 => "1111111110100010",
59581 => "1111111110100010",
59582 => "1111111110100010",
59583 => "1111111110100010",
59584 => "1111111110100010",
59585 => "1111111110100010",
59586 => "1111111110100010",
59587 => "1111111110100010",
59588 => "1111111110100010",
59589 => "1111111110100010",
59590 => "1111111110100010",
59591 => "1111111110100010",
59592 => "1111111110100010",
59593 => "1111111110100010",
59594 => "1111111110100010",
59595 => "1111111110100010",
59596 => "1111111110100010",
59597 => "1111111110100010",
59598 => "1111111110100010",
59599 => "1111111110100010",
59600 => "1111111110100010",
59601 => "1111111110100010",
59602 => "1111111110100010",
59603 => "1111111110100010",
59604 => "1111111110100010",
59605 => "1111111110100010",
59606 => "1111111110100010",
59607 => "1111111110100010",
59608 => "1111111110100010",
59609 => "1111111110100010",
59610 => "1111111110100010",
59611 => "1111111110100010",
59612 => "1111111110100010",
59613 => "1111111110100010",
59614 => "1111111110100010",
59615 => "1111111110100010",
59616 => "1111111110100010",
59617 => "1111111110100010",
59618 => "1111111110100010",
59619 => "1111111110100010",
59620 => "1111111110100010",
59621 => "1111111110100010",
59622 => "1111111110100011",
59623 => "1111111110100011",
59624 => "1111111110100011",
59625 => "1111111110100011",
59626 => "1111111110100011",
59627 => "1111111110100011",
59628 => "1111111110100011",
59629 => "1111111110100011",
59630 => "1111111110100011",
59631 => "1111111110100011",
59632 => "1111111110100011",
59633 => "1111111110100011",
59634 => "1111111110100011",
59635 => "1111111110100011",
59636 => "1111111110100011",
59637 => "1111111110100011",
59638 => "1111111110100011",
59639 => "1111111110100011",
59640 => "1111111110100011",
59641 => "1111111110100011",
59642 => "1111111110100011",
59643 => "1111111110100011",
59644 => "1111111110100011",
59645 => "1111111110100011",
59646 => "1111111110100011",
59647 => "1111111110100011",
59648 => "1111111110100011",
59649 => "1111111110100011",
59650 => "1111111110100011",
59651 => "1111111110100011",
59652 => "1111111110100011",
59653 => "1111111110100011",
59654 => "1111111110100011",
59655 => "1111111110100011",
59656 => "1111111110100011",
59657 => "1111111110100011",
59658 => "1111111110100011",
59659 => "1111111110100011",
59660 => "1111111110100011",
59661 => "1111111110100011",
59662 => "1111111110100011",
59663 => "1111111110100011",
59664 => "1111111110100011",
59665 => "1111111110100011",
59666 => "1111111110100011",
59667 => "1111111110100100",
59668 => "1111111110100100",
59669 => "1111111110100100",
59670 => "1111111110100100",
59671 => "1111111110100100",
59672 => "1111111110100100",
59673 => "1111111110100100",
59674 => "1111111110100100",
59675 => "1111111110100100",
59676 => "1111111110100100",
59677 => "1111111110100100",
59678 => "1111111110100100",
59679 => "1111111110100100",
59680 => "1111111110100100",
59681 => "1111111110100100",
59682 => "1111111110100100",
59683 => "1111111110100100",
59684 => "1111111110100100",
59685 => "1111111110100100",
59686 => "1111111110100100",
59687 => "1111111110100100",
59688 => "1111111110100100",
59689 => "1111111110100100",
59690 => "1111111110100100",
59691 => "1111111110100100",
59692 => "1111111110100100",
59693 => "1111111110100100",
59694 => "1111111110100100",
59695 => "1111111110100100",
59696 => "1111111110100100",
59697 => "1111111110100100",
59698 => "1111111110100100",
59699 => "1111111110100100",
59700 => "1111111110100100",
59701 => "1111111110100100",
59702 => "1111111110100100",
59703 => "1111111110100100",
59704 => "1111111110100100",
59705 => "1111111110100100",
59706 => "1111111110100100",
59707 => "1111111110100100",
59708 => "1111111110100100",
59709 => "1111111110100100",
59710 => "1111111110100100",
59711 => "1111111110100100",
59712 => "1111111110100101",
59713 => "1111111110100101",
59714 => "1111111110100101",
59715 => "1111111110100101",
59716 => "1111111110100101",
59717 => "1111111110100101",
59718 => "1111111110100101",
59719 => "1111111110100101",
59720 => "1111111110100101",
59721 => "1111111110100101",
59722 => "1111111110100101",
59723 => "1111111110100101",
59724 => "1111111110100101",
59725 => "1111111110100101",
59726 => "1111111110100101",
59727 => "1111111110100101",
59728 => "1111111110100101",
59729 => "1111111110100101",
59730 => "1111111110100101",
59731 => "1111111110100101",
59732 => "1111111110100101",
59733 => "1111111110100101",
59734 => "1111111110100101",
59735 => "1111111110100101",
59736 => "1111111110100101",
59737 => "1111111110100101",
59738 => "1111111110100101",
59739 => "1111111110100101",
59740 => "1111111110100101",
59741 => "1111111110100101",
59742 => "1111111110100101",
59743 => "1111111110100101",
59744 => "1111111110100101",
59745 => "1111111110100101",
59746 => "1111111110100101",
59747 => "1111111110100101",
59748 => "1111111110100101",
59749 => "1111111110100101",
59750 => "1111111110100101",
59751 => "1111111110100101",
59752 => "1111111110100101",
59753 => "1111111110100101",
59754 => "1111111110100101",
59755 => "1111111110100101",
59756 => "1111111110100101",
59757 => "1111111110100110",
59758 => "1111111110100110",
59759 => "1111111110100110",
59760 => "1111111110100110",
59761 => "1111111110100110",
59762 => "1111111110100110",
59763 => "1111111110100110",
59764 => "1111111110100110",
59765 => "1111111110100110",
59766 => "1111111110100110",
59767 => "1111111110100110",
59768 => "1111111110100110",
59769 => "1111111110100110",
59770 => "1111111110100110",
59771 => "1111111110100110",
59772 => "1111111110100110",
59773 => "1111111110100110",
59774 => "1111111110100110",
59775 => "1111111110100110",
59776 => "1111111110100110",
59777 => "1111111110100110",
59778 => "1111111110100110",
59779 => "1111111110100110",
59780 => "1111111110100110",
59781 => "1111111110100110",
59782 => "1111111110100110",
59783 => "1111111110100110",
59784 => "1111111110100110",
59785 => "1111111110100110",
59786 => "1111111110100110",
59787 => "1111111110100110",
59788 => "1111111110100110",
59789 => "1111111110100110",
59790 => "1111111110100110",
59791 => "1111111110100110",
59792 => "1111111110100110",
59793 => "1111111110100110",
59794 => "1111111110100110",
59795 => "1111111110100110",
59796 => "1111111110100110",
59797 => "1111111110100110",
59798 => "1111111110100110",
59799 => "1111111110100110",
59800 => "1111111110100110",
59801 => "1111111110100110",
59802 => "1111111110100110",
59803 => "1111111110100111",
59804 => "1111111110100111",
59805 => "1111111110100111",
59806 => "1111111110100111",
59807 => "1111111110100111",
59808 => "1111111110100111",
59809 => "1111111110100111",
59810 => "1111111110100111",
59811 => "1111111110100111",
59812 => "1111111110100111",
59813 => "1111111110100111",
59814 => "1111111110100111",
59815 => "1111111110100111",
59816 => "1111111110100111",
59817 => "1111111110100111",
59818 => "1111111110100111",
59819 => "1111111110100111",
59820 => "1111111110100111",
59821 => "1111111110100111",
59822 => "1111111110100111",
59823 => "1111111110100111",
59824 => "1111111110100111",
59825 => "1111111110100111",
59826 => "1111111110100111",
59827 => "1111111110100111",
59828 => "1111111110100111",
59829 => "1111111110100111",
59830 => "1111111110100111",
59831 => "1111111110100111",
59832 => "1111111110100111",
59833 => "1111111110100111",
59834 => "1111111110100111",
59835 => "1111111110100111",
59836 => "1111111110100111",
59837 => "1111111110100111",
59838 => "1111111110100111",
59839 => "1111111110100111",
59840 => "1111111110100111",
59841 => "1111111110100111",
59842 => "1111111110100111",
59843 => "1111111110100111",
59844 => "1111111110100111",
59845 => "1111111110100111",
59846 => "1111111110100111",
59847 => "1111111110100111",
59848 => "1111111110100111",
59849 => "1111111110101000",
59850 => "1111111110101000",
59851 => "1111111110101000",
59852 => "1111111110101000",
59853 => "1111111110101000",
59854 => "1111111110101000",
59855 => "1111111110101000",
59856 => "1111111110101000",
59857 => "1111111110101000",
59858 => "1111111110101000",
59859 => "1111111110101000",
59860 => "1111111110101000",
59861 => "1111111110101000",
59862 => "1111111110101000",
59863 => "1111111110101000",
59864 => "1111111110101000",
59865 => "1111111110101000",
59866 => "1111111110101000",
59867 => "1111111110101000",
59868 => "1111111110101000",
59869 => "1111111110101000",
59870 => "1111111110101000",
59871 => "1111111110101000",
59872 => "1111111110101000",
59873 => "1111111110101000",
59874 => "1111111110101000",
59875 => "1111111110101000",
59876 => "1111111110101000",
59877 => "1111111110101000",
59878 => "1111111110101000",
59879 => "1111111110101000",
59880 => "1111111110101000",
59881 => "1111111110101000",
59882 => "1111111110101000",
59883 => "1111111110101000",
59884 => "1111111110101000",
59885 => "1111111110101000",
59886 => "1111111110101000",
59887 => "1111111110101000",
59888 => "1111111110101000",
59889 => "1111111110101000",
59890 => "1111111110101000",
59891 => "1111111110101000",
59892 => "1111111110101000",
59893 => "1111111110101000",
59894 => "1111111110101000",
59895 => "1111111110101000",
59896 => "1111111110101001",
59897 => "1111111110101001",
59898 => "1111111110101001",
59899 => "1111111110101001",
59900 => "1111111110101001",
59901 => "1111111110101001",
59902 => "1111111110101001",
59903 => "1111111110101001",
59904 => "1111111110101001",
59905 => "1111111110101001",
59906 => "1111111110101001",
59907 => "1111111110101001",
59908 => "1111111110101001",
59909 => "1111111110101001",
59910 => "1111111110101001",
59911 => "1111111110101001",
59912 => "1111111110101001",
59913 => "1111111110101001",
59914 => "1111111110101001",
59915 => "1111111110101001",
59916 => "1111111110101001",
59917 => "1111111110101001",
59918 => "1111111110101001",
59919 => "1111111110101001",
59920 => "1111111110101001",
59921 => "1111111110101001",
59922 => "1111111110101001",
59923 => "1111111110101001",
59924 => "1111111110101001",
59925 => "1111111110101001",
59926 => "1111111110101001",
59927 => "1111111110101001",
59928 => "1111111110101001",
59929 => "1111111110101001",
59930 => "1111111110101001",
59931 => "1111111110101001",
59932 => "1111111110101001",
59933 => "1111111110101001",
59934 => "1111111110101001",
59935 => "1111111110101001",
59936 => "1111111110101001",
59937 => "1111111110101001",
59938 => "1111111110101001",
59939 => "1111111110101001",
59940 => "1111111110101001",
59941 => "1111111110101001",
59942 => "1111111110101001",
59943 => "1111111110101010",
59944 => "1111111110101010",
59945 => "1111111110101010",
59946 => "1111111110101010",
59947 => "1111111110101010",
59948 => "1111111110101010",
59949 => "1111111110101010",
59950 => "1111111110101010",
59951 => "1111111110101010",
59952 => "1111111110101010",
59953 => "1111111110101010",
59954 => "1111111110101010",
59955 => "1111111110101010",
59956 => "1111111110101010",
59957 => "1111111110101010",
59958 => "1111111110101010",
59959 => "1111111110101010",
59960 => "1111111110101010",
59961 => "1111111110101010",
59962 => "1111111110101010",
59963 => "1111111110101010",
59964 => "1111111110101010",
59965 => "1111111110101010",
59966 => "1111111110101010",
59967 => "1111111110101010",
59968 => "1111111110101010",
59969 => "1111111110101010",
59970 => "1111111110101010",
59971 => "1111111110101010",
59972 => "1111111110101010",
59973 => "1111111110101010",
59974 => "1111111110101010",
59975 => "1111111110101010",
59976 => "1111111110101010",
59977 => "1111111110101010",
59978 => "1111111110101010",
59979 => "1111111110101010",
59980 => "1111111110101010",
59981 => "1111111110101010",
59982 => "1111111110101010",
59983 => "1111111110101010",
59984 => "1111111110101010",
59985 => "1111111110101010",
59986 => "1111111110101010",
59987 => "1111111110101010",
59988 => "1111111110101010",
59989 => "1111111110101010",
59990 => "1111111110101010",
59991 => "1111111110101011",
59992 => "1111111110101011",
59993 => "1111111110101011",
59994 => "1111111110101011",
59995 => "1111111110101011",
59996 => "1111111110101011",
59997 => "1111111110101011",
59998 => "1111111110101011",
59999 => "1111111110101011",
60000 => "1111111110101011",
60001 => "1111111110101011",
60002 => "1111111110101011",
60003 => "1111111110101011",
60004 => "1111111110101011",
60005 => "1111111110101011",
60006 => "1111111110101011",
60007 => "1111111110101011",
60008 => "1111111110101011",
60009 => "1111111110101011",
60010 => "1111111110101011",
60011 => "1111111110101011",
60012 => "1111111110101011",
60013 => "1111111110101011",
60014 => "1111111110101011",
60015 => "1111111110101011",
60016 => "1111111110101011",
60017 => "1111111110101011",
60018 => "1111111110101011",
60019 => "1111111110101011",
60020 => "1111111110101011",
60021 => "1111111110101011",
60022 => "1111111110101011",
60023 => "1111111110101011",
60024 => "1111111110101011",
60025 => "1111111110101011",
60026 => "1111111110101011",
60027 => "1111111110101011",
60028 => "1111111110101011",
60029 => "1111111110101011",
60030 => "1111111110101011",
60031 => "1111111110101011",
60032 => "1111111110101011",
60033 => "1111111110101011",
60034 => "1111111110101011",
60035 => "1111111110101011",
60036 => "1111111110101011",
60037 => "1111111110101011",
60038 => "1111111110101011",
60039 => "1111111110101011",
60040 => "1111111110101100",
60041 => "1111111110101100",
60042 => "1111111110101100",
60043 => "1111111110101100",
60044 => "1111111110101100",
60045 => "1111111110101100",
60046 => "1111111110101100",
60047 => "1111111110101100",
60048 => "1111111110101100",
60049 => "1111111110101100",
60050 => "1111111110101100",
60051 => "1111111110101100",
60052 => "1111111110101100",
60053 => "1111111110101100",
60054 => "1111111110101100",
60055 => "1111111110101100",
60056 => "1111111110101100",
60057 => "1111111110101100",
60058 => "1111111110101100",
60059 => "1111111110101100",
60060 => "1111111110101100",
60061 => "1111111110101100",
60062 => "1111111110101100",
60063 => "1111111110101100",
60064 => "1111111110101100",
60065 => "1111111110101100",
60066 => "1111111110101100",
60067 => "1111111110101100",
60068 => "1111111110101100",
60069 => "1111111110101100",
60070 => "1111111110101100",
60071 => "1111111110101100",
60072 => "1111111110101100",
60073 => "1111111110101100",
60074 => "1111111110101100",
60075 => "1111111110101100",
60076 => "1111111110101100",
60077 => "1111111110101100",
60078 => "1111111110101100",
60079 => "1111111110101100",
60080 => "1111111110101100",
60081 => "1111111110101100",
60082 => "1111111110101100",
60083 => "1111111110101100",
60084 => "1111111110101100",
60085 => "1111111110101100",
60086 => "1111111110101100",
60087 => "1111111110101100",
60088 => "1111111110101100",
60089 => "1111111110101101",
60090 => "1111111110101101",
60091 => "1111111110101101",
60092 => "1111111110101101",
60093 => "1111111110101101",
60094 => "1111111110101101",
60095 => "1111111110101101",
60096 => "1111111110101101",
60097 => "1111111110101101",
60098 => "1111111110101101",
60099 => "1111111110101101",
60100 => "1111111110101101",
60101 => "1111111110101101",
60102 => "1111111110101101",
60103 => "1111111110101101",
60104 => "1111111110101101",
60105 => "1111111110101101",
60106 => "1111111110101101",
60107 => "1111111110101101",
60108 => "1111111110101101",
60109 => "1111111110101101",
60110 => "1111111110101101",
60111 => "1111111110101101",
60112 => "1111111110101101",
60113 => "1111111110101101",
60114 => "1111111110101101",
60115 => "1111111110101101",
60116 => "1111111110101101",
60117 => "1111111110101101",
60118 => "1111111110101101",
60119 => "1111111110101101",
60120 => "1111111110101101",
60121 => "1111111110101101",
60122 => "1111111110101101",
60123 => "1111111110101101",
60124 => "1111111110101101",
60125 => "1111111110101101",
60126 => "1111111110101101",
60127 => "1111111110101101",
60128 => "1111111110101101",
60129 => "1111111110101101",
60130 => "1111111110101101",
60131 => "1111111110101101",
60132 => "1111111110101101",
60133 => "1111111110101101",
60134 => "1111111110101101",
60135 => "1111111110101101",
60136 => "1111111110101101",
60137 => "1111111110101101",
60138 => "1111111110101101",
60139 => "1111111110101110",
60140 => "1111111110101110",
60141 => "1111111110101110",
60142 => "1111111110101110",
60143 => "1111111110101110",
60144 => "1111111110101110",
60145 => "1111111110101110",
60146 => "1111111110101110",
60147 => "1111111110101110",
60148 => "1111111110101110",
60149 => "1111111110101110",
60150 => "1111111110101110",
60151 => "1111111110101110",
60152 => "1111111110101110",
60153 => "1111111110101110",
60154 => "1111111110101110",
60155 => "1111111110101110",
60156 => "1111111110101110",
60157 => "1111111110101110",
60158 => "1111111110101110",
60159 => "1111111110101110",
60160 => "1111111110101110",
60161 => "1111111110101110",
60162 => "1111111110101110",
60163 => "1111111110101110",
60164 => "1111111110101110",
60165 => "1111111110101110",
60166 => "1111111110101110",
60167 => "1111111110101110",
60168 => "1111111110101110",
60169 => "1111111110101110",
60170 => "1111111110101110",
60171 => "1111111110101110",
60172 => "1111111110101110",
60173 => "1111111110101110",
60174 => "1111111110101110",
60175 => "1111111110101110",
60176 => "1111111110101110",
60177 => "1111111110101110",
60178 => "1111111110101110",
60179 => "1111111110101110",
60180 => "1111111110101110",
60181 => "1111111110101110",
60182 => "1111111110101110",
60183 => "1111111110101110",
60184 => "1111111110101110",
60185 => "1111111110101110",
60186 => "1111111110101110",
60187 => "1111111110101110",
60188 => "1111111110101110",
60189 => "1111111110101111",
60190 => "1111111110101111",
60191 => "1111111110101111",
60192 => "1111111110101111",
60193 => "1111111110101111",
60194 => "1111111110101111",
60195 => "1111111110101111",
60196 => "1111111110101111",
60197 => "1111111110101111",
60198 => "1111111110101111",
60199 => "1111111110101111",
60200 => "1111111110101111",
60201 => "1111111110101111",
60202 => "1111111110101111",
60203 => "1111111110101111",
60204 => "1111111110101111",
60205 => "1111111110101111",
60206 => "1111111110101111",
60207 => "1111111110101111",
60208 => "1111111110101111",
60209 => "1111111110101111",
60210 => "1111111110101111",
60211 => "1111111110101111",
60212 => "1111111110101111",
60213 => "1111111110101111",
60214 => "1111111110101111",
60215 => "1111111110101111",
60216 => "1111111110101111",
60217 => "1111111110101111",
60218 => "1111111110101111",
60219 => "1111111110101111",
60220 => "1111111110101111",
60221 => "1111111110101111",
60222 => "1111111110101111",
60223 => "1111111110101111",
60224 => "1111111110101111",
60225 => "1111111110101111",
60226 => "1111111110101111",
60227 => "1111111110101111",
60228 => "1111111110101111",
60229 => "1111111110101111",
60230 => "1111111110101111",
60231 => "1111111110101111",
60232 => "1111111110101111",
60233 => "1111111110101111",
60234 => "1111111110101111",
60235 => "1111111110101111",
60236 => "1111111110101111",
60237 => "1111111110101111",
60238 => "1111111110101111",
60239 => "1111111110101111",
60240 => "1111111110110000",
60241 => "1111111110110000",
60242 => "1111111110110000",
60243 => "1111111110110000",
60244 => "1111111110110000",
60245 => "1111111110110000",
60246 => "1111111110110000",
60247 => "1111111110110000",
60248 => "1111111110110000",
60249 => "1111111110110000",
60250 => "1111111110110000",
60251 => "1111111110110000",
60252 => "1111111110110000",
60253 => "1111111110110000",
60254 => "1111111110110000",
60255 => "1111111110110000",
60256 => "1111111110110000",
60257 => "1111111110110000",
60258 => "1111111110110000",
60259 => "1111111110110000",
60260 => "1111111110110000",
60261 => "1111111110110000",
60262 => "1111111110110000",
60263 => "1111111110110000",
60264 => "1111111110110000",
60265 => "1111111110110000",
60266 => "1111111110110000",
60267 => "1111111110110000",
60268 => "1111111110110000",
60269 => "1111111110110000",
60270 => "1111111110110000",
60271 => "1111111110110000",
60272 => "1111111110110000",
60273 => "1111111110110000",
60274 => "1111111110110000",
60275 => "1111111110110000",
60276 => "1111111110110000",
60277 => "1111111110110000",
60278 => "1111111110110000",
60279 => "1111111110110000",
60280 => "1111111110110000",
60281 => "1111111110110000",
60282 => "1111111110110000",
60283 => "1111111110110000",
60284 => "1111111110110000",
60285 => "1111111110110000",
60286 => "1111111110110000",
60287 => "1111111110110000",
60288 => "1111111110110000",
60289 => "1111111110110000",
60290 => "1111111110110000",
60291 => "1111111110110001",
60292 => "1111111110110001",
60293 => "1111111110110001",
60294 => "1111111110110001",
60295 => "1111111110110001",
60296 => "1111111110110001",
60297 => "1111111110110001",
60298 => "1111111110110001",
60299 => "1111111110110001",
60300 => "1111111110110001",
60301 => "1111111110110001",
60302 => "1111111110110001",
60303 => "1111111110110001",
60304 => "1111111110110001",
60305 => "1111111110110001",
60306 => "1111111110110001",
60307 => "1111111110110001",
60308 => "1111111110110001",
60309 => "1111111110110001",
60310 => "1111111110110001",
60311 => "1111111110110001",
60312 => "1111111110110001",
60313 => "1111111110110001",
60314 => "1111111110110001",
60315 => "1111111110110001",
60316 => "1111111110110001",
60317 => "1111111110110001",
60318 => "1111111110110001",
60319 => "1111111110110001",
60320 => "1111111110110001",
60321 => "1111111110110001",
60322 => "1111111110110001",
60323 => "1111111110110001",
60324 => "1111111110110001",
60325 => "1111111110110001",
60326 => "1111111110110001",
60327 => "1111111110110001",
60328 => "1111111110110001",
60329 => "1111111110110001",
60330 => "1111111110110001",
60331 => "1111111110110001",
60332 => "1111111110110001",
60333 => "1111111110110001",
60334 => "1111111110110001",
60335 => "1111111110110001",
60336 => "1111111110110001",
60337 => "1111111110110001",
60338 => "1111111110110001",
60339 => "1111111110110001",
60340 => "1111111110110001",
60341 => "1111111110110001",
60342 => "1111111110110001",
60343 => "1111111110110001",
60344 => "1111111110110010",
60345 => "1111111110110010",
60346 => "1111111110110010",
60347 => "1111111110110010",
60348 => "1111111110110010",
60349 => "1111111110110010",
60350 => "1111111110110010",
60351 => "1111111110110010",
60352 => "1111111110110010",
60353 => "1111111110110010",
60354 => "1111111110110010",
60355 => "1111111110110010",
60356 => "1111111110110010",
60357 => "1111111110110010",
60358 => "1111111110110010",
60359 => "1111111110110010",
60360 => "1111111110110010",
60361 => "1111111110110010",
60362 => "1111111110110010",
60363 => "1111111110110010",
60364 => "1111111110110010",
60365 => "1111111110110010",
60366 => "1111111110110010",
60367 => "1111111110110010",
60368 => "1111111110110010",
60369 => "1111111110110010",
60370 => "1111111110110010",
60371 => "1111111110110010",
60372 => "1111111110110010",
60373 => "1111111110110010",
60374 => "1111111110110010",
60375 => "1111111110110010",
60376 => "1111111110110010",
60377 => "1111111110110010",
60378 => "1111111110110010",
60379 => "1111111110110010",
60380 => "1111111110110010",
60381 => "1111111110110010",
60382 => "1111111110110010",
60383 => "1111111110110010",
60384 => "1111111110110010",
60385 => "1111111110110010",
60386 => "1111111110110010",
60387 => "1111111110110010",
60388 => "1111111110110010",
60389 => "1111111110110010",
60390 => "1111111110110010",
60391 => "1111111110110010",
60392 => "1111111110110010",
60393 => "1111111110110010",
60394 => "1111111110110010",
60395 => "1111111110110010",
60396 => "1111111110110010",
60397 => "1111111110110011",
60398 => "1111111110110011",
60399 => "1111111110110011",
60400 => "1111111110110011",
60401 => "1111111110110011",
60402 => "1111111110110011",
60403 => "1111111110110011",
60404 => "1111111110110011",
60405 => "1111111110110011",
60406 => "1111111110110011",
60407 => "1111111110110011",
60408 => "1111111110110011",
60409 => "1111111110110011",
60410 => "1111111110110011",
60411 => "1111111110110011",
60412 => "1111111110110011",
60413 => "1111111110110011",
60414 => "1111111110110011",
60415 => "1111111110110011",
60416 => "1111111110110011",
60417 => "1111111110110011",
60418 => "1111111110110011",
60419 => "1111111110110011",
60420 => "1111111110110011",
60421 => "1111111110110011",
60422 => "1111111110110011",
60423 => "1111111110110011",
60424 => "1111111110110011",
60425 => "1111111110110011",
60426 => "1111111110110011",
60427 => "1111111110110011",
60428 => "1111111110110011",
60429 => "1111111110110011",
60430 => "1111111110110011",
60431 => "1111111110110011",
60432 => "1111111110110011",
60433 => "1111111110110011",
60434 => "1111111110110011",
60435 => "1111111110110011",
60436 => "1111111110110011",
60437 => "1111111110110011",
60438 => "1111111110110011",
60439 => "1111111110110011",
60440 => "1111111110110011",
60441 => "1111111110110011",
60442 => "1111111110110011",
60443 => "1111111110110011",
60444 => "1111111110110011",
60445 => "1111111110110011",
60446 => "1111111110110011",
60447 => "1111111110110011",
60448 => "1111111110110011",
60449 => "1111111110110011",
60450 => "1111111110110100",
60451 => "1111111110110100",
60452 => "1111111110110100",
60453 => "1111111110110100",
60454 => "1111111110110100",
60455 => "1111111110110100",
60456 => "1111111110110100",
60457 => "1111111110110100",
60458 => "1111111110110100",
60459 => "1111111110110100",
60460 => "1111111110110100",
60461 => "1111111110110100",
60462 => "1111111110110100",
60463 => "1111111110110100",
60464 => "1111111110110100",
60465 => "1111111110110100",
60466 => "1111111110110100",
60467 => "1111111110110100",
60468 => "1111111110110100",
60469 => "1111111110110100",
60470 => "1111111110110100",
60471 => "1111111110110100",
60472 => "1111111110110100",
60473 => "1111111110110100",
60474 => "1111111110110100",
60475 => "1111111110110100",
60476 => "1111111110110100",
60477 => "1111111110110100",
60478 => "1111111110110100",
60479 => "1111111110110100",
60480 => "1111111110110100",
60481 => "1111111110110100",
60482 => "1111111110110100",
60483 => "1111111110110100",
60484 => "1111111110110100",
60485 => "1111111110110100",
60486 => "1111111110110100",
60487 => "1111111110110100",
60488 => "1111111110110100",
60489 => "1111111110110100",
60490 => "1111111110110100",
60491 => "1111111110110100",
60492 => "1111111110110100",
60493 => "1111111110110100",
60494 => "1111111110110100",
60495 => "1111111110110100",
60496 => "1111111110110100",
60497 => "1111111110110100",
60498 => "1111111110110100",
60499 => "1111111110110100",
60500 => "1111111110110100",
60501 => "1111111110110100",
60502 => "1111111110110100",
60503 => "1111111110110100",
60504 => "1111111110110100",
60505 => "1111111110110101",
60506 => "1111111110110101",
60507 => "1111111110110101",
60508 => "1111111110110101",
60509 => "1111111110110101",
60510 => "1111111110110101",
60511 => "1111111110110101",
60512 => "1111111110110101",
60513 => "1111111110110101",
60514 => "1111111110110101",
60515 => "1111111110110101",
60516 => "1111111110110101",
60517 => "1111111110110101",
60518 => "1111111110110101",
60519 => "1111111110110101",
60520 => "1111111110110101",
60521 => "1111111110110101",
60522 => "1111111110110101",
60523 => "1111111110110101",
60524 => "1111111110110101",
60525 => "1111111110110101",
60526 => "1111111110110101",
60527 => "1111111110110101",
60528 => "1111111110110101",
60529 => "1111111110110101",
60530 => "1111111110110101",
60531 => "1111111110110101",
60532 => "1111111110110101",
60533 => "1111111110110101",
60534 => "1111111110110101",
60535 => "1111111110110101",
60536 => "1111111110110101",
60537 => "1111111110110101",
60538 => "1111111110110101",
60539 => "1111111110110101",
60540 => "1111111110110101",
60541 => "1111111110110101",
60542 => "1111111110110101",
60543 => "1111111110110101",
60544 => "1111111110110101",
60545 => "1111111110110101",
60546 => "1111111110110101",
60547 => "1111111110110101",
60548 => "1111111110110101",
60549 => "1111111110110101",
60550 => "1111111110110101",
60551 => "1111111110110101",
60552 => "1111111110110101",
60553 => "1111111110110101",
60554 => "1111111110110101",
60555 => "1111111110110101",
60556 => "1111111110110101",
60557 => "1111111110110101",
60558 => "1111111110110101",
60559 => "1111111110110101",
60560 => "1111111110110110",
60561 => "1111111110110110",
60562 => "1111111110110110",
60563 => "1111111110110110",
60564 => "1111111110110110",
60565 => "1111111110110110",
60566 => "1111111110110110",
60567 => "1111111110110110",
60568 => "1111111110110110",
60569 => "1111111110110110",
60570 => "1111111110110110",
60571 => "1111111110110110",
60572 => "1111111110110110",
60573 => "1111111110110110",
60574 => "1111111110110110",
60575 => "1111111110110110",
60576 => "1111111110110110",
60577 => "1111111110110110",
60578 => "1111111110110110",
60579 => "1111111110110110",
60580 => "1111111110110110",
60581 => "1111111110110110",
60582 => "1111111110110110",
60583 => "1111111110110110",
60584 => "1111111110110110",
60585 => "1111111110110110",
60586 => "1111111110110110",
60587 => "1111111110110110",
60588 => "1111111110110110",
60589 => "1111111110110110",
60590 => "1111111110110110",
60591 => "1111111110110110",
60592 => "1111111110110110",
60593 => "1111111110110110",
60594 => "1111111110110110",
60595 => "1111111110110110",
60596 => "1111111110110110",
60597 => "1111111110110110",
60598 => "1111111110110110",
60599 => "1111111110110110",
60600 => "1111111110110110",
60601 => "1111111110110110",
60602 => "1111111110110110",
60603 => "1111111110110110",
60604 => "1111111110110110",
60605 => "1111111110110110",
60606 => "1111111110110110",
60607 => "1111111110110110",
60608 => "1111111110110110",
60609 => "1111111110110110",
60610 => "1111111110110110",
60611 => "1111111110110110",
60612 => "1111111110110110",
60613 => "1111111110110110",
60614 => "1111111110110110",
60615 => "1111111110110111",
60616 => "1111111110110111",
60617 => "1111111110110111",
60618 => "1111111110110111",
60619 => "1111111110110111",
60620 => "1111111110110111",
60621 => "1111111110110111",
60622 => "1111111110110111",
60623 => "1111111110110111",
60624 => "1111111110110111",
60625 => "1111111110110111",
60626 => "1111111110110111",
60627 => "1111111110110111",
60628 => "1111111110110111",
60629 => "1111111110110111",
60630 => "1111111110110111",
60631 => "1111111110110111",
60632 => "1111111110110111",
60633 => "1111111110110111",
60634 => "1111111110110111",
60635 => "1111111110110111",
60636 => "1111111110110111",
60637 => "1111111110110111",
60638 => "1111111110110111",
60639 => "1111111110110111",
60640 => "1111111110110111",
60641 => "1111111110110111",
60642 => "1111111110110111",
60643 => "1111111110110111",
60644 => "1111111110110111",
60645 => "1111111110110111",
60646 => "1111111110110111",
60647 => "1111111110110111",
60648 => "1111111110110111",
60649 => "1111111110110111",
60650 => "1111111110110111",
60651 => "1111111110110111",
60652 => "1111111110110111",
60653 => "1111111110110111",
60654 => "1111111110110111",
60655 => "1111111110110111",
60656 => "1111111110110111",
60657 => "1111111110110111",
60658 => "1111111110110111",
60659 => "1111111110110111",
60660 => "1111111110110111",
60661 => "1111111110110111",
60662 => "1111111110110111",
60663 => "1111111110110111",
60664 => "1111111110110111",
60665 => "1111111110110111",
60666 => "1111111110110111",
60667 => "1111111110110111",
60668 => "1111111110110111",
60669 => "1111111110110111",
60670 => "1111111110110111",
60671 => "1111111110110111",
60672 => "1111111110111000",
60673 => "1111111110111000",
60674 => "1111111110111000",
60675 => "1111111110111000",
60676 => "1111111110111000",
60677 => "1111111110111000",
60678 => "1111111110111000",
60679 => "1111111110111000",
60680 => "1111111110111000",
60681 => "1111111110111000",
60682 => "1111111110111000",
60683 => "1111111110111000",
60684 => "1111111110111000",
60685 => "1111111110111000",
60686 => "1111111110111000",
60687 => "1111111110111000",
60688 => "1111111110111000",
60689 => "1111111110111000",
60690 => "1111111110111000",
60691 => "1111111110111000",
60692 => "1111111110111000",
60693 => "1111111110111000",
60694 => "1111111110111000",
60695 => "1111111110111000",
60696 => "1111111110111000",
60697 => "1111111110111000",
60698 => "1111111110111000",
60699 => "1111111110111000",
60700 => "1111111110111000",
60701 => "1111111110111000",
60702 => "1111111110111000",
60703 => "1111111110111000",
60704 => "1111111110111000",
60705 => "1111111110111000",
60706 => "1111111110111000",
60707 => "1111111110111000",
60708 => "1111111110111000",
60709 => "1111111110111000",
60710 => "1111111110111000",
60711 => "1111111110111000",
60712 => "1111111110111000",
60713 => "1111111110111000",
60714 => "1111111110111000",
60715 => "1111111110111000",
60716 => "1111111110111000",
60717 => "1111111110111000",
60718 => "1111111110111000",
60719 => "1111111110111000",
60720 => "1111111110111000",
60721 => "1111111110111000",
60722 => "1111111110111000",
60723 => "1111111110111000",
60724 => "1111111110111000",
60725 => "1111111110111000",
60726 => "1111111110111000",
60727 => "1111111110111000",
60728 => "1111111110111000",
60729 => "1111111110111001",
60730 => "1111111110111001",
60731 => "1111111110111001",
60732 => "1111111110111001",
60733 => "1111111110111001",
60734 => "1111111110111001",
60735 => "1111111110111001",
60736 => "1111111110111001",
60737 => "1111111110111001",
60738 => "1111111110111001",
60739 => "1111111110111001",
60740 => "1111111110111001",
60741 => "1111111110111001",
60742 => "1111111110111001",
60743 => "1111111110111001",
60744 => "1111111110111001",
60745 => "1111111110111001",
60746 => "1111111110111001",
60747 => "1111111110111001",
60748 => "1111111110111001",
60749 => "1111111110111001",
60750 => "1111111110111001",
60751 => "1111111110111001",
60752 => "1111111110111001",
60753 => "1111111110111001",
60754 => "1111111110111001",
60755 => "1111111110111001",
60756 => "1111111110111001",
60757 => "1111111110111001",
60758 => "1111111110111001",
60759 => "1111111110111001",
60760 => "1111111110111001",
60761 => "1111111110111001",
60762 => "1111111110111001",
60763 => "1111111110111001",
60764 => "1111111110111001",
60765 => "1111111110111001",
60766 => "1111111110111001",
60767 => "1111111110111001",
60768 => "1111111110111001",
60769 => "1111111110111001",
60770 => "1111111110111001",
60771 => "1111111110111001",
60772 => "1111111110111001",
60773 => "1111111110111001",
60774 => "1111111110111001",
60775 => "1111111110111001",
60776 => "1111111110111001",
60777 => "1111111110111001",
60778 => "1111111110111001",
60779 => "1111111110111001",
60780 => "1111111110111001",
60781 => "1111111110111001",
60782 => "1111111110111001",
60783 => "1111111110111001",
60784 => "1111111110111001",
60785 => "1111111110111001",
60786 => "1111111110111001",
60787 => "1111111110111010",
60788 => "1111111110111010",
60789 => "1111111110111010",
60790 => "1111111110111010",
60791 => "1111111110111010",
60792 => "1111111110111010",
60793 => "1111111110111010",
60794 => "1111111110111010",
60795 => "1111111110111010",
60796 => "1111111110111010",
60797 => "1111111110111010",
60798 => "1111111110111010",
60799 => "1111111110111010",
60800 => "1111111110111010",
60801 => "1111111110111010",
60802 => "1111111110111010",
60803 => "1111111110111010",
60804 => "1111111110111010",
60805 => "1111111110111010",
60806 => "1111111110111010",
60807 => "1111111110111010",
60808 => "1111111110111010",
60809 => "1111111110111010",
60810 => "1111111110111010",
60811 => "1111111110111010",
60812 => "1111111110111010",
60813 => "1111111110111010",
60814 => "1111111110111010",
60815 => "1111111110111010",
60816 => "1111111110111010",
60817 => "1111111110111010",
60818 => "1111111110111010",
60819 => "1111111110111010",
60820 => "1111111110111010",
60821 => "1111111110111010",
60822 => "1111111110111010",
60823 => "1111111110111010",
60824 => "1111111110111010",
60825 => "1111111110111010",
60826 => "1111111110111010",
60827 => "1111111110111010",
60828 => "1111111110111010",
60829 => "1111111110111010",
60830 => "1111111110111010",
60831 => "1111111110111010",
60832 => "1111111110111010",
60833 => "1111111110111010",
60834 => "1111111110111010",
60835 => "1111111110111010",
60836 => "1111111110111010",
60837 => "1111111110111010",
60838 => "1111111110111010",
60839 => "1111111110111010",
60840 => "1111111110111010",
60841 => "1111111110111010",
60842 => "1111111110111010",
60843 => "1111111110111010",
60844 => "1111111110111010",
60845 => "1111111110111010",
60846 => "1111111110111011",
60847 => "1111111110111011",
60848 => "1111111110111011",
60849 => "1111111110111011",
60850 => "1111111110111011",
60851 => "1111111110111011",
60852 => "1111111110111011",
60853 => "1111111110111011",
60854 => "1111111110111011",
60855 => "1111111110111011",
60856 => "1111111110111011",
60857 => "1111111110111011",
60858 => "1111111110111011",
60859 => "1111111110111011",
60860 => "1111111110111011",
60861 => "1111111110111011",
60862 => "1111111110111011",
60863 => "1111111110111011",
60864 => "1111111110111011",
60865 => "1111111110111011",
60866 => "1111111110111011",
60867 => "1111111110111011",
60868 => "1111111110111011",
60869 => "1111111110111011",
60870 => "1111111110111011",
60871 => "1111111110111011",
60872 => "1111111110111011",
60873 => "1111111110111011",
60874 => "1111111110111011",
60875 => "1111111110111011",
60876 => "1111111110111011",
60877 => "1111111110111011",
60878 => "1111111110111011",
60879 => "1111111110111011",
60880 => "1111111110111011",
60881 => "1111111110111011",
60882 => "1111111110111011",
60883 => "1111111110111011",
60884 => "1111111110111011",
60885 => "1111111110111011",
60886 => "1111111110111011",
60887 => "1111111110111011",
60888 => "1111111110111011",
60889 => "1111111110111011",
60890 => "1111111110111011",
60891 => "1111111110111011",
60892 => "1111111110111011",
60893 => "1111111110111011",
60894 => "1111111110111011",
60895 => "1111111110111011",
60896 => "1111111110111011",
60897 => "1111111110111011",
60898 => "1111111110111011",
60899 => "1111111110111011",
60900 => "1111111110111011",
60901 => "1111111110111011",
60902 => "1111111110111011",
60903 => "1111111110111011",
60904 => "1111111110111011",
60905 => "1111111110111011",
60906 => "1111111110111100",
60907 => "1111111110111100",
60908 => "1111111110111100",
60909 => "1111111110111100",
60910 => "1111111110111100",
60911 => "1111111110111100",
60912 => "1111111110111100",
60913 => "1111111110111100",
60914 => "1111111110111100",
60915 => "1111111110111100",
60916 => "1111111110111100",
60917 => "1111111110111100",
60918 => "1111111110111100",
60919 => "1111111110111100",
60920 => "1111111110111100",
60921 => "1111111110111100",
60922 => "1111111110111100",
60923 => "1111111110111100",
60924 => "1111111110111100",
60925 => "1111111110111100",
60926 => "1111111110111100",
60927 => "1111111110111100",
60928 => "1111111110111100",
60929 => "1111111110111100",
60930 => "1111111110111100",
60931 => "1111111110111100",
60932 => "1111111110111100",
60933 => "1111111110111100",
60934 => "1111111110111100",
60935 => "1111111110111100",
60936 => "1111111110111100",
60937 => "1111111110111100",
60938 => "1111111110111100",
60939 => "1111111110111100",
60940 => "1111111110111100",
60941 => "1111111110111100",
60942 => "1111111110111100",
60943 => "1111111110111100",
60944 => "1111111110111100",
60945 => "1111111110111100",
60946 => "1111111110111100",
60947 => "1111111110111100",
60948 => "1111111110111100",
60949 => "1111111110111100",
60950 => "1111111110111100",
60951 => "1111111110111100",
60952 => "1111111110111100",
60953 => "1111111110111100",
60954 => "1111111110111100",
60955 => "1111111110111100",
60956 => "1111111110111100",
60957 => "1111111110111100",
60958 => "1111111110111100",
60959 => "1111111110111100",
60960 => "1111111110111100",
60961 => "1111111110111100",
60962 => "1111111110111100",
60963 => "1111111110111100",
60964 => "1111111110111100",
60965 => "1111111110111100",
60966 => "1111111110111100",
60967 => "1111111110111101",
60968 => "1111111110111101",
60969 => "1111111110111101",
60970 => "1111111110111101",
60971 => "1111111110111101",
60972 => "1111111110111101",
60973 => "1111111110111101",
60974 => "1111111110111101",
60975 => "1111111110111101",
60976 => "1111111110111101",
60977 => "1111111110111101",
60978 => "1111111110111101",
60979 => "1111111110111101",
60980 => "1111111110111101",
60981 => "1111111110111101",
60982 => "1111111110111101",
60983 => "1111111110111101",
60984 => "1111111110111101",
60985 => "1111111110111101",
60986 => "1111111110111101",
60987 => "1111111110111101",
60988 => "1111111110111101",
60989 => "1111111110111101",
60990 => "1111111110111101",
60991 => "1111111110111101",
60992 => "1111111110111101",
60993 => "1111111110111101",
60994 => "1111111110111101",
60995 => "1111111110111101",
60996 => "1111111110111101",
60997 => "1111111110111101",
60998 => "1111111110111101",
60999 => "1111111110111101",
61000 => "1111111110111101",
61001 => "1111111110111101",
61002 => "1111111110111101",
61003 => "1111111110111101",
61004 => "1111111110111101",
61005 => "1111111110111101",
61006 => "1111111110111101",
61007 => "1111111110111101",
61008 => "1111111110111101",
61009 => "1111111110111101",
61010 => "1111111110111101",
61011 => "1111111110111101",
61012 => "1111111110111101",
61013 => "1111111110111101",
61014 => "1111111110111101",
61015 => "1111111110111101",
61016 => "1111111110111101",
61017 => "1111111110111101",
61018 => "1111111110111101",
61019 => "1111111110111101",
61020 => "1111111110111101",
61021 => "1111111110111101",
61022 => "1111111110111101",
61023 => "1111111110111101",
61024 => "1111111110111101",
61025 => "1111111110111101",
61026 => "1111111110111101",
61027 => "1111111110111101",
61028 => "1111111110111101",
61029 => "1111111110111110",
61030 => "1111111110111110",
61031 => "1111111110111110",
61032 => "1111111110111110",
61033 => "1111111110111110",
61034 => "1111111110111110",
61035 => "1111111110111110",
61036 => "1111111110111110",
61037 => "1111111110111110",
61038 => "1111111110111110",
61039 => "1111111110111110",
61040 => "1111111110111110",
61041 => "1111111110111110",
61042 => "1111111110111110",
61043 => "1111111110111110",
61044 => "1111111110111110",
61045 => "1111111110111110",
61046 => "1111111110111110",
61047 => "1111111110111110",
61048 => "1111111110111110",
61049 => "1111111110111110",
61050 => "1111111110111110",
61051 => "1111111110111110",
61052 => "1111111110111110",
61053 => "1111111110111110",
61054 => "1111111110111110",
61055 => "1111111110111110",
61056 => "1111111110111110",
61057 => "1111111110111110",
61058 => "1111111110111110",
61059 => "1111111110111110",
61060 => "1111111110111110",
61061 => "1111111110111110",
61062 => "1111111110111110",
61063 => "1111111110111110",
61064 => "1111111110111110",
61065 => "1111111110111110",
61066 => "1111111110111110",
61067 => "1111111110111110",
61068 => "1111111110111110",
61069 => "1111111110111110",
61070 => "1111111110111110",
61071 => "1111111110111110",
61072 => "1111111110111110",
61073 => "1111111110111110",
61074 => "1111111110111110",
61075 => "1111111110111110",
61076 => "1111111110111110",
61077 => "1111111110111110",
61078 => "1111111110111110",
61079 => "1111111110111110",
61080 => "1111111110111110",
61081 => "1111111110111110",
61082 => "1111111110111110",
61083 => "1111111110111110",
61084 => "1111111110111110",
61085 => "1111111110111110",
61086 => "1111111110111110",
61087 => "1111111110111110",
61088 => "1111111110111110",
61089 => "1111111110111110",
61090 => "1111111110111110",
61091 => "1111111110111111",
61092 => "1111111110111111",
61093 => "1111111110111111",
61094 => "1111111110111111",
61095 => "1111111110111111",
61096 => "1111111110111111",
61097 => "1111111110111111",
61098 => "1111111110111111",
61099 => "1111111110111111",
61100 => "1111111110111111",
61101 => "1111111110111111",
61102 => "1111111110111111",
61103 => "1111111110111111",
61104 => "1111111110111111",
61105 => "1111111110111111",
61106 => "1111111110111111",
61107 => "1111111110111111",
61108 => "1111111110111111",
61109 => "1111111110111111",
61110 => "1111111110111111",
61111 => "1111111110111111",
61112 => "1111111110111111",
61113 => "1111111110111111",
61114 => "1111111110111111",
61115 => "1111111110111111",
61116 => "1111111110111111",
61117 => "1111111110111111",
61118 => "1111111110111111",
61119 => "1111111110111111",
61120 => "1111111110111111",
61121 => "1111111110111111",
61122 => "1111111110111111",
61123 => "1111111110111111",
61124 => "1111111110111111",
61125 => "1111111110111111",
61126 => "1111111110111111",
61127 => "1111111110111111",
61128 => "1111111110111111",
61129 => "1111111110111111",
61130 => "1111111110111111",
61131 => "1111111110111111",
61132 => "1111111110111111",
61133 => "1111111110111111",
61134 => "1111111110111111",
61135 => "1111111110111111",
61136 => "1111111110111111",
61137 => "1111111110111111",
61138 => "1111111110111111",
61139 => "1111111110111111",
61140 => "1111111110111111",
61141 => "1111111110111111",
61142 => "1111111110111111",
61143 => "1111111110111111",
61144 => "1111111110111111",
61145 => "1111111110111111",
61146 => "1111111110111111",
61147 => "1111111110111111",
61148 => "1111111110111111",
61149 => "1111111110111111",
61150 => "1111111110111111",
61151 => "1111111110111111",
61152 => "1111111110111111",
61153 => "1111111110111111",
61154 => "1111111110111111",
61155 => "1111111111000000",
61156 => "1111111111000000",
61157 => "1111111111000000",
61158 => "1111111111000000",
61159 => "1111111111000000",
61160 => "1111111111000000",
61161 => "1111111111000000",
61162 => "1111111111000000",
61163 => "1111111111000000",
61164 => "1111111111000000",
61165 => "1111111111000000",
61166 => "1111111111000000",
61167 => "1111111111000000",
61168 => "1111111111000000",
61169 => "1111111111000000",
61170 => "1111111111000000",
61171 => "1111111111000000",
61172 => "1111111111000000",
61173 => "1111111111000000",
61174 => "1111111111000000",
61175 => "1111111111000000",
61176 => "1111111111000000",
61177 => "1111111111000000",
61178 => "1111111111000000",
61179 => "1111111111000000",
61180 => "1111111111000000",
61181 => "1111111111000000",
61182 => "1111111111000000",
61183 => "1111111111000000",
61184 => "1111111111000000",
61185 => "1111111111000000",
61186 => "1111111111000000",
61187 => "1111111111000000",
61188 => "1111111111000000",
61189 => "1111111111000000",
61190 => "1111111111000000",
61191 => "1111111111000000",
61192 => "1111111111000000",
61193 => "1111111111000000",
61194 => "1111111111000000",
61195 => "1111111111000000",
61196 => "1111111111000000",
61197 => "1111111111000000",
61198 => "1111111111000000",
61199 => "1111111111000000",
61200 => "1111111111000000",
61201 => "1111111111000000",
61202 => "1111111111000000",
61203 => "1111111111000000",
61204 => "1111111111000000",
61205 => "1111111111000000",
61206 => "1111111111000000",
61207 => "1111111111000000",
61208 => "1111111111000000",
61209 => "1111111111000000",
61210 => "1111111111000000",
61211 => "1111111111000000",
61212 => "1111111111000000",
61213 => "1111111111000000",
61214 => "1111111111000000",
61215 => "1111111111000000",
61216 => "1111111111000000",
61217 => "1111111111000000",
61218 => "1111111111000000",
61219 => "1111111111000001",
61220 => "1111111111000001",
61221 => "1111111111000001",
61222 => "1111111111000001",
61223 => "1111111111000001",
61224 => "1111111111000001",
61225 => "1111111111000001",
61226 => "1111111111000001",
61227 => "1111111111000001",
61228 => "1111111111000001",
61229 => "1111111111000001",
61230 => "1111111111000001",
61231 => "1111111111000001",
61232 => "1111111111000001",
61233 => "1111111111000001",
61234 => "1111111111000001",
61235 => "1111111111000001",
61236 => "1111111111000001",
61237 => "1111111111000001",
61238 => "1111111111000001",
61239 => "1111111111000001",
61240 => "1111111111000001",
61241 => "1111111111000001",
61242 => "1111111111000001",
61243 => "1111111111000001",
61244 => "1111111111000001",
61245 => "1111111111000001",
61246 => "1111111111000001",
61247 => "1111111111000001",
61248 => "1111111111000001",
61249 => "1111111111000001",
61250 => "1111111111000001",
61251 => "1111111111000001",
61252 => "1111111111000001",
61253 => "1111111111000001",
61254 => "1111111111000001",
61255 => "1111111111000001",
61256 => "1111111111000001",
61257 => "1111111111000001",
61258 => "1111111111000001",
61259 => "1111111111000001",
61260 => "1111111111000001",
61261 => "1111111111000001",
61262 => "1111111111000001",
61263 => "1111111111000001",
61264 => "1111111111000001",
61265 => "1111111111000001",
61266 => "1111111111000001",
61267 => "1111111111000001",
61268 => "1111111111000001",
61269 => "1111111111000001",
61270 => "1111111111000001",
61271 => "1111111111000001",
61272 => "1111111111000001",
61273 => "1111111111000001",
61274 => "1111111111000001",
61275 => "1111111111000001",
61276 => "1111111111000001",
61277 => "1111111111000001",
61278 => "1111111111000001",
61279 => "1111111111000001",
61280 => "1111111111000001",
61281 => "1111111111000001",
61282 => "1111111111000001",
61283 => "1111111111000001",
61284 => "1111111111000001",
61285 => "1111111111000010",
61286 => "1111111111000010",
61287 => "1111111111000010",
61288 => "1111111111000010",
61289 => "1111111111000010",
61290 => "1111111111000010",
61291 => "1111111111000010",
61292 => "1111111111000010",
61293 => "1111111111000010",
61294 => "1111111111000010",
61295 => "1111111111000010",
61296 => "1111111111000010",
61297 => "1111111111000010",
61298 => "1111111111000010",
61299 => "1111111111000010",
61300 => "1111111111000010",
61301 => "1111111111000010",
61302 => "1111111111000010",
61303 => "1111111111000010",
61304 => "1111111111000010",
61305 => "1111111111000010",
61306 => "1111111111000010",
61307 => "1111111111000010",
61308 => "1111111111000010",
61309 => "1111111111000010",
61310 => "1111111111000010",
61311 => "1111111111000010",
61312 => "1111111111000010",
61313 => "1111111111000010",
61314 => "1111111111000010",
61315 => "1111111111000010",
61316 => "1111111111000010",
61317 => "1111111111000010",
61318 => "1111111111000010",
61319 => "1111111111000010",
61320 => "1111111111000010",
61321 => "1111111111000010",
61322 => "1111111111000010",
61323 => "1111111111000010",
61324 => "1111111111000010",
61325 => "1111111111000010",
61326 => "1111111111000010",
61327 => "1111111111000010",
61328 => "1111111111000010",
61329 => "1111111111000010",
61330 => "1111111111000010",
61331 => "1111111111000010",
61332 => "1111111111000010",
61333 => "1111111111000010",
61334 => "1111111111000010",
61335 => "1111111111000010",
61336 => "1111111111000010",
61337 => "1111111111000010",
61338 => "1111111111000010",
61339 => "1111111111000010",
61340 => "1111111111000010",
61341 => "1111111111000010",
61342 => "1111111111000010",
61343 => "1111111111000010",
61344 => "1111111111000010",
61345 => "1111111111000010",
61346 => "1111111111000010",
61347 => "1111111111000010",
61348 => "1111111111000010",
61349 => "1111111111000010",
61350 => "1111111111000010",
61351 => "1111111111000010",
61352 => "1111111111000011",
61353 => "1111111111000011",
61354 => "1111111111000011",
61355 => "1111111111000011",
61356 => "1111111111000011",
61357 => "1111111111000011",
61358 => "1111111111000011",
61359 => "1111111111000011",
61360 => "1111111111000011",
61361 => "1111111111000011",
61362 => "1111111111000011",
61363 => "1111111111000011",
61364 => "1111111111000011",
61365 => "1111111111000011",
61366 => "1111111111000011",
61367 => "1111111111000011",
61368 => "1111111111000011",
61369 => "1111111111000011",
61370 => "1111111111000011",
61371 => "1111111111000011",
61372 => "1111111111000011",
61373 => "1111111111000011",
61374 => "1111111111000011",
61375 => "1111111111000011",
61376 => "1111111111000011",
61377 => "1111111111000011",
61378 => "1111111111000011",
61379 => "1111111111000011",
61380 => "1111111111000011",
61381 => "1111111111000011",
61382 => "1111111111000011",
61383 => "1111111111000011",
61384 => "1111111111000011",
61385 => "1111111111000011",
61386 => "1111111111000011",
61387 => "1111111111000011",
61388 => "1111111111000011",
61389 => "1111111111000011",
61390 => "1111111111000011",
61391 => "1111111111000011",
61392 => "1111111111000011",
61393 => "1111111111000011",
61394 => "1111111111000011",
61395 => "1111111111000011",
61396 => "1111111111000011",
61397 => "1111111111000011",
61398 => "1111111111000011",
61399 => "1111111111000011",
61400 => "1111111111000011",
61401 => "1111111111000011",
61402 => "1111111111000011",
61403 => "1111111111000011",
61404 => "1111111111000011",
61405 => "1111111111000011",
61406 => "1111111111000011",
61407 => "1111111111000011",
61408 => "1111111111000011",
61409 => "1111111111000011",
61410 => "1111111111000011",
61411 => "1111111111000011",
61412 => "1111111111000011",
61413 => "1111111111000011",
61414 => "1111111111000011",
61415 => "1111111111000011",
61416 => "1111111111000011",
61417 => "1111111111000011",
61418 => "1111111111000011",
61419 => "1111111111000100",
61420 => "1111111111000100",
61421 => "1111111111000100",
61422 => "1111111111000100",
61423 => "1111111111000100",
61424 => "1111111111000100",
61425 => "1111111111000100",
61426 => "1111111111000100",
61427 => "1111111111000100",
61428 => "1111111111000100",
61429 => "1111111111000100",
61430 => "1111111111000100",
61431 => "1111111111000100",
61432 => "1111111111000100",
61433 => "1111111111000100",
61434 => "1111111111000100",
61435 => "1111111111000100",
61436 => "1111111111000100",
61437 => "1111111111000100",
61438 => "1111111111000100",
61439 => "1111111111000100",
61440 => "1111111111000100",
61441 => "1111111111000100",
61442 => "1111111111000100",
61443 => "1111111111000100",
61444 => "1111111111000100",
61445 => "1111111111000100",
61446 => "1111111111000100",
61447 => "1111111111000100",
61448 => "1111111111000100",
61449 => "1111111111000100",
61450 => "1111111111000100",
61451 => "1111111111000100",
61452 => "1111111111000100",
61453 => "1111111111000100",
61454 => "1111111111000100",
61455 => "1111111111000100",
61456 => "1111111111000100",
61457 => "1111111111000100",
61458 => "1111111111000100",
61459 => "1111111111000100",
61460 => "1111111111000100",
61461 => "1111111111000100",
61462 => "1111111111000100",
61463 => "1111111111000100",
61464 => "1111111111000100",
61465 => "1111111111000100",
61466 => "1111111111000100",
61467 => "1111111111000100",
61468 => "1111111111000100",
61469 => "1111111111000100",
61470 => "1111111111000100",
61471 => "1111111111000100",
61472 => "1111111111000100",
61473 => "1111111111000100",
61474 => "1111111111000100",
61475 => "1111111111000100",
61476 => "1111111111000100",
61477 => "1111111111000100",
61478 => "1111111111000100",
61479 => "1111111111000100",
61480 => "1111111111000100",
61481 => "1111111111000100",
61482 => "1111111111000100",
61483 => "1111111111000100",
61484 => "1111111111000100",
61485 => "1111111111000100",
61486 => "1111111111000100",
61487 => "1111111111000100",
61488 => "1111111111000101",
61489 => "1111111111000101",
61490 => "1111111111000101",
61491 => "1111111111000101",
61492 => "1111111111000101",
61493 => "1111111111000101",
61494 => "1111111111000101",
61495 => "1111111111000101",
61496 => "1111111111000101",
61497 => "1111111111000101",
61498 => "1111111111000101",
61499 => "1111111111000101",
61500 => "1111111111000101",
61501 => "1111111111000101",
61502 => "1111111111000101",
61503 => "1111111111000101",
61504 => "1111111111000101",
61505 => "1111111111000101",
61506 => "1111111111000101",
61507 => "1111111111000101",
61508 => "1111111111000101",
61509 => "1111111111000101",
61510 => "1111111111000101",
61511 => "1111111111000101",
61512 => "1111111111000101",
61513 => "1111111111000101",
61514 => "1111111111000101",
61515 => "1111111111000101",
61516 => "1111111111000101",
61517 => "1111111111000101",
61518 => "1111111111000101",
61519 => "1111111111000101",
61520 => "1111111111000101",
61521 => "1111111111000101",
61522 => "1111111111000101",
61523 => "1111111111000101",
61524 => "1111111111000101",
61525 => "1111111111000101",
61526 => "1111111111000101",
61527 => "1111111111000101",
61528 => "1111111111000101",
61529 => "1111111111000101",
61530 => "1111111111000101",
61531 => "1111111111000101",
61532 => "1111111111000101",
61533 => "1111111111000101",
61534 => "1111111111000101",
61535 => "1111111111000101",
61536 => "1111111111000101",
61537 => "1111111111000101",
61538 => "1111111111000101",
61539 => "1111111111000101",
61540 => "1111111111000101",
61541 => "1111111111000101",
61542 => "1111111111000101",
61543 => "1111111111000101",
61544 => "1111111111000101",
61545 => "1111111111000101",
61546 => "1111111111000101",
61547 => "1111111111000101",
61548 => "1111111111000101",
61549 => "1111111111000101",
61550 => "1111111111000101",
61551 => "1111111111000101",
61552 => "1111111111000101",
61553 => "1111111111000101",
61554 => "1111111111000101",
61555 => "1111111111000101",
61556 => "1111111111000101",
61557 => "1111111111000101",
61558 => "1111111111000110",
61559 => "1111111111000110",
61560 => "1111111111000110",
61561 => "1111111111000110",
61562 => "1111111111000110",
61563 => "1111111111000110",
61564 => "1111111111000110",
61565 => "1111111111000110",
61566 => "1111111111000110",
61567 => "1111111111000110",
61568 => "1111111111000110",
61569 => "1111111111000110",
61570 => "1111111111000110",
61571 => "1111111111000110",
61572 => "1111111111000110",
61573 => "1111111111000110",
61574 => "1111111111000110",
61575 => "1111111111000110",
61576 => "1111111111000110",
61577 => "1111111111000110",
61578 => "1111111111000110",
61579 => "1111111111000110",
61580 => "1111111111000110",
61581 => "1111111111000110",
61582 => "1111111111000110",
61583 => "1111111111000110",
61584 => "1111111111000110",
61585 => "1111111111000110",
61586 => "1111111111000110",
61587 => "1111111111000110",
61588 => "1111111111000110",
61589 => "1111111111000110",
61590 => "1111111111000110",
61591 => "1111111111000110",
61592 => "1111111111000110",
61593 => "1111111111000110",
61594 => "1111111111000110",
61595 => "1111111111000110",
61596 => "1111111111000110",
61597 => "1111111111000110",
61598 => "1111111111000110",
61599 => "1111111111000110",
61600 => "1111111111000110",
61601 => "1111111111000110",
61602 => "1111111111000110",
61603 => "1111111111000110",
61604 => "1111111111000110",
61605 => "1111111111000110",
61606 => "1111111111000110",
61607 => "1111111111000110",
61608 => "1111111111000110",
61609 => "1111111111000110",
61610 => "1111111111000110",
61611 => "1111111111000110",
61612 => "1111111111000110",
61613 => "1111111111000110",
61614 => "1111111111000110",
61615 => "1111111111000110",
61616 => "1111111111000110",
61617 => "1111111111000110",
61618 => "1111111111000110",
61619 => "1111111111000110",
61620 => "1111111111000110",
61621 => "1111111111000110",
61622 => "1111111111000110",
61623 => "1111111111000110",
61624 => "1111111111000110",
61625 => "1111111111000110",
61626 => "1111111111000110",
61627 => "1111111111000110",
61628 => "1111111111000110",
61629 => "1111111111000110",
61630 => "1111111111000111",
61631 => "1111111111000111",
61632 => "1111111111000111",
61633 => "1111111111000111",
61634 => "1111111111000111",
61635 => "1111111111000111",
61636 => "1111111111000111",
61637 => "1111111111000111",
61638 => "1111111111000111",
61639 => "1111111111000111",
61640 => "1111111111000111",
61641 => "1111111111000111",
61642 => "1111111111000111",
61643 => "1111111111000111",
61644 => "1111111111000111",
61645 => "1111111111000111",
61646 => "1111111111000111",
61647 => "1111111111000111",
61648 => "1111111111000111",
61649 => "1111111111000111",
61650 => "1111111111000111",
61651 => "1111111111000111",
61652 => "1111111111000111",
61653 => "1111111111000111",
61654 => "1111111111000111",
61655 => "1111111111000111",
61656 => "1111111111000111",
61657 => "1111111111000111",
61658 => "1111111111000111",
61659 => "1111111111000111",
61660 => "1111111111000111",
61661 => "1111111111000111",
61662 => "1111111111000111",
61663 => "1111111111000111",
61664 => "1111111111000111",
61665 => "1111111111000111",
61666 => "1111111111000111",
61667 => "1111111111000111",
61668 => "1111111111000111",
61669 => "1111111111000111",
61670 => "1111111111000111",
61671 => "1111111111000111",
61672 => "1111111111000111",
61673 => "1111111111000111",
61674 => "1111111111000111",
61675 => "1111111111000111",
61676 => "1111111111000111",
61677 => "1111111111000111",
61678 => "1111111111000111",
61679 => "1111111111000111",
61680 => "1111111111000111",
61681 => "1111111111000111",
61682 => "1111111111000111",
61683 => "1111111111000111",
61684 => "1111111111000111",
61685 => "1111111111000111",
61686 => "1111111111000111",
61687 => "1111111111000111",
61688 => "1111111111000111",
61689 => "1111111111000111",
61690 => "1111111111000111",
61691 => "1111111111000111",
61692 => "1111111111000111",
61693 => "1111111111000111",
61694 => "1111111111000111",
61695 => "1111111111000111",
61696 => "1111111111000111",
61697 => "1111111111000111",
61698 => "1111111111000111",
61699 => "1111111111000111",
61700 => "1111111111000111",
61701 => "1111111111000111",
61702 => "1111111111001000",
61703 => "1111111111001000",
61704 => "1111111111001000",
61705 => "1111111111001000",
61706 => "1111111111001000",
61707 => "1111111111001000",
61708 => "1111111111001000",
61709 => "1111111111001000",
61710 => "1111111111001000",
61711 => "1111111111001000",
61712 => "1111111111001000",
61713 => "1111111111001000",
61714 => "1111111111001000",
61715 => "1111111111001000",
61716 => "1111111111001000",
61717 => "1111111111001000",
61718 => "1111111111001000",
61719 => "1111111111001000",
61720 => "1111111111001000",
61721 => "1111111111001000",
61722 => "1111111111001000",
61723 => "1111111111001000",
61724 => "1111111111001000",
61725 => "1111111111001000",
61726 => "1111111111001000",
61727 => "1111111111001000",
61728 => "1111111111001000",
61729 => "1111111111001000",
61730 => "1111111111001000",
61731 => "1111111111001000",
61732 => "1111111111001000",
61733 => "1111111111001000",
61734 => "1111111111001000",
61735 => "1111111111001000",
61736 => "1111111111001000",
61737 => "1111111111001000",
61738 => "1111111111001000",
61739 => "1111111111001000",
61740 => "1111111111001000",
61741 => "1111111111001000",
61742 => "1111111111001000",
61743 => "1111111111001000",
61744 => "1111111111001000",
61745 => "1111111111001000",
61746 => "1111111111001000",
61747 => "1111111111001000",
61748 => "1111111111001000",
61749 => "1111111111001000",
61750 => "1111111111001000",
61751 => "1111111111001000",
61752 => "1111111111001000",
61753 => "1111111111001000",
61754 => "1111111111001000",
61755 => "1111111111001000",
61756 => "1111111111001000",
61757 => "1111111111001000",
61758 => "1111111111001000",
61759 => "1111111111001000",
61760 => "1111111111001000",
61761 => "1111111111001000",
61762 => "1111111111001000",
61763 => "1111111111001000",
61764 => "1111111111001000",
61765 => "1111111111001000",
61766 => "1111111111001000",
61767 => "1111111111001000",
61768 => "1111111111001000",
61769 => "1111111111001000",
61770 => "1111111111001000",
61771 => "1111111111001000",
61772 => "1111111111001000",
61773 => "1111111111001000",
61774 => "1111111111001000",
61775 => "1111111111001000",
61776 => "1111111111001001",
61777 => "1111111111001001",
61778 => "1111111111001001",
61779 => "1111111111001001",
61780 => "1111111111001001",
61781 => "1111111111001001",
61782 => "1111111111001001",
61783 => "1111111111001001",
61784 => "1111111111001001",
61785 => "1111111111001001",
61786 => "1111111111001001",
61787 => "1111111111001001",
61788 => "1111111111001001",
61789 => "1111111111001001",
61790 => "1111111111001001",
61791 => "1111111111001001",
61792 => "1111111111001001",
61793 => "1111111111001001",
61794 => "1111111111001001",
61795 => "1111111111001001",
61796 => "1111111111001001",
61797 => "1111111111001001",
61798 => "1111111111001001",
61799 => "1111111111001001",
61800 => "1111111111001001",
61801 => "1111111111001001",
61802 => "1111111111001001",
61803 => "1111111111001001",
61804 => "1111111111001001",
61805 => "1111111111001001",
61806 => "1111111111001001",
61807 => "1111111111001001",
61808 => "1111111111001001",
61809 => "1111111111001001",
61810 => "1111111111001001",
61811 => "1111111111001001",
61812 => "1111111111001001",
61813 => "1111111111001001",
61814 => "1111111111001001",
61815 => "1111111111001001",
61816 => "1111111111001001",
61817 => "1111111111001001",
61818 => "1111111111001001",
61819 => "1111111111001001",
61820 => "1111111111001001",
61821 => "1111111111001001",
61822 => "1111111111001001",
61823 => "1111111111001001",
61824 => "1111111111001001",
61825 => "1111111111001001",
61826 => "1111111111001001",
61827 => "1111111111001001",
61828 => "1111111111001001",
61829 => "1111111111001001",
61830 => "1111111111001001",
61831 => "1111111111001001",
61832 => "1111111111001001",
61833 => "1111111111001001",
61834 => "1111111111001001",
61835 => "1111111111001001",
61836 => "1111111111001001",
61837 => "1111111111001001",
61838 => "1111111111001001",
61839 => "1111111111001001",
61840 => "1111111111001001",
61841 => "1111111111001001",
61842 => "1111111111001001",
61843 => "1111111111001001",
61844 => "1111111111001001",
61845 => "1111111111001001",
61846 => "1111111111001001",
61847 => "1111111111001001",
61848 => "1111111111001001",
61849 => "1111111111001001",
61850 => "1111111111001001",
61851 => "1111111111001010",
61852 => "1111111111001010",
61853 => "1111111111001010",
61854 => "1111111111001010",
61855 => "1111111111001010",
61856 => "1111111111001010",
61857 => "1111111111001010",
61858 => "1111111111001010",
61859 => "1111111111001010",
61860 => "1111111111001010",
61861 => "1111111111001010",
61862 => "1111111111001010",
61863 => "1111111111001010",
61864 => "1111111111001010",
61865 => "1111111111001010",
61866 => "1111111111001010",
61867 => "1111111111001010",
61868 => "1111111111001010",
61869 => "1111111111001010",
61870 => "1111111111001010",
61871 => "1111111111001010",
61872 => "1111111111001010",
61873 => "1111111111001010",
61874 => "1111111111001010",
61875 => "1111111111001010",
61876 => "1111111111001010",
61877 => "1111111111001010",
61878 => "1111111111001010",
61879 => "1111111111001010",
61880 => "1111111111001010",
61881 => "1111111111001010",
61882 => "1111111111001010",
61883 => "1111111111001010",
61884 => "1111111111001010",
61885 => "1111111111001010",
61886 => "1111111111001010",
61887 => "1111111111001010",
61888 => "1111111111001010",
61889 => "1111111111001010",
61890 => "1111111111001010",
61891 => "1111111111001010",
61892 => "1111111111001010",
61893 => "1111111111001010",
61894 => "1111111111001010",
61895 => "1111111111001010",
61896 => "1111111111001010",
61897 => "1111111111001010",
61898 => "1111111111001010",
61899 => "1111111111001010",
61900 => "1111111111001010",
61901 => "1111111111001010",
61902 => "1111111111001010",
61903 => "1111111111001010",
61904 => "1111111111001010",
61905 => "1111111111001010",
61906 => "1111111111001010",
61907 => "1111111111001010",
61908 => "1111111111001010",
61909 => "1111111111001010",
61910 => "1111111111001010",
61911 => "1111111111001010",
61912 => "1111111111001010",
61913 => "1111111111001010",
61914 => "1111111111001010",
61915 => "1111111111001010",
61916 => "1111111111001010",
61917 => "1111111111001010",
61918 => "1111111111001010",
61919 => "1111111111001010",
61920 => "1111111111001010",
61921 => "1111111111001010",
61922 => "1111111111001010",
61923 => "1111111111001010",
61924 => "1111111111001010",
61925 => "1111111111001010",
61926 => "1111111111001010",
61927 => "1111111111001010",
61928 => "1111111111001011",
61929 => "1111111111001011",
61930 => "1111111111001011",
61931 => "1111111111001011",
61932 => "1111111111001011",
61933 => "1111111111001011",
61934 => "1111111111001011",
61935 => "1111111111001011",
61936 => "1111111111001011",
61937 => "1111111111001011",
61938 => "1111111111001011",
61939 => "1111111111001011",
61940 => "1111111111001011",
61941 => "1111111111001011",
61942 => "1111111111001011",
61943 => "1111111111001011",
61944 => "1111111111001011",
61945 => "1111111111001011",
61946 => "1111111111001011",
61947 => "1111111111001011",
61948 => "1111111111001011",
61949 => "1111111111001011",
61950 => "1111111111001011",
61951 => "1111111111001011",
61952 => "1111111111001011",
61953 => "1111111111001011",
61954 => "1111111111001011",
61955 => "1111111111001011",
61956 => "1111111111001011",
61957 => "1111111111001011",
61958 => "1111111111001011",
61959 => "1111111111001011",
61960 => "1111111111001011",
61961 => "1111111111001011",
61962 => "1111111111001011",
61963 => "1111111111001011",
61964 => "1111111111001011",
61965 => "1111111111001011",
61966 => "1111111111001011",
61967 => "1111111111001011",
61968 => "1111111111001011",
61969 => "1111111111001011",
61970 => "1111111111001011",
61971 => "1111111111001011",
61972 => "1111111111001011",
61973 => "1111111111001011",
61974 => "1111111111001011",
61975 => "1111111111001011",
61976 => "1111111111001011",
61977 => "1111111111001011",
61978 => "1111111111001011",
61979 => "1111111111001011",
61980 => "1111111111001011",
61981 => "1111111111001011",
61982 => "1111111111001011",
61983 => "1111111111001011",
61984 => "1111111111001011",
61985 => "1111111111001011",
61986 => "1111111111001011",
61987 => "1111111111001011",
61988 => "1111111111001011",
61989 => "1111111111001011",
61990 => "1111111111001011",
61991 => "1111111111001011",
61992 => "1111111111001011",
61993 => "1111111111001011",
61994 => "1111111111001011",
61995 => "1111111111001011",
61996 => "1111111111001011",
61997 => "1111111111001011",
61998 => "1111111111001011",
61999 => "1111111111001011",
62000 => "1111111111001011",
62001 => "1111111111001011",
62002 => "1111111111001011",
62003 => "1111111111001011",
62004 => "1111111111001011",
62005 => "1111111111001011",
62006 => "1111111111001100",
62007 => "1111111111001100",
62008 => "1111111111001100",
62009 => "1111111111001100",
62010 => "1111111111001100",
62011 => "1111111111001100",
62012 => "1111111111001100",
62013 => "1111111111001100",
62014 => "1111111111001100",
62015 => "1111111111001100",
62016 => "1111111111001100",
62017 => "1111111111001100",
62018 => "1111111111001100",
62019 => "1111111111001100",
62020 => "1111111111001100",
62021 => "1111111111001100",
62022 => "1111111111001100",
62023 => "1111111111001100",
62024 => "1111111111001100",
62025 => "1111111111001100",
62026 => "1111111111001100",
62027 => "1111111111001100",
62028 => "1111111111001100",
62029 => "1111111111001100",
62030 => "1111111111001100",
62031 => "1111111111001100",
62032 => "1111111111001100",
62033 => "1111111111001100",
62034 => "1111111111001100",
62035 => "1111111111001100",
62036 => "1111111111001100",
62037 => "1111111111001100",
62038 => "1111111111001100",
62039 => "1111111111001100",
62040 => "1111111111001100",
62041 => "1111111111001100",
62042 => "1111111111001100",
62043 => "1111111111001100",
62044 => "1111111111001100",
62045 => "1111111111001100",
62046 => "1111111111001100",
62047 => "1111111111001100",
62048 => "1111111111001100",
62049 => "1111111111001100",
62050 => "1111111111001100",
62051 => "1111111111001100",
62052 => "1111111111001100",
62053 => "1111111111001100",
62054 => "1111111111001100",
62055 => "1111111111001100",
62056 => "1111111111001100",
62057 => "1111111111001100",
62058 => "1111111111001100",
62059 => "1111111111001100",
62060 => "1111111111001100",
62061 => "1111111111001100",
62062 => "1111111111001100",
62063 => "1111111111001100",
62064 => "1111111111001100",
62065 => "1111111111001100",
62066 => "1111111111001100",
62067 => "1111111111001100",
62068 => "1111111111001100",
62069 => "1111111111001100",
62070 => "1111111111001100",
62071 => "1111111111001100",
62072 => "1111111111001100",
62073 => "1111111111001100",
62074 => "1111111111001100",
62075 => "1111111111001100",
62076 => "1111111111001100",
62077 => "1111111111001100",
62078 => "1111111111001100",
62079 => "1111111111001100",
62080 => "1111111111001100",
62081 => "1111111111001100",
62082 => "1111111111001100",
62083 => "1111111111001100",
62084 => "1111111111001100",
62085 => "1111111111001100",
62086 => "1111111111001101",
62087 => "1111111111001101",
62088 => "1111111111001101",
62089 => "1111111111001101",
62090 => "1111111111001101",
62091 => "1111111111001101",
62092 => "1111111111001101",
62093 => "1111111111001101",
62094 => "1111111111001101",
62095 => "1111111111001101",
62096 => "1111111111001101",
62097 => "1111111111001101",
62098 => "1111111111001101",
62099 => "1111111111001101",
62100 => "1111111111001101",
62101 => "1111111111001101",
62102 => "1111111111001101",
62103 => "1111111111001101",
62104 => "1111111111001101",
62105 => "1111111111001101",
62106 => "1111111111001101",
62107 => "1111111111001101",
62108 => "1111111111001101",
62109 => "1111111111001101",
62110 => "1111111111001101",
62111 => "1111111111001101",
62112 => "1111111111001101",
62113 => "1111111111001101",
62114 => "1111111111001101",
62115 => "1111111111001101",
62116 => "1111111111001101",
62117 => "1111111111001101",
62118 => "1111111111001101",
62119 => "1111111111001101",
62120 => "1111111111001101",
62121 => "1111111111001101",
62122 => "1111111111001101",
62123 => "1111111111001101",
62124 => "1111111111001101",
62125 => "1111111111001101",
62126 => "1111111111001101",
62127 => "1111111111001101",
62128 => "1111111111001101",
62129 => "1111111111001101",
62130 => "1111111111001101",
62131 => "1111111111001101",
62132 => "1111111111001101",
62133 => "1111111111001101",
62134 => "1111111111001101",
62135 => "1111111111001101",
62136 => "1111111111001101",
62137 => "1111111111001101",
62138 => "1111111111001101",
62139 => "1111111111001101",
62140 => "1111111111001101",
62141 => "1111111111001101",
62142 => "1111111111001101",
62143 => "1111111111001101",
62144 => "1111111111001101",
62145 => "1111111111001101",
62146 => "1111111111001101",
62147 => "1111111111001101",
62148 => "1111111111001101",
62149 => "1111111111001101",
62150 => "1111111111001101",
62151 => "1111111111001101",
62152 => "1111111111001101",
62153 => "1111111111001101",
62154 => "1111111111001101",
62155 => "1111111111001101",
62156 => "1111111111001101",
62157 => "1111111111001101",
62158 => "1111111111001101",
62159 => "1111111111001101",
62160 => "1111111111001101",
62161 => "1111111111001101",
62162 => "1111111111001101",
62163 => "1111111111001101",
62164 => "1111111111001101",
62165 => "1111111111001101",
62166 => "1111111111001101",
62167 => "1111111111001110",
62168 => "1111111111001110",
62169 => "1111111111001110",
62170 => "1111111111001110",
62171 => "1111111111001110",
62172 => "1111111111001110",
62173 => "1111111111001110",
62174 => "1111111111001110",
62175 => "1111111111001110",
62176 => "1111111111001110",
62177 => "1111111111001110",
62178 => "1111111111001110",
62179 => "1111111111001110",
62180 => "1111111111001110",
62181 => "1111111111001110",
62182 => "1111111111001110",
62183 => "1111111111001110",
62184 => "1111111111001110",
62185 => "1111111111001110",
62186 => "1111111111001110",
62187 => "1111111111001110",
62188 => "1111111111001110",
62189 => "1111111111001110",
62190 => "1111111111001110",
62191 => "1111111111001110",
62192 => "1111111111001110",
62193 => "1111111111001110",
62194 => "1111111111001110",
62195 => "1111111111001110",
62196 => "1111111111001110",
62197 => "1111111111001110",
62198 => "1111111111001110",
62199 => "1111111111001110",
62200 => "1111111111001110",
62201 => "1111111111001110",
62202 => "1111111111001110",
62203 => "1111111111001110",
62204 => "1111111111001110",
62205 => "1111111111001110",
62206 => "1111111111001110",
62207 => "1111111111001110",
62208 => "1111111111001110",
62209 => "1111111111001110",
62210 => "1111111111001110",
62211 => "1111111111001110",
62212 => "1111111111001110",
62213 => "1111111111001110",
62214 => "1111111111001110",
62215 => "1111111111001110",
62216 => "1111111111001110",
62217 => "1111111111001110",
62218 => "1111111111001110",
62219 => "1111111111001110",
62220 => "1111111111001110",
62221 => "1111111111001110",
62222 => "1111111111001110",
62223 => "1111111111001110",
62224 => "1111111111001110",
62225 => "1111111111001110",
62226 => "1111111111001110",
62227 => "1111111111001110",
62228 => "1111111111001110",
62229 => "1111111111001110",
62230 => "1111111111001110",
62231 => "1111111111001110",
62232 => "1111111111001110",
62233 => "1111111111001110",
62234 => "1111111111001110",
62235 => "1111111111001110",
62236 => "1111111111001110",
62237 => "1111111111001110",
62238 => "1111111111001110",
62239 => "1111111111001110",
62240 => "1111111111001110",
62241 => "1111111111001110",
62242 => "1111111111001110",
62243 => "1111111111001110",
62244 => "1111111111001110",
62245 => "1111111111001110",
62246 => "1111111111001110",
62247 => "1111111111001110",
62248 => "1111111111001110",
62249 => "1111111111001110",
62250 => "1111111111001111",
62251 => "1111111111001111",
62252 => "1111111111001111",
62253 => "1111111111001111",
62254 => "1111111111001111",
62255 => "1111111111001111",
62256 => "1111111111001111",
62257 => "1111111111001111",
62258 => "1111111111001111",
62259 => "1111111111001111",
62260 => "1111111111001111",
62261 => "1111111111001111",
62262 => "1111111111001111",
62263 => "1111111111001111",
62264 => "1111111111001111",
62265 => "1111111111001111",
62266 => "1111111111001111",
62267 => "1111111111001111",
62268 => "1111111111001111",
62269 => "1111111111001111",
62270 => "1111111111001111",
62271 => "1111111111001111",
62272 => "1111111111001111",
62273 => "1111111111001111",
62274 => "1111111111001111",
62275 => "1111111111001111",
62276 => "1111111111001111",
62277 => "1111111111001111",
62278 => "1111111111001111",
62279 => "1111111111001111",
62280 => "1111111111001111",
62281 => "1111111111001111",
62282 => "1111111111001111",
62283 => "1111111111001111",
62284 => "1111111111001111",
62285 => "1111111111001111",
62286 => "1111111111001111",
62287 => "1111111111001111",
62288 => "1111111111001111",
62289 => "1111111111001111",
62290 => "1111111111001111",
62291 => "1111111111001111",
62292 => "1111111111001111",
62293 => "1111111111001111",
62294 => "1111111111001111",
62295 => "1111111111001111",
62296 => "1111111111001111",
62297 => "1111111111001111",
62298 => "1111111111001111",
62299 => "1111111111001111",
62300 => "1111111111001111",
62301 => "1111111111001111",
62302 => "1111111111001111",
62303 => "1111111111001111",
62304 => "1111111111001111",
62305 => "1111111111001111",
62306 => "1111111111001111",
62307 => "1111111111001111",
62308 => "1111111111001111",
62309 => "1111111111001111",
62310 => "1111111111001111",
62311 => "1111111111001111",
62312 => "1111111111001111",
62313 => "1111111111001111",
62314 => "1111111111001111",
62315 => "1111111111001111",
62316 => "1111111111001111",
62317 => "1111111111001111",
62318 => "1111111111001111",
62319 => "1111111111001111",
62320 => "1111111111001111",
62321 => "1111111111001111",
62322 => "1111111111001111",
62323 => "1111111111001111",
62324 => "1111111111001111",
62325 => "1111111111001111",
62326 => "1111111111001111",
62327 => "1111111111001111",
62328 => "1111111111001111",
62329 => "1111111111001111",
62330 => "1111111111001111",
62331 => "1111111111001111",
62332 => "1111111111001111",
62333 => "1111111111001111",
62334 => "1111111111010000",
62335 => "1111111111010000",
62336 => "1111111111010000",
62337 => "1111111111010000",
62338 => "1111111111010000",
62339 => "1111111111010000",
62340 => "1111111111010000",
62341 => "1111111111010000",
62342 => "1111111111010000",
62343 => "1111111111010000",
62344 => "1111111111010000",
62345 => "1111111111010000",
62346 => "1111111111010000",
62347 => "1111111111010000",
62348 => "1111111111010000",
62349 => "1111111111010000",
62350 => "1111111111010000",
62351 => "1111111111010000",
62352 => "1111111111010000",
62353 => "1111111111010000",
62354 => "1111111111010000",
62355 => "1111111111010000",
62356 => "1111111111010000",
62357 => "1111111111010000",
62358 => "1111111111010000",
62359 => "1111111111010000",
62360 => "1111111111010000",
62361 => "1111111111010000",
62362 => "1111111111010000",
62363 => "1111111111010000",
62364 => "1111111111010000",
62365 => "1111111111010000",
62366 => "1111111111010000",
62367 => "1111111111010000",
62368 => "1111111111010000",
62369 => "1111111111010000",
62370 => "1111111111010000",
62371 => "1111111111010000",
62372 => "1111111111010000",
62373 => "1111111111010000",
62374 => "1111111111010000",
62375 => "1111111111010000",
62376 => "1111111111010000",
62377 => "1111111111010000",
62378 => "1111111111010000",
62379 => "1111111111010000",
62380 => "1111111111010000",
62381 => "1111111111010000",
62382 => "1111111111010000",
62383 => "1111111111010000",
62384 => "1111111111010000",
62385 => "1111111111010000",
62386 => "1111111111010000",
62387 => "1111111111010000",
62388 => "1111111111010000",
62389 => "1111111111010000",
62390 => "1111111111010000",
62391 => "1111111111010000",
62392 => "1111111111010000",
62393 => "1111111111010000",
62394 => "1111111111010000",
62395 => "1111111111010000",
62396 => "1111111111010000",
62397 => "1111111111010000",
62398 => "1111111111010000",
62399 => "1111111111010000",
62400 => "1111111111010000",
62401 => "1111111111010000",
62402 => "1111111111010000",
62403 => "1111111111010000",
62404 => "1111111111010000",
62405 => "1111111111010000",
62406 => "1111111111010000",
62407 => "1111111111010000",
62408 => "1111111111010000",
62409 => "1111111111010000",
62410 => "1111111111010000",
62411 => "1111111111010000",
62412 => "1111111111010000",
62413 => "1111111111010000",
62414 => "1111111111010000",
62415 => "1111111111010000",
62416 => "1111111111010000",
62417 => "1111111111010000",
62418 => "1111111111010000",
62419 => "1111111111010000",
62420 => "1111111111010001",
62421 => "1111111111010001",
62422 => "1111111111010001",
62423 => "1111111111010001",
62424 => "1111111111010001",
62425 => "1111111111010001",
62426 => "1111111111010001",
62427 => "1111111111010001",
62428 => "1111111111010001",
62429 => "1111111111010001",
62430 => "1111111111010001",
62431 => "1111111111010001",
62432 => "1111111111010001",
62433 => "1111111111010001",
62434 => "1111111111010001",
62435 => "1111111111010001",
62436 => "1111111111010001",
62437 => "1111111111010001",
62438 => "1111111111010001",
62439 => "1111111111010001",
62440 => "1111111111010001",
62441 => "1111111111010001",
62442 => "1111111111010001",
62443 => "1111111111010001",
62444 => "1111111111010001",
62445 => "1111111111010001",
62446 => "1111111111010001",
62447 => "1111111111010001",
62448 => "1111111111010001",
62449 => "1111111111010001",
62450 => "1111111111010001",
62451 => "1111111111010001",
62452 => "1111111111010001",
62453 => "1111111111010001",
62454 => "1111111111010001",
62455 => "1111111111010001",
62456 => "1111111111010001",
62457 => "1111111111010001",
62458 => "1111111111010001",
62459 => "1111111111010001",
62460 => "1111111111010001",
62461 => "1111111111010001",
62462 => "1111111111010001",
62463 => "1111111111010001",
62464 => "1111111111010001",
62465 => "1111111111010001",
62466 => "1111111111010001",
62467 => "1111111111010001",
62468 => "1111111111010001",
62469 => "1111111111010001",
62470 => "1111111111010001",
62471 => "1111111111010001",
62472 => "1111111111010001",
62473 => "1111111111010001",
62474 => "1111111111010001",
62475 => "1111111111010001",
62476 => "1111111111010001",
62477 => "1111111111010001",
62478 => "1111111111010001",
62479 => "1111111111010001",
62480 => "1111111111010001",
62481 => "1111111111010001",
62482 => "1111111111010001",
62483 => "1111111111010001",
62484 => "1111111111010001",
62485 => "1111111111010001",
62486 => "1111111111010001",
62487 => "1111111111010001",
62488 => "1111111111010001",
62489 => "1111111111010001",
62490 => "1111111111010001",
62491 => "1111111111010001",
62492 => "1111111111010001",
62493 => "1111111111010001",
62494 => "1111111111010001",
62495 => "1111111111010001",
62496 => "1111111111010001",
62497 => "1111111111010001",
62498 => "1111111111010001",
62499 => "1111111111010001",
62500 => "1111111111010001",
62501 => "1111111111010001",
62502 => "1111111111010001",
62503 => "1111111111010001",
62504 => "1111111111010001",
62505 => "1111111111010001",
62506 => "1111111111010001",
62507 => "1111111111010001",
62508 => "1111111111010001",
62509 => "1111111111010010",
62510 => "1111111111010010",
62511 => "1111111111010010",
62512 => "1111111111010010",
62513 => "1111111111010010",
62514 => "1111111111010010",
62515 => "1111111111010010",
62516 => "1111111111010010",
62517 => "1111111111010010",
62518 => "1111111111010010",
62519 => "1111111111010010",
62520 => "1111111111010010",
62521 => "1111111111010010",
62522 => "1111111111010010",
62523 => "1111111111010010",
62524 => "1111111111010010",
62525 => "1111111111010010",
62526 => "1111111111010010",
62527 => "1111111111010010",
62528 => "1111111111010010",
62529 => "1111111111010010",
62530 => "1111111111010010",
62531 => "1111111111010010",
62532 => "1111111111010010",
62533 => "1111111111010010",
62534 => "1111111111010010",
62535 => "1111111111010010",
62536 => "1111111111010010",
62537 => "1111111111010010",
62538 => "1111111111010010",
62539 => "1111111111010010",
62540 => "1111111111010010",
62541 => "1111111111010010",
62542 => "1111111111010010",
62543 => "1111111111010010",
62544 => "1111111111010010",
62545 => "1111111111010010",
62546 => "1111111111010010",
62547 => "1111111111010010",
62548 => "1111111111010010",
62549 => "1111111111010010",
62550 => "1111111111010010",
62551 => "1111111111010010",
62552 => "1111111111010010",
62553 => "1111111111010010",
62554 => "1111111111010010",
62555 => "1111111111010010",
62556 => "1111111111010010",
62557 => "1111111111010010",
62558 => "1111111111010010",
62559 => "1111111111010010",
62560 => "1111111111010010",
62561 => "1111111111010010",
62562 => "1111111111010010",
62563 => "1111111111010010",
62564 => "1111111111010010",
62565 => "1111111111010010",
62566 => "1111111111010010",
62567 => "1111111111010010",
62568 => "1111111111010010",
62569 => "1111111111010010",
62570 => "1111111111010010",
62571 => "1111111111010010",
62572 => "1111111111010010",
62573 => "1111111111010010",
62574 => "1111111111010010",
62575 => "1111111111010010",
62576 => "1111111111010010",
62577 => "1111111111010010",
62578 => "1111111111010010",
62579 => "1111111111010010",
62580 => "1111111111010010",
62581 => "1111111111010010",
62582 => "1111111111010010",
62583 => "1111111111010010",
62584 => "1111111111010010",
62585 => "1111111111010010",
62586 => "1111111111010010",
62587 => "1111111111010010",
62588 => "1111111111010010",
62589 => "1111111111010010",
62590 => "1111111111010010",
62591 => "1111111111010010",
62592 => "1111111111010010",
62593 => "1111111111010010",
62594 => "1111111111010010",
62595 => "1111111111010010",
62596 => "1111111111010010",
62597 => "1111111111010010",
62598 => "1111111111010010",
62599 => "1111111111010011",
62600 => "1111111111010011",
62601 => "1111111111010011",
62602 => "1111111111010011",
62603 => "1111111111010011",
62604 => "1111111111010011",
62605 => "1111111111010011",
62606 => "1111111111010011",
62607 => "1111111111010011",
62608 => "1111111111010011",
62609 => "1111111111010011",
62610 => "1111111111010011",
62611 => "1111111111010011",
62612 => "1111111111010011",
62613 => "1111111111010011",
62614 => "1111111111010011",
62615 => "1111111111010011",
62616 => "1111111111010011",
62617 => "1111111111010011",
62618 => "1111111111010011",
62619 => "1111111111010011",
62620 => "1111111111010011",
62621 => "1111111111010011",
62622 => "1111111111010011",
62623 => "1111111111010011",
62624 => "1111111111010011",
62625 => "1111111111010011",
62626 => "1111111111010011",
62627 => "1111111111010011",
62628 => "1111111111010011",
62629 => "1111111111010011",
62630 => "1111111111010011",
62631 => "1111111111010011",
62632 => "1111111111010011",
62633 => "1111111111010011",
62634 => "1111111111010011",
62635 => "1111111111010011",
62636 => "1111111111010011",
62637 => "1111111111010011",
62638 => "1111111111010011",
62639 => "1111111111010011",
62640 => "1111111111010011",
62641 => "1111111111010011",
62642 => "1111111111010011",
62643 => "1111111111010011",
62644 => "1111111111010011",
62645 => "1111111111010011",
62646 => "1111111111010011",
62647 => "1111111111010011",
62648 => "1111111111010011",
62649 => "1111111111010011",
62650 => "1111111111010011",
62651 => "1111111111010011",
62652 => "1111111111010011",
62653 => "1111111111010011",
62654 => "1111111111010011",
62655 => "1111111111010011",
62656 => "1111111111010011",
62657 => "1111111111010011",
62658 => "1111111111010011",
62659 => "1111111111010011",
62660 => "1111111111010011",
62661 => "1111111111010011",
62662 => "1111111111010011",
62663 => "1111111111010011",
62664 => "1111111111010011",
62665 => "1111111111010011",
62666 => "1111111111010011",
62667 => "1111111111010011",
62668 => "1111111111010011",
62669 => "1111111111010011",
62670 => "1111111111010011",
62671 => "1111111111010011",
62672 => "1111111111010011",
62673 => "1111111111010011",
62674 => "1111111111010011",
62675 => "1111111111010011",
62676 => "1111111111010011",
62677 => "1111111111010011",
62678 => "1111111111010011",
62679 => "1111111111010011",
62680 => "1111111111010011",
62681 => "1111111111010011",
62682 => "1111111111010011",
62683 => "1111111111010011",
62684 => "1111111111010011",
62685 => "1111111111010011",
62686 => "1111111111010011",
62687 => "1111111111010011",
62688 => "1111111111010011",
62689 => "1111111111010011",
62690 => "1111111111010011",
62691 => "1111111111010100",
62692 => "1111111111010100",
62693 => "1111111111010100",
62694 => "1111111111010100",
62695 => "1111111111010100",
62696 => "1111111111010100",
62697 => "1111111111010100",
62698 => "1111111111010100",
62699 => "1111111111010100",
62700 => "1111111111010100",
62701 => "1111111111010100",
62702 => "1111111111010100",
62703 => "1111111111010100",
62704 => "1111111111010100",
62705 => "1111111111010100",
62706 => "1111111111010100",
62707 => "1111111111010100",
62708 => "1111111111010100",
62709 => "1111111111010100",
62710 => "1111111111010100",
62711 => "1111111111010100",
62712 => "1111111111010100",
62713 => "1111111111010100",
62714 => "1111111111010100",
62715 => "1111111111010100",
62716 => "1111111111010100",
62717 => "1111111111010100",
62718 => "1111111111010100",
62719 => "1111111111010100",
62720 => "1111111111010100",
62721 => "1111111111010100",
62722 => "1111111111010100",
62723 => "1111111111010100",
62724 => "1111111111010100",
62725 => "1111111111010100",
62726 => "1111111111010100",
62727 => "1111111111010100",
62728 => "1111111111010100",
62729 => "1111111111010100",
62730 => "1111111111010100",
62731 => "1111111111010100",
62732 => "1111111111010100",
62733 => "1111111111010100",
62734 => "1111111111010100",
62735 => "1111111111010100",
62736 => "1111111111010100",
62737 => "1111111111010100",
62738 => "1111111111010100",
62739 => "1111111111010100",
62740 => "1111111111010100",
62741 => "1111111111010100",
62742 => "1111111111010100",
62743 => "1111111111010100",
62744 => "1111111111010100",
62745 => "1111111111010100",
62746 => "1111111111010100",
62747 => "1111111111010100",
62748 => "1111111111010100",
62749 => "1111111111010100",
62750 => "1111111111010100",
62751 => "1111111111010100",
62752 => "1111111111010100",
62753 => "1111111111010100",
62754 => "1111111111010100",
62755 => "1111111111010100",
62756 => "1111111111010100",
62757 => "1111111111010100",
62758 => "1111111111010100",
62759 => "1111111111010100",
62760 => "1111111111010100",
62761 => "1111111111010100",
62762 => "1111111111010100",
62763 => "1111111111010100",
62764 => "1111111111010100",
62765 => "1111111111010100",
62766 => "1111111111010100",
62767 => "1111111111010100",
62768 => "1111111111010100",
62769 => "1111111111010100",
62770 => "1111111111010100",
62771 => "1111111111010100",
62772 => "1111111111010100",
62773 => "1111111111010100",
62774 => "1111111111010100",
62775 => "1111111111010100",
62776 => "1111111111010100",
62777 => "1111111111010100",
62778 => "1111111111010100",
62779 => "1111111111010100",
62780 => "1111111111010100",
62781 => "1111111111010100",
62782 => "1111111111010100",
62783 => "1111111111010100",
62784 => "1111111111010100",
62785 => "1111111111010101",
62786 => "1111111111010101",
62787 => "1111111111010101",
62788 => "1111111111010101",
62789 => "1111111111010101",
62790 => "1111111111010101",
62791 => "1111111111010101",
62792 => "1111111111010101",
62793 => "1111111111010101",
62794 => "1111111111010101",
62795 => "1111111111010101",
62796 => "1111111111010101",
62797 => "1111111111010101",
62798 => "1111111111010101",
62799 => "1111111111010101",
62800 => "1111111111010101",
62801 => "1111111111010101",
62802 => "1111111111010101",
62803 => "1111111111010101",
62804 => "1111111111010101",
62805 => "1111111111010101",
62806 => "1111111111010101",
62807 => "1111111111010101",
62808 => "1111111111010101",
62809 => "1111111111010101",
62810 => "1111111111010101",
62811 => "1111111111010101",
62812 => "1111111111010101",
62813 => "1111111111010101",
62814 => "1111111111010101",
62815 => "1111111111010101",
62816 => "1111111111010101",
62817 => "1111111111010101",
62818 => "1111111111010101",
62819 => "1111111111010101",
62820 => "1111111111010101",
62821 => "1111111111010101",
62822 => "1111111111010101",
62823 => "1111111111010101",
62824 => "1111111111010101",
62825 => "1111111111010101",
62826 => "1111111111010101",
62827 => "1111111111010101",
62828 => "1111111111010101",
62829 => "1111111111010101",
62830 => "1111111111010101",
62831 => "1111111111010101",
62832 => "1111111111010101",
62833 => "1111111111010101",
62834 => "1111111111010101",
62835 => "1111111111010101",
62836 => "1111111111010101",
62837 => "1111111111010101",
62838 => "1111111111010101",
62839 => "1111111111010101",
62840 => "1111111111010101",
62841 => "1111111111010101",
62842 => "1111111111010101",
62843 => "1111111111010101",
62844 => "1111111111010101",
62845 => "1111111111010101",
62846 => "1111111111010101",
62847 => "1111111111010101",
62848 => "1111111111010101",
62849 => "1111111111010101",
62850 => "1111111111010101",
62851 => "1111111111010101",
62852 => "1111111111010101",
62853 => "1111111111010101",
62854 => "1111111111010101",
62855 => "1111111111010101",
62856 => "1111111111010101",
62857 => "1111111111010101",
62858 => "1111111111010101",
62859 => "1111111111010101",
62860 => "1111111111010101",
62861 => "1111111111010101",
62862 => "1111111111010101",
62863 => "1111111111010101",
62864 => "1111111111010101",
62865 => "1111111111010101",
62866 => "1111111111010101",
62867 => "1111111111010101",
62868 => "1111111111010101",
62869 => "1111111111010101",
62870 => "1111111111010101",
62871 => "1111111111010101",
62872 => "1111111111010101",
62873 => "1111111111010101",
62874 => "1111111111010101",
62875 => "1111111111010101",
62876 => "1111111111010101",
62877 => "1111111111010101",
62878 => "1111111111010101",
62879 => "1111111111010101",
62880 => "1111111111010101",
62881 => "1111111111010101",
62882 => "1111111111010110",
62883 => "1111111111010110",
62884 => "1111111111010110",
62885 => "1111111111010110",
62886 => "1111111111010110",
62887 => "1111111111010110",
62888 => "1111111111010110",
62889 => "1111111111010110",
62890 => "1111111111010110",
62891 => "1111111111010110",
62892 => "1111111111010110",
62893 => "1111111111010110",
62894 => "1111111111010110",
62895 => "1111111111010110",
62896 => "1111111111010110",
62897 => "1111111111010110",
62898 => "1111111111010110",
62899 => "1111111111010110",
62900 => "1111111111010110",
62901 => "1111111111010110",
62902 => "1111111111010110",
62903 => "1111111111010110",
62904 => "1111111111010110",
62905 => "1111111111010110",
62906 => "1111111111010110",
62907 => "1111111111010110",
62908 => "1111111111010110",
62909 => "1111111111010110",
62910 => "1111111111010110",
62911 => "1111111111010110",
62912 => "1111111111010110",
62913 => "1111111111010110",
62914 => "1111111111010110",
62915 => "1111111111010110",
62916 => "1111111111010110",
62917 => "1111111111010110",
62918 => "1111111111010110",
62919 => "1111111111010110",
62920 => "1111111111010110",
62921 => "1111111111010110",
62922 => "1111111111010110",
62923 => "1111111111010110",
62924 => "1111111111010110",
62925 => "1111111111010110",
62926 => "1111111111010110",
62927 => "1111111111010110",
62928 => "1111111111010110",
62929 => "1111111111010110",
62930 => "1111111111010110",
62931 => "1111111111010110",
62932 => "1111111111010110",
62933 => "1111111111010110",
62934 => "1111111111010110",
62935 => "1111111111010110",
62936 => "1111111111010110",
62937 => "1111111111010110",
62938 => "1111111111010110",
62939 => "1111111111010110",
62940 => "1111111111010110",
62941 => "1111111111010110",
62942 => "1111111111010110",
62943 => "1111111111010110",
62944 => "1111111111010110",
62945 => "1111111111010110",
62946 => "1111111111010110",
62947 => "1111111111010110",
62948 => "1111111111010110",
62949 => "1111111111010110",
62950 => "1111111111010110",
62951 => "1111111111010110",
62952 => "1111111111010110",
62953 => "1111111111010110",
62954 => "1111111111010110",
62955 => "1111111111010110",
62956 => "1111111111010110",
62957 => "1111111111010110",
62958 => "1111111111010110",
62959 => "1111111111010110",
62960 => "1111111111010110",
62961 => "1111111111010110",
62962 => "1111111111010110",
62963 => "1111111111010110",
62964 => "1111111111010110",
62965 => "1111111111010110",
62966 => "1111111111010110",
62967 => "1111111111010110",
62968 => "1111111111010110",
62969 => "1111111111010110",
62970 => "1111111111010110",
62971 => "1111111111010110",
62972 => "1111111111010110",
62973 => "1111111111010110",
62974 => "1111111111010110",
62975 => "1111111111010110",
62976 => "1111111111010110",
62977 => "1111111111010110",
62978 => "1111111111010110",
62979 => "1111111111010110",
62980 => "1111111111010111",
62981 => "1111111111010111",
62982 => "1111111111010111",
62983 => "1111111111010111",
62984 => "1111111111010111",
62985 => "1111111111010111",
62986 => "1111111111010111",
62987 => "1111111111010111",
62988 => "1111111111010111",
62989 => "1111111111010111",
62990 => "1111111111010111",
62991 => "1111111111010111",
62992 => "1111111111010111",
62993 => "1111111111010111",
62994 => "1111111111010111",
62995 => "1111111111010111",
62996 => "1111111111010111",
62997 => "1111111111010111",
62998 => "1111111111010111",
62999 => "1111111111010111",
63000 => "1111111111010111",
63001 => "1111111111010111",
63002 => "1111111111010111",
63003 => "1111111111010111",
63004 => "1111111111010111",
63005 => "1111111111010111",
63006 => "1111111111010111",
63007 => "1111111111010111",
63008 => "1111111111010111",
63009 => "1111111111010111",
63010 => "1111111111010111",
63011 => "1111111111010111",
63012 => "1111111111010111",
63013 => "1111111111010111",
63014 => "1111111111010111",
63015 => "1111111111010111",
63016 => "1111111111010111",
63017 => "1111111111010111",
63018 => "1111111111010111",
63019 => "1111111111010111",
63020 => "1111111111010111",
63021 => "1111111111010111",
63022 => "1111111111010111",
63023 => "1111111111010111",
63024 => "1111111111010111",
63025 => "1111111111010111",
63026 => "1111111111010111",
63027 => "1111111111010111",
63028 => "1111111111010111",
63029 => "1111111111010111",
63030 => "1111111111010111",
63031 => "1111111111010111",
63032 => "1111111111010111",
63033 => "1111111111010111",
63034 => "1111111111010111",
63035 => "1111111111010111",
63036 => "1111111111010111",
63037 => "1111111111010111",
63038 => "1111111111010111",
63039 => "1111111111010111",
63040 => "1111111111010111",
63041 => "1111111111010111",
63042 => "1111111111010111",
63043 => "1111111111010111",
63044 => "1111111111010111",
63045 => "1111111111010111",
63046 => "1111111111010111",
63047 => "1111111111010111",
63048 => "1111111111010111",
63049 => "1111111111010111",
63050 => "1111111111010111",
63051 => "1111111111010111",
63052 => "1111111111010111",
63053 => "1111111111010111",
63054 => "1111111111010111",
63055 => "1111111111010111",
63056 => "1111111111010111",
63057 => "1111111111010111",
63058 => "1111111111010111",
63059 => "1111111111010111",
63060 => "1111111111010111",
63061 => "1111111111010111",
63062 => "1111111111010111",
63063 => "1111111111010111",
63064 => "1111111111010111",
63065 => "1111111111010111",
63066 => "1111111111010111",
63067 => "1111111111010111",
63068 => "1111111111010111",
63069 => "1111111111010111",
63070 => "1111111111010111",
63071 => "1111111111010111",
63072 => "1111111111010111",
63073 => "1111111111010111",
63074 => "1111111111010111",
63075 => "1111111111010111",
63076 => "1111111111010111",
63077 => "1111111111010111",
63078 => "1111111111010111",
63079 => "1111111111010111",
63080 => "1111111111010111",
63081 => "1111111111011000",
63082 => "1111111111011000",
63083 => "1111111111011000",
63084 => "1111111111011000",
63085 => "1111111111011000",
63086 => "1111111111011000",
63087 => "1111111111011000",
63088 => "1111111111011000",
63089 => "1111111111011000",
63090 => "1111111111011000",
63091 => "1111111111011000",
63092 => "1111111111011000",
63093 => "1111111111011000",
63094 => "1111111111011000",
63095 => "1111111111011000",
63096 => "1111111111011000",
63097 => "1111111111011000",
63098 => "1111111111011000",
63099 => "1111111111011000",
63100 => "1111111111011000",
63101 => "1111111111011000",
63102 => "1111111111011000",
63103 => "1111111111011000",
63104 => "1111111111011000",
63105 => "1111111111011000",
63106 => "1111111111011000",
63107 => "1111111111011000",
63108 => "1111111111011000",
63109 => "1111111111011000",
63110 => "1111111111011000",
63111 => "1111111111011000",
63112 => "1111111111011000",
63113 => "1111111111011000",
63114 => "1111111111011000",
63115 => "1111111111011000",
63116 => "1111111111011000",
63117 => "1111111111011000",
63118 => "1111111111011000",
63119 => "1111111111011000",
63120 => "1111111111011000",
63121 => "1111111111011000",
63122 => "1111111111011000",
63123 => "1111111111011000",
63124 => "1111111111011000",
63125 => "1111111111011000",
63126 => "1111111111011000",
63127 => "1111111111011000",
63128 => "1111111111011000",
63129 => "1111111111011000",
63130 => "1111111111011000",
63131 => "1111111111011000",
63132 => "1111111111011000",
63133 => "1111111111011000",
63134 => "1111111111011000",
63135 => "1111111111011000",
63136 => "1111111111011000",
63137 => "1111111111011000",
63138 => "1111111111011000",
63139 => "1111111111011000",
63140 => "1111111111011000",
63141 => "1111111111011000",
63142 => "1111111111011000",
63143 => "1111111111011000",
63144 => "1111111111011000",
63145 => "1111111111011000",
63146 => "1111111111011000",
63147 => "1111111111011000",
63148 => "1111111111011000",
63149 => "1111111111011000",
63150 => "1111111111011000",
63151 => "1111111111011000",
63152 => "1111111111011000",
63153 => "1111111111011000",
63154 => "1111111111011000",
63155 => "1111111111011000",
63156 => "1111111111011000",
63157 => "1111111111011000",
63158 => "1111111111011000",
63159 => "1111111111011000",
63160 => "1111111111011000",
63161 => "1111111111011000",
63162 => "1111111111011000",
63163 => "1111111111011000",
63164 => "1111111111011000",
63165 => "1111111111011000",
63166 => "1111111111011000",
63167 => "1111111111011000",
63168 => "1111111111011000",
63169 => "1111111111011000",
63170 => "1111111111011000",
63171 => "1111111111011000",
63172 => "1111111111011000",
63173 => "1111111111011000",
63174 => "1111111111011000",
63175 => "1111111111011000",
63176 => "1111111111011000",
63177 => "1111111111011000",
63178 => "1111111111011000",
63179 => "1111111111011000",
63180 => "1111111111011000",
63181 => "1111111111011000",
63182 => "1111111111011000",
63183 => "1111111111011000",
63184 => "1111111111011000",
63185 => "1111111111011001",
63186 => "1111111111011001",
63187 => "1111111111011001",
63188 => "1111111111011001",
63189 => "1111111111011001",
63190 => "1111111111011001",
63191 => "1111111111011001",
63192 => "1111111111011001",
63193 => "1111111111011001",
63194 => "1111111111011001",
63195 => "1111111111011001",
63196 => "1111111111011001",
63197 => "1111111111011001",
63198 => "1111111111011001",
63199 => "1111111111011001",
63200 => "1111111111011001",
63201 => "1111111111011001",
63202 => "1111111111011001",
63203 => "1111111111011001",
63204 => "1111111111011001",
63205 => "1111111111011001",
63206 => "1111111111011001",
63207 => "1111111111011001",
63208 => "1111111111011001",
63209 => "1111111111011001",
63210 => "1111111111011001",
63211 => "1111111111011001",
63212 => "1111111111011001",
63213 => "1111111111011001",
63214 => "1111111111011001",
63215 => "1111111111011001",
63216 => "1111111111011001",
63217 => "1111111111011001",
63218 => "1111111111011001",
63219 => "1111111111011001",
63220 => "1111111111011001",
63221 => "1111111111011001",
63222 => "1111111111011001",
63223 => "1111111111011001",
63224 => "1111111111011001",
63225 => "1111111111011001",
63226 => "1111111111011001",
63227 => "1111111111011001",
63228 => "1111111111011001",
63229 => "1111111111011001",
63230 => "1111111111011001",
63231 => "1111111111011001",
63232 => "1111111111011001",
63233 => "1111111111011001",
63234 => "1111111111011001",
63235 => "1111111111011001",
63236 => "1111111111011001",
63237 => "1111111111011001",
63238 => "1111111111011001",
63239 => "1111111111011001",
63240 => "1111111111011001",
63241 => "1111111111011001",
63242 => "1111111111011001",
63243 => "1111111111011001",
63244 => "1111111111011001",
63245 => "1111111111011001",
63246 => "1111111111011001",
63247 => "1111111111011001",
63248 => "1111111111011001",
63249 => "1111111111011001",
63250 => "1111111111011001",
63251 => "1111111111011001",
63252 => "1111111111011001",
63253 => "1111111111011001",
63254 => "1111111111011001",
63255 => "1111111111011001",
63256 => "1111111111011001",
63257 => "1111111111011001",
63258 => "1111111111011001",
63259 => "1111111111011001",
63260 => "1111111111011001",
63261 => "1111111111011001",
63262 => "1111111111011001",
63263 => "1111111111011001",
63264 => "1111111111011001",
63265 => "1111111111011001",
63266 => "1111111111011001",
63267 => "1111111111011001",
63268 => "1111111111011001",
63269 => "1111111111011001",
63270 => "1111111111011001",
63271 => "1111111111011001",
63272 => "1111111111011001",
63273 => "1111111111011001",
63274 => "1111111111011001",
63275 => "1111111111011001",
63276 => "1111111111011001",
63277 => "1111111111011001",
63278 => "1111111111011001",
63279 => "1111111111011001",
63280 => "1111111111011001",
63281 => "1111111111011001",
63282 => "1111111111011001",
63283 => "1111111111011001",
63284 => "1111111111011001",
63285 => "1111111111011001",
63286 => "1111111111011001",
63287 => "1111111111011001",
63288 => "1111111111011001",
63289 => "1111111111011001",
63290 => "1111111111011001",
63291 => "1111111111011001",
63292 => "1111111111011010",
63293 => "1111111111011010",
63294 => "1111111111011010",
63295 => "1111111111011010",
63296 => "1111111111011010",
63297 => "1111111111011010",
63298 => "1111111111011010",
63299 => "1111111111011010",
63300 => "1111111111011010",
63301 => "1111111111011010",
63302 => "1111111111011010",
63303 => "1111111111011010",
63304 => "1111111111011010",
63305 => "1111111111011010",
63306 => "1111111111011010",
63307 => "1111111111011010",
63308 => "1111111111011010",
63309 => "1111111111011010",
63310 => "1111111111011010",
63311 => "1111111111011010",
63312 => "1111111111011010",
63313 => "1111111111011010",
63314 => "1111111111011010",
63315 => "1111111111011010",
63316 => "1111111111011010",
63317 => "1111111111011010",
63318 => "1111111111011010",
63319 => "1111111111011010",
63320 => "1111111111011010",
63321 => "1111111111011010",
63322 => "1111111111011010",
63323 => "1111111111011010",
63324 => "1111111111011010",
63325 => "1111111111011010",
63326 => "1111111111011010",
63327 => "1111111111011010",
63328 => "1111111111011010",
63329 => "1111111111011010",
63330 => "1111111111011010",
63331 => "1111111111011010",
63332 => "1111111111011010",
63333 => "1111111111011010",
63334 => "1111111111011010",
63335 => "1111111111011010",
63336 => "1111111111011010",
63337 => "1111111111011010",
63338 => "1111111111011010",
63339 => "1111111111011010",
63340 => "1111111111011010",
63341 => "1111111111011010",
63342 => "1111111111011010",
63343 => "1111111111011010",
63344 => "1111111111011010",
63345 => "1111111111011010",
63346 => "1111111111011010",
63347 => "1111111111011010",
63348 => "1111111111011010",
63349 => "1111111111011010",
63350 => "1111111111011010",
63351 => "1111111111011010",
63352 => "1111111111011010",
63353 => "1111111111011010",
63354 => "1111111111011010",
63355 => "1111111111011010",
63356 => "1111111111011010",
63357 => "1111111111011010",
63358 => "1111111111011010",
63359 => "1111111111011010",
63360 => "1111111111011010",
63361 => "1111111111011010",
63362 => "1111111111011010",
63363 => "1111111111011010",
63364 => "1111111111011010",
63365 => "1111111111011010",
63366 => "1111111111011010",
63367 => "1111111111011010",
63368 => "1111111111011010",
63369 => "1111111111011010",
63370 => "1111111111011010",
63371 => "1111111111011010",
63372 => "1111111111011010",
63373 => "1111111111011010",
63374 => "1111111111011010",
63375 => "1111111111011010",
63376 => "1111111111011010",
63377 => "1111111111011010",
63378 => "1111111111011010",
63379 => "1111111111011010",
63380 => "1111111111011010",
63381 => "1111111111011010",
63382 => "1111111111011010",
63383 => "1111111111011010",
63384 => "1111111111011010",
63385 => "1111111111011010",
63386 => "1111111111011010",
63387 => "1111111111011010",
63388 => "1111111111011010",
63389 => "1111111111011010",
63390 => "1111111111011010",
63391 => "1111111111011010",
63392 => "1111111111011010",
63393 => "1111111111011010",
63394 => "1111111111011010",
63395 => "1111111111011010",
63396 => "1111111111011010",
63397 => "1111111111011010",
63398 => "1111111111011010",
63399 => "1111111111011010",
63400 => "1111111111011010",
63401 => "1111111111011011",
63402 => "1111111111011011",
63403 => "1111111111011011",
63404 => "1111111111011011",
63405 => "1111111111011011",
63406 => "1111111111011011",
63407 => "1111111111011011",
63408 => "1111111111011011",
63409 => "1111111111011011",
63410 => "1111111111011011",
63411 => "1111111111011011",
63412 => "1111111111011011",
63413 => "1111111111011011",
63414 => "1111111111011011",
63415 => "1111111111011011",
63416 => "1111111111011011",
63417 => "1111111111011011",
63418 => "1111111111011011",
63419 => "1111111111011011",
63420 => "1111111111011011",
63421 => "1111111111011011",
63422 => "1111111111011011",
63423 => "1111111111011011",
63424 => "1111111111011011",
63425 => "1111111111011011",
63426 => "1111111111011011",
63427 => "1111111111011011",
63428 => "1111111111011011",
63429 => "1111111111011011",
63430 => "1111111111011011",
63431 => "1111111111011011",
63432 => "1111111111011011",
63433 => "1111111111011011",
63434 => "1111111111011011",
63435 => "1111111111011011",
63436 => "1111111111011011",
63437 => "1111111111011011",
63438 => "1111111111011011",
63439 => "1111111111011011",
63440 => "1111111111011011",
63441 => "1111111111011011",
63442 => "1111111111011011",
63443 => "1111111111011011",
63444 => "1111111111011011",
63445 => "1111111111011011",
63446 => "1111111111011011",
63447 => "1111111111011011",
63448 => "1111111111011011",
63449 => "1111111111011011",
63450 => "1111111111011011",
63451 => "1111111111011011",
63452 => "1111111111011011",
63453 => "1111111111011011",
63454 => "1111111111011011",
63455 => "1111111111011011",
63456 => "1111111111011011",
63457 => "1111111111011011",
63458 => "1111111111011011",
63459 => "1111111111011011",
63460 => "1111111111011011",
63461 => "1111111111011011",
63462 => "1111111111011011",
63463 => "1111111111011011",
63464 => "1111111111011011",
63465 => "1111111111011011",
63466 => "1111111111011011",
63467 => "1111111111011011",
63468 => "1111111111011011",
63469 => "1111111111011011",
63470 => "1111111111011011",
63471 => "1111111111011011",
63472 => "1111111111011011",
63473 => "1111111111011011",
63474 => "1111111111011011",
63475 => "1111111111011011",
63476 => "1111111111011011",
63477 => "1111111111011011",
63478 => "1111111111011011",
63479 => "1111111111011011",
63480 => "1111111111011011",
63481 => "1111111111011011",
63482 => "1111111111011011",
63483 => "1111111111011011",
63484 => "1111111111011011",
63485 => "1111111111011011",
63486 => "1111111111011011",
63487 => "1111111111011011",
63488 => "1111111111011011",
63489 => "1111111111011011",
63490 => "1111111111011011",
63491 => "1111111111011011",
63492 => "1111111111011011",
63493 => "1111111111011011",
63494 => "1111111111011011",
63495 => "1111111111011011",
63496 => "1111111111011011",
63497 => "1111111111011011",
63498 => "1111111111011011",
63499 => "1111111111011011",
63500 => "1111111111011011",
63501 => "1111111111011011",
63502 => "1111111111011011",
63503 => "1111111111011011",
63504 => "1111111111011011",
63505 => "1111111111011011",
63506 => "1111111111011011",
63507 => "1111111111011011",
63508 => "1111111111011011",
63509 => "1111111111011011",
63510 => "1111111111011011",
63511 => "1111111111011011",
63512 => "1111111111011011",
63513 => "1111111111011100",
63514 => "1111111111011100",
63515 => "1111111111011100",
63516 => "1111111111011100",
63517 => "1111111111011100",
63518 => "1111111111011100",
63519 => "1111111111011100",
63520 => "1111111111011100",
63521 => "1111111111011100",
63522 => "1111111111011100",
63523 => "1111111111011100",
63524 => "1111111111011100",
63525 => "1111111111011100",
63526 => "1111111111011100",
63527 => "1111111111011100",
63528 => "1111111111011100",
63529 => "1111111111011100",
63530 => "1111111111011100",
63531 => "1111111111011100",
63532 => "1111111111011100",
63533 => "1111111111011100",
63534 => "1111111111011100",
63535 => "1111111111011100",
63536 => "1111111111011100",
63537 => "1111111111011100",
63538 => "1111111111011100",
63539 => "1111111111011100",
63540 => "1111111111011100",
63541 => "1111111111011100",
63542 => "1111111111011100",
63543 => "1111111111011100",
63544 => "1111111111011100",
63545 => "1111111111011100",
63546 => "1111111111011100",
63547 => "1111111111011100",
63548 => "1111111111011100",
63549 => "1111111111011100",
63550 => "1111111111011100",
63551 => "1111111111011100",
63552 => "1111111111011100",
63553 => "1111111111011100",
63554 => "1111111111011100",
63555 => "1111111111011100",
63556 => "1111111111011100",
63557 => "1111111111011100",
63558 => "1111111111011100",
63559 => "1111111111011100",
63560 => "1111111111011100",
63561 => "1111111111011100",
63562 => "1111111111011100",
63563 => "1111111111011100",
63564 => "1111111111011100",
63565 => "1111111111011100",
63566 => "1111111111011100",
63567 => "1111111111011100",
63568 => "1111111111011100",
63569 => "1111111111011100",
63570 => "1111111111011100",
63571 => "1111111111011100",
63572 => "1111111111011100",
63573 => "1111111111011100",
63574 => "1111111111011100",
63575 => "1111111111011100",
63576 => "1111111111011100",
63577 => "1111111111011100",
63578 => "1111111111011100",
63579 => "1111111111011100",
63580 => "1111111111011100",
63581 => "1111111111011100",
63582 => "1111111111011100",
63583 => "1111111111011100",
63584 => "1111111111011100",
63585 => "1111111111011100",
63586 => "1111111111011100",
63587 => "1111111111011100",
63588 => "1111111111011100",
63589 => "1111111111011100",
63590 => "1111111111011100",
63591 => "1111111111011100",
63592 => "1111111111011100",
63593 => "1111111111011100",
63594 => "1111111111011100",
63595 => "1111111111011100",
63596 => "1111111111011100",
63597 => "1111111111011100",
63598 => "1111111111011100",
63599 => "1111111111011100",
63600 => "1111111111011100",
63601 => "1111111111011100",
63602 => "1111111111011100",
63603 => "1111111111011100",
63604 => "1111111111011100",
63605 => "1111111111011100",
63606 => "1111111111011100",
63607 => "1111111111011100",
63608 => "1111111111011100",
63609 => "1111111111011100",
63610 => "1111111111011100",
63611 => "1111111111011100",
63612 => "1111111111011100",
63613 => "1111111111011100",
63614 => "1111111111011100",
63615 => "1111111111011100",
63616 => "1111111111011100",
63617 => "1111111111011100",
63618 => "1111111111011100",
63619 => "1111111111011100",
63620 => "1111111111011100",
63621 => "1111111111011100",
63622 => "1111111111011100",
63623 => "1111111111011100",
63624 => "1111111111011100",
63625 => "1111111111011100",
63626 => "1111111111011100",
63627 => "1111111111011100",
63628 => "1111111111011100",
63629 => "1111111111011101",
63630 => "1111111111011101",
63631 => "1111111111011101",
63632 => "1111111111011101",
63633 => "1111111111011101",
63634 => "1111111111011101",
63635 => "1111111111011101",
63636 => "1111111111011101",
63637 => "1111111111011101",
63638 => "1111111111011101",
63639 => "1111111111011101",
63640 => "1111111111011101",
63641 => "1111111111011101",
63642 => "1111111111011101",
63643 => "1111111111011101",
63644 => "1111111111011101",
63645 => "1111111111011101",
63646 => "1111111111011101",
63647 => "1111111111011101",
63648 => "1111111111011101",
63649 => "1111111111011101",
63650 => "1111111111011101",
63651 => "1111111111011101",
63652 => "1111111111011101",
63653 => "1111111111011101",
63654 => "1111111111011101",
63655 => "1111111111011101",
63656 => "1111111111011101",
63657 => "1111111111011101",
63658 => "1111111111011101",
63659 => "1111111111011101",
63660 => "1111111111011101",
63661 => "1111111111011101",
63662 => "1111111111011101",
63663 => "1111111111011101",
63664 => "1111111111011101",
63665 => "1111111111011101",
63666 => "1111111111011101",
63667 => "1111111111011101",
63668 => "1111111111011101",
63669 => "1111111111011101",
63670 => "1111111111011101",
63671 => "1111111111011101",
63672 => "1111111111011101",
63673 => "1111111111011101",
63674 => "1111111111011101",
63675 => "1111111111011101",
63676 => "1111111111011101",
63677 => "1111111111011101",
63678 => "1111111111011101",
63679 => "1111111111011101",
63680 => "1111111111011101",
63681 => "1111111111011101",
63682 => "1111111111011101",
63683 => "1111111111011101",
63684 => "1111111111011101",
63685 => "1111111111011101",
63686 => "1111111111011101",
63687 => "1111111111011101",
63688 => "1111111111011101",
63689 => "1111111111011101",
63690 => "1111111111011101",
63691 => "1111111111011101",
63692 => "1111111111011101",
63693 => "1111111111011101",
63694 => "1111111111011101",
63695 => "1111111111011101",
63696 => "1111111111011101",
63697 => "1111111111011101",
63698 => "1111111111011101",
63699 => "1111111111011101",
63700 => "1111111111011101",
63701 => "1111111111011101",
63702 => "1111111111011101",
63703 => "1111111111011101",
63704 => "1111111111011101",
63705 => "1111111111011101",
63706 => "1111111111011101",
63707 => "1111111111011101",
63708 => "1111111111011101",
63709 => "1111111111011101",
63710 => "1111111111011101",
63711 => "1111111111011101",
63712 => "1111111111011101",
63713 => "1111111111011101",
63714 => "1111111111011101",
63715 => "1111111111011101",
63716 => "1111111111011101",
63717 => "1111111111011101",
63718 => "1111111111011101",
63719 => "1111111111011101",
63720 => "1111111111011101",
63721 => "1111111111011101",
63722 => "1111111111011101",
63723 => "1111111111011101",
63724 => "1111111111011101",
63725 => "1111111111011101",
63726 => "1111111111011101",
63727 => "1111111111011101",
63728 => "1111111111011101",
63729 => "1111111111011101",
63730 => "1111111111011101",
63731 => "1111111111011101",
63732 => "1111111111011101",
63733 => "1111111111011101",
63734 => "1111111111011101",
63735 => "1111111111011101",
63736 => "1111111111011101",
63737 => "1111111111011101",
63738 => "1111111111011101",
63739 => "1111111111011101",
63740 => "1111111111011101",
63741 => "1111111111011101",
63742 => "1111111111011101",
63743 => "1111111111011101",
63744 => "1111111111011101",
63745 => "1111111111011101",
63746 => "1111111111011101",
63747 => "1111111111011101",
63748 => "1111111111011110",
63749 => "1111111111011110",
63750 => "1111111111011110",
63751 => "1111111111011110",
63752 => "1111111111011110",
63753 => "1111111111011110",
63754 => "1111111111011110",
63755 => "1111111111011110",
63756 => "1111111111011110",
63757 => "1111111111011110",
63758 => "1111111111011110",
63759 => "1111111111011110",
63760 => "1111111111011110",
63761 => "1111111111011110",
63762 => "1111111111011110",
63763 => "1111111111011110",
63764 => "1111111111011110",
63765 => "1111111111011110",
63766 => "1111111111011110",
63767 => "1111111111011110",
63768 => "1111111111011110",
63769 => "1111111111011110",
63770 => "1111111111011110",
63771 => "1111111111011110",
63772 => "1111111111011110",
63773 => "1111111111011110",
63774 => "1111111111011110",
63775 => "1111111111011110",
63776 => "1111111111011110",
63777 => "1111111111011110",
63778 => "1111111111011110",
63779 => "1111111111011110",
63780 => "1111111111011110",
63781 => "1111111111011110",
63782 => "1111111111011110",
63783 => "1111111111011110",
63784 => "1111111111011110",
63785 => "1111111111011110",
63786 => "1111111111011110",
63787 => "1111111111011110",
63788 => "1111111111011110",
63789 => "1111111111011110",
63790 => "1111111111011110",
63791 => "1111111111011110",
63792 => "1111111111011110",
63793 => "1111111111011110",
63794 => "1111111111011110",
63795 => "1111111111011110",
63796 => "1111111111011110",
63797 => "1111111111011110",
63798 => "1111111111011110",
63799 => "1111111111011110",
63800 => "1111111111011110",
63801 => "1111111111011110",
63802 => "1111111111011110",
63803 => "1111111111011110",
63804 => "1111111111011110",
63805 => "1111111111011110",
63806 => "1111111111011110",
63807 => "1111111111011110",
63808 => "1111111111011110",
63809 => "1111111111011110",
63810 => "1111111111011110",
63811 => "1111111111011110",
63812 => "1111111111011110",
63813 => "1111111111011110",
63814 => "1111111111011110",
63815 => "1111111111011110",
63816 => "1111111111011110",
63817 => "1111111111011110",
63818 => "1111111111011110",
63819 => "1111111111011110",
63820 => "1111111111011110",
63821 => "1111111111011110",
63822 => "1111111111011110",
63823 => "1111111111011110",
63824 => "1111111111011110",
63825 => "1111111111011110",
63826 => "1111111111011110",
63827 => "1111111111011110",
63828 => "1111111111011110",
63829 => "1111111111011110",
63830 => "1111111111011110",
63831 => "1111111111011110",
63832 => "1111111111011110",
63833 => "1111111111011110",
63834 => "1111111111011110",
63835 => "1111111111011110",
63836 => "1111111111011110",
63837 => "1111111111011110",
63838 => "1111111111011110",
63839 => "1111111111011110",
63840 => "1111111111011110",
63841 => "1111111111011110",
63842 => "1111111111011110",
63843 => "1111111111011110",
63844 => "1111111111011110",
63845 => "1111111111011110",
63846 => "1111111111011110",
63847 => "1111111111011110",
63848 => "1111111111011110",
63849 => "1111111111011110",
63850 => "1111111111011110",
63851 => "1111111111011110",
63852 => "1111111111011110",
63853 => "1111111111011110",
63854 => "1111111111011110",
63855 => "1111111111011110",
63856 => "1111111111011110",
63857 => "1111111111011110",
63858 => "1111111111011110",
63859 => "1111111111011110",
63860 => "1111111111011110",
63861 => "1111111111011110",
63862 => "1111111111011110",
63863 => "1111111111011110",
63864 => "1111111111011110",
63865 => "1111111111011110",
63866 => "1111111111011110",
63867 => "1111111111011110",
63868 => "1111111111011110",
63869 => "1111111111011110",
63870 => "1111111111011111",
63871 => "1111111111011111",
63872 => "1111111111011111",
63873 => "1111111111011111",
63874 => "1111111111011111",
63875 => "1111111111011111",
63876 => "1111111111011111",
63877 => "1111111111011111",
63878 => "1111111111011111",
63879 => "1111111111011111",
63880 => "1111111111011111",
63881 => "1111111111011111",
63882 => "1111111111011111",
63883 => "1111111111011111",
63884 => "1111111111011111",
63885 => "1111111111011111",
63886 => "1111111111011111",
63887 => "1111111111011111",
63888 => "1111111111011111",
63889 => "1111111111011111",
63890 => "1111111111011111",
63891 => "1111111111011111",
63892 => "1111111111011111",
63893 => "1111111111011111",
63894 => "1111111111011111",
63895 => "1111111111011111",
63896 => "1111111111011111",
63897 => "1111111111011111",
63898 => "1111111111011111",
63899 => "1111111111011111",
63900 => "1111111111011111",
63901 => "1111111111011111",
63902 => "1111111111011111",
63903 => "1111111111011111",
63904 => "1111111111011111",
63905 => "1111111111011111",
63906 => "1111111111011111",
63907 => "1111111111011111",
63908 => "1111111111011111",
63909 => "1111111111011111",
63910 => "1111111111011111",
63911 => "1111111111011111",
63912 => "1111111111011111",
63913 => "1111111111011111",
63914 => "1111111111011111",
63915 => "1111111111011111",
63916 => "1111111111011111",
63917 => "1111111111011111",
63918 => "1111111111011111",
63919 => "1111111111011111",
63920 => "1111111111011111",
63921 => "1111111111011111",
63922 => "1111111111011111",
63923 => "1111111111011111",
63924 => "1111111111011111",
63925 => "1111111111011111",
63926 => "1111111111011111",
63927 => "1111111111011111",
63928 => "1111111111011111",
63929 => "1111111111011111",
63930 => "1111111111011111",
63931 => "1111111111011111",
63932 => "1111111111011111",
63933 => "1111111111011111",
63934 => "1111111111011111",
63935 => "1111111111011111",
63936 => "1111111111011111",
63937 => "1111111111011111",
63938 => "1111111111011111",
63939 => "1111111111011111",
63940 => "1111111111011111",
63941 => "1111111111011111",
63942 => "1111111111011111",
63943 => "1111111111011111",
63944 => "1111111111011111",
63945 => "1111111111011111",
63946 => "1111111111011111",
63947 => "1111111111011111",
63948 => "1111111111011111",
63949 => "1111111111011111",
63950 => "1111111111011111",
63951 => "1111111111011111",
63952 => "1111111111011111",
63953 => "1111111111011111",
63954 => "1111111111011111",
63955 => "1111111111011111",
63956 => "1111111111011111",
63957 => "1111111111011111",
63958 => "1111111111011111",
63959 => "1111111111011111",
63960 => "1111111111011111",
63961 => "1111111111011111",
63962 => "1111111111011111",
63963 => "1111111111011111",
63964 => "1111111111011111",
63965 => "1111111111011111",
63966 => "1111111111011111",
63967 => "1111111111011111",
63968 => "1111111111011111",
63969 => "1111111111011111",
63970 => "1111111111011111",
63971 => "1111111111011111",
63972 => "1111111111011111",
63973 => "1111111111011111",
63974 => "1111111111011111",
63975 => "1111111111011111",
63976 => "1111111111011111",
63977 => "1111111111011111",
63978 => "1111111111011111",
63979 => "1111111111011111",
63980 => "1111111111011111",
63981 => "1111111111011111",
63982 => "1111111111011111",
63983 => "1111111111011111",
63984 => "1111111111011111",
63985 => "1111111111011111",
63986 => "1111111111011111",
63987 => "1111111111011111",
63988 => "1111111111011111",
63989 => "1111111111011111",
63990 => "1111111111011111",
63991 => "1111111111011111",
63992 => "1111111111011111",
63993 => "1111111111011111",
63994 => "1111111111011111",
63995 => "1111111111011111",
63996 => "1111111111100000",
63997 => "1111111111100000",
63998 => "1111111111100000",
63999 => "1111111111100000",
64000 => "1111111111100000",
64001 => "1111111111100000",
64002 => "1111111111100000",
64003 => "1111111111100000",
64004 => "1111111111100000",
64005 => "1111111111100000",
64006 => "1111111111100000",
64007 => "1111111111100000",
64008 => "1111111111100000",
64009 => "1111111111100000",
64010 => "1111111111100000",
64011 => "1111111111100000",
64012 => "1111111111100000",
64013 => "1111111111100000",
64014 => "1111111111100000",
64015 => "1111111111100000",
64016 => "1111111111100000",
64017 => "1111111111100000",
64018 => "1111111111100000",
64019 => "1111111111100000",
64020 => "1111111111100000",
64021 => "1111111111100000",
64022 => "1111111111100000",
64023 => "1111111111100000",
64024 => "1111111111100000",
64025 => "1111111111100000",
64026 => "1111111111100000",
64027 => "1111111111100000",
64028 => "1111111111100000",
64029 => "1111111111100000",
64030 => "1111111111100000",
64031 => "1111111111100000",
64032 => "1111111111100000",
64033 => "1111111111100000",
64034 => "1111111111100000",
64035 => "1111111111100000",
64036 => "1111111111100000",
64037 => "1111111111100000",
64038 => "1111111111100000",
64039 => "1111111111100000",
64040 => "1111111111100000",
64041 => "1111111111100000",
64042 => "1111111111100000",
64043 => "1111111111100000",
64044 => "1111111111100000",
64045 => "1111111111100000",
64046 => "1111111111100000",
64047 => "1111111111100000",
64048 => "1111111111100000",
64049 => "1111111111100000",
64050 => "1111111111100000",
64051 => "1111111111100000",
64052 => "1111111111100000",
64053 => "1111111111100000",
64054 => "1111111111100000",
64055 => "1111111111100000",
64056 => "1111111111100000",
64057 => "1111111111100000",
64058 => "1111111111100000",
64059 => "1111111111100000",
64060 => "1111111111100000",
64061 => "1111111111100000",
64062 => "1111111111100000",
64063 => "1111111111100000",
64064 => "1111111111100000",
64065 => "1111111111100000",
64066 => "1111111111100000",
64067 => "1111111111100000",
64068 => "1111111111100000",
64069 => "1111111111100000",
64070 => "1111111111100000",
64071 => "1111111111100000",
64072 => "1111111111100000",
64073 => "1111111111100000",
64074 => "1111111111100000",
64075 => "1111111111100000",
64076 => "1111111111100000",
64077 => "1111111111100000",
64078 => "1111111111100000",
64079 => "1111111111100000",
64080 => "1111111111100000",
64081 => "1111111111100000",
64082 => "1111111111100000",
64083 => "1111111111100000",
64084 => "1111111111100000",
64085 => "1111111111100000",
64086 => "1111111111100000",
64087 => "1111111111100000",
64088 => "1111111111100000",
64089 => "1111111111100000",
64090 => "1111111111100000",
64091 => "1111111111100000",
64092 => "1111111111100000",
64093 => "1111111111100000",
64094 => "1111111111100000",
64095 => "1111111111100000",
64096 => "1111111111100000",
64097 => "1111111111100000",
64098 => "1111111111100000",
64099 => "1111111111100000",
64100 => "1111111111100000",
64101 => "1111111111100000",
64102 => "1111111111100000",
64103 => "1111111111100000",
64104 => "1111111111100000",
64105 => "1111111111100000",
64106 => "1111111111100000",
64107 => "1111111111100000",
64108 => "1111111111100000",
64109 => "1111111111100000",
64110 => "1111111111100000",
64111 => "1111111111100000",
64112 => "1111111111100000",
64113 => "1111111111100000",
64114 => "1111111111100000",
64115 => "1111111111100000",
64116 => "1111111111100000",
64117 => "1111111111100000",
64118 => "1111111111100000",
64119 => "1111111111100000",
64120 => "1111111111100000",
64121 => "1111111111100000",
64122 => "1111111111100000",
64123 => "1111111111100000",
64124 => "1111111111100000",
64125 => "1111111111100000",
64126 => "1111111111100001",
64127 => "1111111111100001",
64128 => "1111111111100001",
64129 => "1111111111100001",
64130 => "1111111111100001",
64131 => "1111111111100001",
64132 => "1111111111100001",
64133 => "1111111111100001",
64134 => "1111111111100001",
64135 => "1111111111100001",
64136 => "1111111111100001",
64137 => "1111111111100001",
64138 => "1111111111100001",
64139 => "1111111111100001",
64140 => "1111111111100001",
64141 => "1111111111100001",
64142 => "1111111111100001",
64143 => "1111111111100001",
64144 => "1111111111100001",
64145 => "1111111111100001",
64146 => "1111111111100001",
64147 => "1111111111100001",
64148 => "1111111111100001",
64149 => "1111111111100001",
64150 => "1111111111100001",
64151 => "1111111111100001",
64152 => "1111111111100001",
64153 => "1111111111100001",
64154 => "1111111111100001",
64155 => "1111111111100001",
64156 => "1111111111100001",
64157 => "1111111111100001",
64158 => "1111111111100001",
64159 => "1111111111100001",
64160 => "1111111111100001",
64161 => "1111111111100001",
64162 => "1111111111100001",
64163 => "1111111111100001",
64164 => "1111111111100001",
64165 => "1111111111100001",
64166 => "1111111111100001",
64167 => "1111111111100001",
64168 => "1111111111100001",
64169 => "1111111111100001",
64170 => "1111111111100001",
64171 => "1111111111100001",
64172 => "1111111111100001",
64173 => "1111111111100001",
64174 => "1111111111100001",
64175 => "1111111111100001",
64176 => "1111111111100001",
64177 => "1111111111100001",
64178 => "1111111111100001",
64179 => "1111111111100001",
64180 => "1111111111100001",
64181 => "1111111111100001",
64182 => "1111111111100001",
64183 => "1111111111100001",
64184 => "1111111111100001",
64185 => "1111111111100001",
64186 => "1111111111100001",
64187 => "1111111111100001",
64188 => "1111111111100001",
64189 => "1111111111100001",
64190 => "1111111111100001",
64191 => "1111111111100001",
64192 => "1111111111100001",
64193 => "1111111111100001",
64194 => "1111111111100001",
64195 => "1111111111100001",
64196 => "1111111111100001",
64197 => "1111111111100001",
64198 => "1111111111100001",
64199 => "1111111111100001",
64200 => "1111111111100001",
64201 => "1111111111100001",
64202 => "1111111111100001",
64203 => "1111111111100001",
64204 => "1111111111100001",
64205 => "1111111111100001",
64206 => "1111111111100001",
64207 => "1111111111100001",
64208 => "1111111111100001",
64209 => "1111111111100001",
64210 => "1111111111100001",
64211 => "1111111111100001",
64212 => "1111111111100001",
64213 => "1111111111100001",
64214 => "1111111111100001",
64215 => "1111111111100001",
64216 => "1111111111100001",
64217 => "1111111111100001",
64218 => "1111111111100001",
64219 => "1111111111100001",
64220 => "1111111111100001",
64221 => "1111111111100001",
64222 => "1111111111100001",
64223 => "1111111111100001",
64224 => "1111111111100001",
64225 => "1111111111100001",
64226 => "1111111111100001",
64227 => "1111111111100001",
64228 => "1111111111100001",
64229 => "1111111111100001",
64230 => "1111111111100001",
64231 => "1111111111100001",
64232 => "1111111111100001",
64233 => "1111111111100001",
64234 => "1111111111100001",
64235 => "1111111111100001",
64236 => "1111111111100001",
64237 => "1111111111100001",
64238 => "1111111111100001",
64239 => "1111111111100001",
64240 => "1111111111100001",
64241 => "1111111111100001",
64242 => "1111111111100001",
64243 => "1111111111100001",
64244 => "1111111111100001",
64245 => "1111111111100001",
64246 => "1111111111100001",
64247 => "1111111111100001",
64248 => "1111111111100001",
64249 => "1111111111100001",
64250 => "1111111111100001",
64251 => "1111111111100001",
64252 => "1111111111100001",
64253 => "1111111111100001",
64254 => "1111111111100001",
64255 => "1111111111100001",
64256 => "1111111111100001",
64257 => "1111111111100001",
64258 => "1111111111100001",
64259 => "1111111111100001",
64260 => "1111111111100010",
64261 => "1111111111100010",
64262 => "1111111111100010",
64263 => "1111111111100010",
64264 => "1111111111100010",
64265 => "1111111111100010",
64266 => "1111111111100010",
64267 => "1111111111100010",
64268 => "1111111111100010",
64269 => "1111111111100010",
64270 => "1111111111100010",
64271 => "1111111111100010",
64272 => "1111111111100010",
64273 => "1111111111100010",
64274 => "1111111111100010",
64275 => "1111111111100010",
64276 => "1111111111100010",
64277 => "1111111111100010",
64278 => "1111111111100010",
64279 => "1111111111100010",
64280 => "1111111111100010",
64281 => "1111111111100010",
64282 => "1111111111100010",
64283 => "1111111111100010",
64284 => "1111111111100010",
64285 => "1111111111100010",
64286 => "1111111111100010",
64287 => "1111111111100010",
64288 => "1111111111100010",
64289 => "1111111111100010",
64290 => "1111111111100010",
64291 => "1111111111100010",
64292 => "1111111111100010",
64293 => "1111111111100010",
64294 => "1111111111100010",
64295 => "1111111111100010",
64296 => "1111111111100010",
64297 => "1111111111100010",
64298 => "1111111111100010",
64299 => "1111111111100010",
64300 => "1111111111100010",
64301 => "1111111111100010",
64302 => "1111111111100010",
64303 => "1111111111100010",
64304 => "1111111111100010",
64305 => "1111111111100010",
64306 => "1111111111100010",
64307 => "1111111111100010",
64308 => "1111111111100010",
64309 => "1111111111100010",
64310 => "1111111111100010",
64311 => "1111111111100010",
64312 => "1111111111100010",
64313 => "1111111111100010",
64314 => "1111111111100010",
64315 => "1111111111100010",
64316 => "1111111111100010",
64317 => "1111111111100010",
64318 => "1111111111100010",
64319 => "1111111111100010",
64320 => "1111111111100010",
64321 => "1111111111100010",
64322 => "1111111111100010",
64323 => "1111111111100010",
64324 => "1111111111100010",
64325 => "1111111111100010",
64326 => "1111111111100010",
64327 => "1111111111100010",
64328 => "1111111111100010",
64329 => "1111111111100010",
64330 => "1111111111100010",
64331 => "1111111111100010",
64332 => "1111111111100010",
64333 => "1111111111100010",
64334 => "1111111111100010",
64335 => "1111111111100010",
64336 => "1111111111100010",
64337 => "1111111111100010",
64338 => "1111111111100010",
64339 => "1111111111100010",
64340 => "1111111111100010",
64341 => "1111111111100010",
64342 => "1111111111100010",
64343 => "1111111111100010",
64344 => "1111111111100010",
64345 => "1111111111100010",
64346 => "1111111111100010",
64347 => "1111111111100010",
64348 => "1111111111100010",
64349 => "1111111111100010",
64350 => "1111111111100010",
64351 => "1111111111100010",
64352 => "1111111111100010",
64353 => "1111111111100010",
64354 => "1111111111100010",
64355 => "1111111111100010",
64356 => "1111111111100010",
64357 => "1111111111100010",
64358 => "1111111111100010",
64359 => "1111111111100010",
64360 => "1111111111100010",
64361 => "1111111111100010",
64362 => "1111111111100010",
64363 => "1111111111100010",
64364 => "1111111111100010",
64365 => "1111111111100010",
64366 => "1111111111100010",
64367 => "1111111111100010",
64368 => "1111111111100010",
64369 => "1111111111100010",
64370 => "1111111111100010",
64371 => "1111111111100010",
64372 => "1111111111100010",
64373 => "1111111111100010",
64374 => "1111111111100010",
64375 => "1111111111100010",
64376 => "1111111111100010",
64377 => "1111111111100010",
64378 => "1111111111100010",
64379 => "1111111111100010",
64380 => "1111111111100010",
64381 => "1111111111100010",
64382 => "1111111111100010",
64383 => "1111111111100010",
64384 => "1111111111100010",
64385 => "1111111111100010",
64386 => "1111111111100010",
64387 => "1111111111100010",
64388 => "1111111111100010",
64389 => "1111111111100010",
64390 => "1111111111100010",
64391 => "1111111111100010",
64392 => "1111111111100010",
64393 => "1111111111100010",
64394 => "1111111111100010",
64395 => "1111111111100010",
64396 => "1111111111100010",
64397 => "1111111111100010",
64398 => "1111111111100010",
64399 => "1111111111100011",
64400 => "1111111111100011",
64401 => "1111111111100011",
64402 => "1111111111100011",
64403 => "1111111111100011",
64404 => "1111111111100011",
64405 => "1111111111100011",
64406 => "1111111111100011",
64407 => "1111111111100011",
64408 => "1111111111100011",
64409 => "1111111111100011",
64410 => "1111111111100011",
64411 => "1111111111100011",
64412 => "1111111111100011",
64413 => "1111111111100011",
64414 => "1111111111100011",
64415 => "1111111111100011",
64416 => "1111111111100011",
64417 => "1111111111100011",
64418 => "1111111111100011",
64419 => "1111111111100011",
64420 => "1111111111100011",
64421 => "1111111111100011",
64422 => "1111111111100011",
64423 => "1111111111100011",
64424 => "1111111111100011",
64425 => "1111111111100011",
64426 => "1111111111100011",
64427 => "1111111111100011",
64428 => "1111111111100011",
64429 => "1111111111100011",
64430 => "1111111111100011",
64431 => "1111111111100011",
64432 => "1111111111100011",
64433 => "1111111111100011",
64434 => "1111111111100011",
64435 => "1111111111100011",
64436 => "1111111111100011",
64437 => "1111111111100011",
64438 => "1111111111100011",
64439 => "1111111111100011",
64440 => "1111111111100011",
64441 => "1111111111100011",
64442 => "1111111111100011",
64443 => "1111111111100011",
64444 => "1111111111100011",
64445 => "1111111111100011",
64446 => "1111111111100011",
64447 => "1111111111100011",
64448 => "1111111111100011",
64449 => "1111111111100011",
64450 => "1111111111100011",
64451 => "1111111111100011",
64452 => "1111111111100011",
64453 => "1111111111100011",
64454 => "1111111111100011",
64455 => "1111111111100011",
64456 => "1111111111100011",
64457 => "1111111111100011",
64458 => "1111111111100011",
64459 => "1111111111100011",
64460 => "1111111111100011",
64461 => "1111111111100011",
64462 => "1111111111100011",
64463 => "1111111111100011",
64464 => "1111111111100011",
64465 => "1111111111100011",
64466 => "1111111111100011",
64467 => "1111111111100011",
64468 => "1111111111100011",
64469 => "1111111111100011",
64470 => "1111111111100011",
64471 => "1111111111100011",
64472 => "1111111111100011",
64473 => "1111111111100011",
64474 => "1111111111100011",
64475 => "1111111111100011",
64476 => "1111111111100011",
64477 => "1111111111100011",
64478 => "1111111111100011",
64479 => "1111111111100011",
64480 => "1111111111100011",
64481 => "1111111111100011",
64482 => "1111111111100011",
64483 => "1111111111100011",
64484 => "1111111111100011",
64485 => "1111111111100011",
64486 => "1111111111100011",
64487 => "1111111111100011",
64488 => "1111111111100011",
64489 => "1111111111100011",
64490 => "1111111111100011",
64491 => "1111111111100011",
64492 => "1111111111100011",
64493 => "1111111111100011",
64494 => "1111111111100011",
64495 => "1111111111100011",
64496 => "1111111111100011",
64497 => "1111111111100011",
64498 => "1111111111100011",
64499 => "1111111111100011",
64500 => "1111111111100011",
64501 => "1111111111100011",
64502 => "1111111111100011",
64503 => "1111111111100011",
64504 => "1111111111100011",
64505 => "1111111111100011",
64506 => "1111111111100011",
64507 => "1111111111100011",
64508 => "1111111111100011",
64509 => "1111111111100011",
64510 => "1111111111100011",
64511 => "1111111111100011",
64512 => "1111111111100011",
64513 => "1111111111100011",
64514 => "1111111111100011",
64515 => "1111111111100011",
64516 => "1111111111100011",
64517 => "1111111111100011",
64518 => "1111111111100011",
64519 => "1111111111100011",
64520 => "1111111111100011",
64521 => "1111111111100011",
64522 => "1111111111100011",
64523 => "1111111111100011",
64524 => "1111111111100011",
64525 => "1111111111100011",
64526 => "1111111111100011",
64527 => "1111111111100011",
64528 => "1111111111100011",
64529 => "1111111111100011",
64530 => "1111111111100011",
64531 => "1111111111100011",
64532 => "1111111111100011",
64533 => "1111111111100011",
64534 => "1111111111100011",
64535 => "1111111111100011",
64536 => "1111111111100011",
64537 => "1111111111100011",
64538 => "1111111111100011",
64539 => "1111111111100011",
64540 => "1111111111100011",
64541 => "1111111111100011",
64542 => "1111111111100011",
64543 => "1111111111100100",
64544 => "1111111111100100",
64545 => "1111111111100100",
64546 => "1111111111100100",
64547 => "1111111111100100",
64548 => "1111111111100100",
64549 => "1111111111100100",
64550 => "1111111111100100",
64551 => "1111111111100100",
64552 => "1111111111100100",
64553 => "1111111111100100",
64554 => "1111111111100100",
64555 => "1111111111100100",
64556 => "1111111111100100",
64557 => "1111111111100100",
64558 => "1111111111100100",
64559 => "1111111111100100",
64560 => "1111111111100100",
64561 => "1111111111100100",
64562 => "1111111111100100",
64563 => "1111111111100100",
64564 => "1111111111100100",
64565 => "1111111111100100",
64566 => "1111111111100100",
64567 => "1111111111100100",
64568 => "1111111111100100",
64569 => "1111111111100100",
64570 => "1111111111100100",
64571 => "1111111111100100",
64572 => "1111111111100100",
64573 => "1111111111100100",
64574 => "1111111111100100",
64575 => "1111111111100100",
64576 => "1111111111100100",
64577 => "1111111111100100",
64578 => "1111111111100100",
64579 => "1111111111100100",
64580 => "1111111111100100",
64581 => "1111111111100100",
64582 => "1111111111100100",
64583 => "1111111111100100",
64584 => "1111111111100100",
64585 => "1111111111100100",
64586 => "1111111111100100",
64587 => "1111111111100100",
64588 => "1111111111100100",
64589 => "1111111111100100",
64590 => "1111111111100100",
64591 => "1111111111100100",
64592 => "1111111111100100",
64593 => "1111111111100100",
64594 => "1111111111100100",
64595 => "1111111111100100",
64596 => "1111111111100100",
64597 => "1111111111100100",
64598 => "1111111111100100",
64599 => "1111111111100100",
64600 => "1111111111100100",
64601 => "1111111111100100",
64602 => "1111111111100100",
64603 => "1111111111100100",
64604 => "1111111111100100",
64605 => "1111111111100100",
64606 => "1111111111100100",
64607 => "1111111111100100",
64608 => "1111111111100100",
64609 => "1111111111100100",
64610 => "1111111111100100",
64611 => "1111111111100100",
64612 => "1111111111100100",
64613 => "1111111111100100",
64614 => "1111111111100100",
64615 => "1111111111100100",
64616 => "1111111111100100",
64617 => "1111111111100100",
64618 => "1111111111100100",
64619 => "1111111111100100",
64620 => "1111111111100100",
64621 => "1111111111100100",
64622 => "1111111111100100",
64623 => "1111111111100100",
64624 => "1111111111100100",
64625 => "1111111111100100",
64626 => "1111111111100100",
64627 => "1111111111100100",
64628 => "1111111111100100",
64629 => "1111111111100100",
64630 => "1111111111100100",
64631 => "1111111111100100",
64632 => "1111111111100100",
64633 => "1111111111100100",
64634 => "1111111111100100",
64635 => "1111111111100100",
64636 => "1111111111100100",
64637 => "1111111111100100",
64638 => "1111111111100100",
64639 => "1111111111100100",
64640 => "1111111111100100",
64641 => "1111111111100100",
64642 => "1111111111100100",
64643 => "1111111111100100",
64644 => "1111111111100100",
64645 => "1111111111100100",
64646 => "1111111111100100",
64647 => "1111111111100100",
64648 => "1111111111100100",
64649 => "1111111111100100",
64650 => "1111111111100100",
64651 => "1111111111100100",
64652 => "1111111111100100",
64653 => "1111111111100100",
64654 => "1111111111100100",
64655 => "1111111111100100",
64656 => "1111111111100100",
64657 => "1111111111100100",
64658 => "1111111111100100",
64659 => "1111111111100100",
64660 => "1111111111100100",
64661 => "1111111111100100",
64662 => "1111111111100100",
64663 => "1111111111100100",
64664 => "1111111111100100",
64665 => "1111111111100100",
64666 => "1111111111100100",
64667 => "1111111111100100",
64668 => "1111111111100100",
64669 => "1111111111100100",
64670 => "1111111111100100",
64671 => "1111111111100100",
64672 => "1111111111100100",
64673 => "1111111111100100",
64674 => "1111111111100100",
64675 => "1111111111100100",
64676 => "1111111111100100",
64677 => "1111111111100100",
64678 => "1111111111100100",
64679 => "1111111111100100",
64680 => "1111111111100100",
64681 => "1111111111100100",
64682 => "1111111111100100",
64683 => "1111111111100100",
64684 => "1111111111100100",
64685 => "1111111111100100",
64686 => "1111111111100100",
64687 => "1111111111100100",
64688 => "1111111111100100",
64689 => "1111111111100100",
64690 => "1111111111100100",
64691 => "1111111111100100",
64692 => "1111111111100101",
64693 => "1111111111100101",
64694 => "1111111111100101",
64695 => "1111111111100101",
64696 => "1111111111100101",
64697 => "1111111111100101",
64698 => "1111111111100101",
64699 => "1111111111100101",
64700 => "1111111111100101",
64701 => "1111111111100101",
64702 => "1111111111100101",
64703 => "1111111111100101",
64704 => "1111111111100101",
64705 => "1111111111100101",
64706 => "1111111111100101",
64707 => "1111111111100101",
64708 => "1111111111100101",
64709 => "1111111111100101",
64710 => "1111111111100101",
64711 => "1111111111100101",
64712 => "1111111111100101",
64713 => "1111111111100101",
64714 => "1111111111100101",
64715 => "1111111111100101",
64716 => "1111111111100101",
64717 => "1111111111100101",
64718 => "1111111111100101",
64719 => "1111111111100101",
64720 => "1111111111100101",
64721 => "1111111111100101",
64722 => "1111111111100101",
64723 => "1111111111100101",
64724 => "1111111111100101",
64725 => "1111111111100101",
64726 => "1111111111100101",
64727 => "1111111111100101",
64728 => "1111111111100101",
64729 => "1111111111100101",
64730 => "1111111111100101",
64731 => "1111111111100101",
64732 => "1111111111100101",
64733 => "1111111111100101",
64734 => "1111111111100101",
64735 => "1111111111100101",
64736 => "1111111111100101",
64737 => "1111111111100101",
64738 => "1111111111100101",
64739 => "1111111111100101",
64740 => "1111111111100101",
64741 => "1111111111100101",
64742 => "1111111111100101",
64743 => "1111111111100101",
64744 => "1111111111100101",
64745 => "1111111111100101",
64746 => "1111111111100101",
64747 => "1111111111100101",
64748 => "1111111111100101",
64749 => "1111111111100101",
64750 => "1111111111100101",
64751 => "1111111111100101",
64752 => "1111111111100101",
64753 => "1111111111100101",
64754 => "1111111111100101",
64755 => "1111111111100101",
64756 => "1111111111100101",
64757 => "1111111111100101",
64758 => "1111111111100101",
64759 => "1111111111100101",
64760 => "1111111111100101",
64761 => "1111111111100101",
64762 => "1111111111100101",
64763 => "1111111111100101",
64764 => "1111111111100101",
64765 => "1111111111100101",
64766 => "1111111111100101",
64767 => "1111111111100101",
64768 => "1111111111100101",
64769 => "1111111111100101",
64770 => "1111111111100101",
64771 => "1111111111100101",
64772 => "1111111111100101",
64773 => "1111111111100101",
64774 => "1111111111100101",
64775 => "1111111111100101",
64776 => "1111111111100101",
64777 => "1111111111100101",
64778 => "1111111111100101",
64779 => "1111111111100101",
64780 => "1111111111100101",
64781 => "1111111111100101",
64782 => "1111111111100101",
64783 => "1111111111100101",
64784 => "1111111111100101",
64785 => "1111111111100101",
64786 => "1111111111100101",
64787 => "1111111111100101",
64788 => "1111111111100101",
64789 => "1111111111100101",
64790 => "1111111111100101",
64791 => "1111111111100101",
64792 => "1111111111100101",
64793 => "1111111111100101",
64794 => "1111111111100101",
64795 => "1111111111100101",
64796 => "1111111111100101",
64797 => "1111111111100101",
64798 => "1111111111100101",
64799 => "1111111111100101",
64800 => "1111111111100101",
64801 => "1111111111100101",
64802 => "1111111111100101",
64803 => "1111111111100101",
64804 => "1111111111100101",
64805 => "1111111111100101",
64806 => "1111111111100101",
64807 => "1111111111100101",
64808 => "1111111111100101",
64809 => "1111111111100101",
64810 => "1111111111100101",
64811 => "1111111111100101",
64812 => "1111111111100101",
64813 => "1111111111100101",
64814 => "1111111111100101",
64815 => "1111111111100101",
64816 => "1111111111100101",
64817 => "1111111111100101",
64818 => "1111111111100101",
64819 => "1111111111100101",
64820 => "1111111111100101",
64821 => "1111111111100101",
64822 => "1111111111100101",
64823 => "1111111111100101",
64824 => "1111111111100101",
64825 => "1111111111100101",
64826 => "1111111111100101",
64827 => "1111111111100101",
64828 => "1111111111100101",
64829 => "1111111111100101",
64830 => "1111111111100101",
64831 => "1111111111100101",
64832 => "1111111111100101",
64833 => "1111111111100101",
64834 => "1111111111100101",
64835 => "1111111111100101",
64836 => "1111111111100101",
64837 => "1111111111100101",
64838 => "1111111111100101",
64839 => "1111111111100101",
64840 => "1111111111100101",
64841 => "1111111111100101",
64842 => "1111111111100101",
64843 => "1111111111100101",
64844 => "1111111111100101",
64845 => "1111111111100101",
64846 => "1111111111100101",
64847 => "1111111111100110",
64848 => "1111111111100110",
64849 => "1111111111100110",
64850 => "1111111111100110",
64851 => "1111111111100110",
64852 => "1111111111100110",
64853 => "1111111111100110",
64854 => "1111111111100110",
64855 => "1111111111100110",
64856 => "1111111111100110",
64857 => "1111111111100110",
64858 => "1111111111100110",
64859 => "1111111111100110",
64860 => "1111111111100110",
64861 => "1111111111100110",
64862 => "1111111111100110",
64863 => "1111111111100110",
64864 => "1111111111100110",
64865 => "1111111111100110",
64866 => "1111111111100110",
64867 => "1111111111100110",
64868 => "1111111111100110",
64869 => "1111111111100110",
64870 => "1111111111100110",
64871 => "1111111111100110",
64872 => "1111111111100110",
64873 => "1111111111100110",
64874 => "1111111111100110",
64875 => "1111111111100110",
64876 => "1111111111100110",
64877 => "1111111111100110",
64878 => "1111111111100110",
64879 => "1111111111100110",
64880 => "1111111111100110",
64881 => "1111111111100110",
64882 => "1111111111100110",
64883 => "1111111111100110",
64884 => "1111111111100110",
64885 => "1111111111100110",
64886 => "1111111111100110",
64887 => "1111111111100110",
64888 => "1111111111100110",
64889 => "1111111111100110",
64890 => "1111111111100110",
64891 => "1111111111100110",
64892 => "1111111111100110",
64893 => "1111111111100110",
64894 => "1111111111100110",
64895 => "1111111111100110",
64896 => "1111111111100110",
64897 => "1111111111100110",
64898 => "1111111111100110",
64899 => "1111111111100110",
64900 => "1111111111100110",
64901 => "1111111111100110",
64902 => "1111111111100110",
64903 => "1111111111100110",
64904 => "1111111111100110",
64905 => "1111111111100110",
64906 => "1111111111100110",
64907 => "1111111111100110",
64908 => "1111111111100110",
64909 => "1111111111100110",
64910 => "1111111111100110",
64911 => "1111111111100110",
64912 => "1111111111100110",
64913 => "1111111111100110",
64914 => "1111111111100110",
64915 => "1111111111100110",
64916 => "1111111111100110",
64917 => "1111111111100110",
64918 => "1111111111100110",
64919 => "1111111111100110",
64920 => "1111111111100110",
64921 => "1111111111100110",
64922 => "1111111111100110",
64923 => "1111111111100110",
64924 => "1111111111100110",
64925 => "1111111111100110",
64926 => "1111111111100110",
64927 => "1111111111100110",
64928 => "1111111111100110",
64929 => "1111111111100110",
64930 => "1111111111100110",
64931 => "1111111111100110",
64932 => "1111111111100110",
64933 => "1111111111100110",
64934 => "1111111111100110",
64935 => "1111111111100110",
64936 => "1111111111100110",
64937 => "1111111111100110",
64938 => "1111111111100110",
64939 => "1111111111100110",
64940 => "1111111111100110",
64941 => "1111111111100110",
64942 => "1111111111100110",
64943 => "1111111111100110",
64944 => "1111111111100110",
64945 => "1111111111100110",
64946 => "1111111111100110",
64947 => "1111111111100110",
64948 => "1111111111100110",
64949 => "1111111111100110",
64950 => "1111111111100110",
64951 => "1111111111100110",
64952 => "1111111111100110",
64953 => "1111111111100110",
64954 => "1111111111100110",
64955 => "1111111111100110",
64956 => "1111111111100110",
64957 => "1111111111100110",
64958 => "1111111111100110",
64959 => "1111111111100110",
64960 => "1111111111100110",
64961 => "1111111111100110",
64962 => "1111111111100110",
64963 => "1111111111100110",
64964 => "1111111111100110",
64965 => "1111111111100110",
64966 => "1111111111100110",
64967 => "1111111111100110",
64968 => "1111111111100110",
64969 => "1111111111100110",
64970 => "1111111111100110",
64971 => "1111111111100110",
64972 => "1111111111100110",
64973 => "1111111111100110",
64974 => "1111111111100110",
64975 => "1111111111100110",
64976 => "1111111111100110",
64977 => "1111111111100110",
64978 => "1111111111100110",
64979 => "1111111111100110",
64980 => "1111111111100110",
64981 => "1111111111100110",
64982 => "1111111111100110",
64983 => "1111111111100110",
64984 => "1111111111100110",
64985 => "1111111111100110",
64986 => "1111111111100110",
64987 => "1111111111100110",
64988 => "1111111111100110",
64989 => "1111111111100110",
64990 => "1111111111100110",
64991 => "1111111111100110",
64992 => "1111111111100110",
64993 => "1111111111100110",
64994 => "1111111111100110",
64995 => "1111111111100110",
64996 => "1111111111100110",
64997 => "1111111111100110",
64998 => "1111111111100110",
64999 => "1111111111100110",
65000 => "1111111111100110",
65001 => "1111111111100110",
65002 => "1111111111100110",
65003 => "1111111111100110",
65004 => "1111111111100110",
65005 => "1111111111100110",
65006 => "1111111111100110",
65007 => "1111111111100110",
65008 => "1111111111100111",
65009 => "1111111111100111",
65010 => "1111111111100111",
65011 => "1111111111100111",
65012 => "1111111111100111",
65013 => "1111111111100111",
65014 => "1111111111100111",
65015 => "1111111111100111",
65016 => "1111111111100111",
65017 => "1111111111100111",
65018 => "1111111111100111",
65019 => "1111111111100111",
65020 => "1111111111100111",
65021 => "1111111111100111",
65022 => "1111111111100111",
65023 => "1111111111100111",
65024 => "1111111111100111",
65025 => "1111111111100111",
65026 => "1111111111100111",
65027 => "1111111111100111",
65028 => "1111111111100111",
65029 => "1111111111100111",
65030 => "1111111111100111",
65031 => "1111111111100111",
65032 => "1111111111100111",
65033 => "1111111111100111",
65034 => "1111111111100111",
65035 => "1111111111100111",
65036 => "1111111111100111",
65037 => "1111111111100111",
65038 => "1111111111100111",
65039 => "1111111111100111",
65040 => "1111111111100111",
65041 => "1111111111100111",
65042 => "1111111111100111",
65043 => "1111111111100111",
65044 => "1111111111100111",
65045 => "1111111111100111",
65046 => "1111111111100111",
65047 => "1111111111100111",
65048 => "1111111111100111",
65049 => "1111111111100111",
65050 => "1111111111100111",
65051 => "1111111111100111",
65052 => "1111111111100111",
65053 => "1111111111100111",
65054 => "1111111111100111",
65055 => "1111111111100111",
65056 => "1111111111100111",
65057 => "1111111111100111",
65058 => "1111111111100111",
65059 => "1111111111100111",
65060 => "1111111111100111",
65061 => "1111111111100111",
65062 => "1111111111100111",
65063 => "1111111111100111",
65064 => "1111111111100111",
65065 => "1111111111100111",
65066 => "1111111111100111",
65067 => "1111111111100111",
65068 => "1111111111100111",
65069 => "1111111111100111",
65070 => "1111111111100111",
65071 => "1111111111100111",
65072 => "1111111111100111",
65073 => "1111111111100111",
65074 => "1111111111100111",
65075 => "1111111111100111",
65076 => "1111111111100111",
65077 => "1111111111100111",
65078 => "1111111111100111",
65079 => "1111111111100111",
65080 => "1111111111100111",
65081 => "1111111111100111",
65082 => "1111111111100111",
65083 => "1111111111100111",
65084 => "1111111111100111",
65085 => "1111111111100111",
65086 => "1111111111100111",
65087 => "1111111111100111",
65088 => "1111111111100111",
65089 => "1111111111100111",
65090 => "1111111111100111",
65091 => "1111111111100111",
65092 => "1111111111100111",
65093 => "1111111111100111",
65094 => "1111111111100111",
65095 => "1111111111100111",
65096 => "1111111111100111",
65097 => "1111111111100111",
65098 => "1111111111100111",
65099 => "1111111111100111",
65100 => "1111111111100111",
65101 => "1111111111100111",
65102 => "1111111111100111",
65103 => "1111111111100111",
65104 => "1111111111100111",
65105 => "1111111111100111",
65106 => "1111111111100111",
65107 => "1111111111100111",
65108 => "1111111111100111",
65109 => "1111111111100111",
65110 => "1111111111100111",
65111 => "1111111111100111",
65112 => "1111111111100111",
65113 => "1111111111100111",
65114 => "1111111111100111",
65115 => "1111111111100111",
65116 => "1111111111100111",
65117 => "1111111111100111",
65118 => "1111111111100111",
65119 => "1111111111100111",
65120 => "1111111111100111",
65121 => "1111111111100111",
65122 => "1111111111100111",
65123 => "1111111111100111",
65124 => "1111111111100111",
65125 => "1111111111100111",
65126 => "1111111111100111",
65127 => "1111111111100111",
65128 => "1111111111100111",
65129 => "1111111111100111",
65130 => "1111111111100111",
65131 => "1111111111100111",
65132 => "1111111111100111",
65133 => "1111111111100111",
65134 => "1111111111100111",
65135 => "1111111111100111",
65136 => "1111111111100111",
65137 => "1111111111100111",
65138 => "1111111111100111",
65139 => "1111111111100111",
65140 => "1111111111100111",
65141 => "1111111111100111",
65142 => "1111111111100111",
65143 => "1111111111100111",
65144 => "1111111111100111",
65145 => "1111111111100111",
65146 => "1111111111100111",
65147 => "1111111111100111",
65148 => "1111111111100111",
65149 => "1111111111100111",
65150 => "1111111111100111",
65151 => "1111111111100111",
65152 => "1111111111100111",
65153 => "1111111111100111",
65154 => "1111111111100111",
65155 => "1111111111100111",
65156 => "1111111111100111",
65157 => "1111111111100111",
65158 => "1111111111100111",
65159 => "1111111111100111",
65160 => "1111111111100111",
65161 => "1111111111100111",
65162 => "1111111111100111",
65163 => "1111111111100111",
65164 => "1111111111100111",
65165 => "1111111111100111",
65166 => "1111111111100111",
65167 => "1111111111100111",
65168 => "1111111111100111",
65169 => "1111111111100111",
65170 => "1111111111100111",
65171 => "1111111111100111",
65172 => "1111111111100111",
65173 => "1111111111100111",
65174 => "1111111111100111",
65175 => "1111111111101000",
65176 => "1111111111101000",
65177 => "1111111111101000",
65178 => "1111111111101000",
65179 => "1111111111101000",
65180 => "1111111111101000",
65181 => "1111111111101000",
65182 => "1111111111101000",
65183 => "1111111111101000",
65184 => "1111111111101000",
65185 => "1111111111101000",
65186 => "1111111111101000",
65187 => "1111111111101000",
65188 => "1111111111101000",
65189 => "1111111111101000",
65190 => "1111111111101000",
65191 => "1111111111101000",
65192 => "1111111111101000",
65193 => "1111111111101000",
65194 => "1111111111101000",
65195 => "1111111111101000",
65196 => "1111111111101000",
65197 => "1111111111101000",
65198 => "1111111111101000",
65199 => "1111111111101000",
65200 => "1111111111101000",
65201 => "1111111111101000",
65202 => "1111111111101000",
65203 => "1111111111101000",
65204 => "1111111111101000",
65205 => "1111111111101000",
65206 => "1111111111101000",
65207 => "1111111111101000",
65208 => "1111111111101000",
65209 => "1111111111101000",
65210 => "1111111111101000",
65211 => "1111111111101000",
65212 => "1111111111101000",
65213 => "1111111111101000",
65214 => "1111111111101000",
65215 => "1111111111101000",
65216 => "1111111111101000",
65217 => "1111111111101000",
65218 => "1111111111101000",
65219 => "1111111111101000",
65220 => "1111111111101000",
65221 => "1111111111101000",
65222 => "1111111111101000",
65223 => "1111111111101000",
65224 => "1111111111101000",
65225 => "1111111111101000",
65226 => "1111111111101000",
65227 => "1111111111101000",
65228 => "1111111111101000",
65229 => "1111111111101000",
65230 => "1111111111101000",
65231 => "1111111111101000",
65232 => "1111111111101000",
65233 => "1111111111101000",
65234 => "1111111111101000",
65235 => "1111111111101000",
65236 => "1111111111101000",
65237 => "1111111111101000",
65238 => "1111111111101000",
65239 => "1111111111101000",
65240 => "1111111111101000",
65241 => "1111111111101000",
65242 => "1111111111101000",
65243 => "1111111111101000",
65244 => "1111111111101000",
65245 => "1111111111101000",
65246 => "1111111111101000",
65247 => "1111111111101000",
65248 => "1111111111101000",
65249 => "1111111111101000",
65250 => "1111111111101000",
65251 => "1111111111101000",
65252 => "1111111111101000",
65253 => "1111111111101000",
65254 => "1111111111101000",
65255 => "1111111111101000",
65256 => "1111111111101000",
65257 => "1111111111101000",
65258 => "1111111111101000",
65259 => "1111111111101000",
65260 => "1111111111101000",
65261 => "1111111111101000",
65262 => "1111111111101000",
65263 => "1111111111101000",
65264 => "1111111111101000",
65265 => "1111111111101000",
65266 => "1111111111101000",
65267 => "1111111111101000",
65268 => "1111111111101000",
65269 => "1111111111101000",
65270 => "1111111111101000",
65271 => "1111111111101000",
65272 => "1111111111101000",
65273 => "1111111111101000",
65274 => "1111111111101000",
65275 => "1111111111101000",
65276 => "1111111111101000",
65277 => "1111111111101000",
65278 => "1111111111101000",
65279 => "1111111111101000",
65280 => "1111111111101000",
65281 => "1111111111101000",
65282 => "1111111111101000",
65283 => "1111111111101000",
65284 => "1111111111101000",
65285 => "1111111111101000",
65286 => "1111111111101000",
65287 => "1111111111101000",
65288 => "1111111111101000",
65289 => "1111111111101000",
65290 => "1111111111101000",
65291 => "1111111111101000",
65292 => "1111111111101000",
65293 => "1111111111101000",
65294 => "1111111111101000",
65295 => "1111111111101000",
65296 => "1111111111101000",
65297 => "1111111111101000",
65298 => "1111111111101000",
65299 => "1111111111101000",
65300 => "1111111111101000",
65301 => "1111111111101000",
65302 => "1111111111101000",
65303 => "1111111111101000",
65304 => "1111111111101000",
65305 => "1111111111101000",
65306 => "1111111111101000",
65307 => "1111111111101000",
65308 => "1111111111101000",
65309 => "1111111111101000",
65310 => "1111111111101000",
65311 => "1111111111101000",
65312 => "1111111111101000",
65313 => "1111111111101000",
65314 => "1111111111101000",
65315 => "1111111111101000",
65316 => "1111111111101000",
65317 => "1111111111101000",
65318 => "1111111111101000",
65319 => "1111111111101000",
65320 => "1111111111101000",
65321 => "1111111111101000",
65322 => "1111111111101000",
65323 => "1111111111101000",
65324 => "1111111111101000",
65325 => "1111111111101000",
65326 => "1111111111101000",
65327 => "1111111111101000",
65328 => "1111111111101000",
65329 => "1111111111101000",
65330 => "1111111111101000",
65331 => "1111111111101000",
65332 => "1111111111101000",
65333 => "1111111111101000",
65334 => "1111111111101000",
65335 => "1111111111101000",
65336 => "1111111111101000",
65337 => "1111111111101000",
65338 => "1111111111101000",
65339 => "1111111111101000",
65340 => "1111111111101000",
65341 => "1111111111101000",
65342 => "1111111111101000",
65343 => "1111111111101000",
65344 => "1111111111101000",
65345 => "1111111111101000",
65346 => "1111111111101000",
65347 => "1111111111101000",
65348 => "1111111111101000",
65349 => "1111111111101001",
65350 => "1111111111101001",
65351 => "1111111111101001",
65352 => "1111111111101001",
65353 => "1111111111101001",
65354 => "1111111111101001",
65355 => "1111111111101001",
65356 => "1111111111101001",
65357 => "1111111111101001",
65358 => "1111111111101001",
65359 => "1111111111101001",
65360 => "1111111111101001",
65361 => "1111111111101001",
65362 => "1111111111101001",
65363 => "1111111111101001",
65364 => "1111111111101001",
65365 => "1111111111101001",
65366 => "1111111111101001",
65367 => "1111111111101001",
65368 => "1111111111101001",
65369 => "1111111111101001",
65370 => "1111111111101001",
65371 => "1111111111101001",
65372 => "1111111111101001",
65373 => "1111111111101001",
65374 => "1111111111101001",
65375 => "1111111111101001",
65376 => "1111111111101001",
65377 => "1111111111101001",
65378 => "1111111111101001",
65379 => "1111111111101001",
65380 => "1111111111101001",
65381 => "1111111111101001",
65382 => "1111111111101001",
65383 => "1111111111101001",
65384 => "1111111111101001",
65385 => "1111111111101001",
65386 => "1111111111101001",
65387 => "1111111111101001",
65388 => "1111111111101001",
65389 => "1111111111101001",
65390 => "1111111111101001",
65391 => "1111111111101001",
65392 => "1111111111101001",
65393 => "1111111111101001",
65394 => "1111111111101001",
65395 => "1111111111101001",
65396 => "1111111111101001",
65397 => "1111111111101001",
65398 => "1111111111101001",
65399 => "1111111111101001",
65400 => "1111111111101001",
65401 => "1111111111101001",
65402 => "1111111111101001",
65403 => "1111111111101001",
65404 => "1111111111101001",
65405 => "1111111111101001",
65406 => "1111111111101001",
65407 => "1111111111101001",
65408 => "1111111111101001",
65409 => "1111111111101001",
65410 => "1111111111101001",
65411 => "1111111111101001",
65412 => "1111111111101001",
65413 => "1111111111101001",
65414 => "1111111111101001",
65415 => "1111111111101001",
65416 => "1111111111101001",
65417 => "1111111111101001",
65418 => "1111111111101001",
65419 => "1111111111101001",
65420 => "1111111111101001",
65421 => "1111111111101001",
65422 => "1111111111101001",
65423 => "1111111111101001",
65424 => "1111111111101001",
65425 => "1111111111101001",
65426 => "1111111111101001",
65427 => "1111111111101001",
65428 => "1111111111101001",
65429 => "1111111111101001",
65430 => "1111111111101001",
65431 => "1111111111101001",
65432 => "1111111111101001",
65433 => "1111111111101001",
65434 => "1111111111101001",
65435 => "1111111111101001",
65436 => "1111111111101001",
65437 => "1111111111101001",
65438 => "1111111111101001",
65439 => "1111111111101001",
65440 => "1111111111101001",
65441 => "1111111111101001",
65442 => "1111111111101001",
65443 => "1111111111101001",
65444 => "1111111111101001",
65445 => "1111111111101001",
65446 => "1111111111101001",
65447 => "1111111111101001",
65448 => "1111111111101001",
65449 => "1111111111101001",
65450 => "1111111111101001",
65451 => "1111111111101001",
65452 => "1111111111101001",
65453 => "1111111111101001",
65454 => "1111111111101001",
65455 => "1111111111101001",
65456 => "1111111111101001",
65457 => "1111111111101001",
65458 => "1111111111101001",
65459 => "1111111111101001",
65460 => "1111111111101001",
65461 => "1111111111101001",
65462 => "1111111111101001",
65463 => "1111111111101001",
65464 => "1111111111101001",
65465 => "1111111111101001",
65466 => "1111111111101001",
65467 => "1111111111101001",
65468 => "1111111111101001",
65469 => "1111111111101001",
65470 => "1111111111101001",
65471 => "1111111111101001",
65472 => "1111111111101001",
65473 => "1111111111101001",
65474 => "1111111111101001",
65475 => "1111111111101001",
65476 => "1111111111101001",
65477 => "1111111111101001",
65478 => "1111111111101001",
65479 => "1111111111101001",
65480 => "1111111111101001",
65481 => "1111111111101001",
65482 => "1111111111101001",
65483 => "1111111111101001",
65484 => "1111111111101001",
65485 => "1111111111101001",
65486 => "1111111111101001",
65487 => "1111111111101001",
65488 => "1111111111101001",
65489 => "1111111111101001",
65490 => "1111111111101001",
65491 => "1111111111101001",
65492 => "1111111111101001",
65493 => "1111111111101001",
65494 => "1111111111101001",
65495 => "1111111111101001",
65496 => "1111111111101001",
65497 => "1111111111101001",
65498 => "1111111111101001",
65499 => "1111111111101001",
65500 => "1111111111101001",
65501 => "1111111111101001",
65502 => "1111111111101001",
65503 => "1111111111101001",
65504 => "1111111111101001",
65505 => "1111111111101001",
65506 => "1111111111101001",
65507 => "1111111111101001",
65508 => "1111111111101001",
65509 => "1111111111101001",
65510 => "1111111111101001",
65511 => "1111111111101001",
65512 => "1111111111101001",
65513 => "1111111111101001",
65514 => "1111111111101001",
65515 => "1111111111101001",
65516 => "1111111111101001",
65517 => "1111111111101001",
65518 => "1111111111101001",
65519 => "1111111111101001",
65520 => "1111111111101001",
65521 => "1111111111101001",
65522 => "1111111111101001",
65523 => "1111111111101001",
65524 => "1111111111101001",
65525 => "1111111111101001",
65526 => "1111111111101001",
65527 => "1111111111101001",
65528 => "1111111111101001",
65529 => "1111111111101001",
65530 => "1111111111101001",
65531 => "1111111111101010",
65532 => "1111111111101010",
65533 => "1111111111101010",
65534 => "1111111111101010",
65535 => "1111111111101010"

    );	 
	 
begin
	
		
	data_val <= lut_data(address);
		
		
		
		
		
		
		
		
		

end archLUT;