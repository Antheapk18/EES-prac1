library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- need entity
entity prac_16bits is
port(

clk: in std_logic; -- this is 50 MHz clock on PIN_V11 
rx : in std_logic; -- PIN_AH27

tx: out std_logic); -- just choose a random PIN_AG28

end prac_16bits;

-- will start with behavioural logic but will need to change to structural
architecture UART of prac_16bits is
	--signal tx_value : std_logic_vector(7 downto 0) := "00000000";
	--signal tx_value2 : std_logic_vector(7 downto 0) := "00000000";
	signal data_reg : std_logic_vector(15 downto 0) := "0000000000000000";
	signal rx_value : std_logic_vector(7 downto 0) := "00000000";
	signal tx_counter : integer := 0;
	signal rx_counter : integer := 0;
	signal baud_counter: integer := 0;
	signal baudReceive_counter: integer := 0;
	signal flag_receive :integer := 0; -- flag to be set when allowed to transmit data back
	signal CounterLUT: integer := 0;
	type lut_array is array (0 to 65535) of std_logic_vector(15 downto 0);
	constant lut_data : lut_array := (
0 => "0000000000001010",
1 => "0000000000001010",
2 => "0000000000001010",
3 => "0000000000001011",
4 => "0000000000001011",
5 => "0000000000001011",
6 => "0000000000001011",
7 => "0000000000001011",
8 => "0000000000001011",
9 => "0000000000001011",
10 => "0000000000001011",
11 => "0000000000001011",
12 => "0000000000001011",
13 => "0000000000001011",
14 => "0000000000001011",
15 => "0000000000001011",
16 => "0000000000001011",
17 => "0000000000001011",
18 => "0000000000001011",
19 => "0000000000001011",
20 => "0000000000001011",
21 => "0000000000001011",
22 => "0000000000001011",
23 => "0000000000001011",
24 => "0000000000001011",
25 => "0000000000001011",
26 => "0000000000001011",
27 => "0000000000001011",
28 => "0000000000001011",
29 => "0000000000001011",
30 => "0000000000001011",
31 => "0000000000001011",
32 => "0000000000001011",
33 => "0000000000001011",
34 => "0000000000001011",
35 => "0000000000001011",
36 => "0000000000001011",
37 => "0000000000001011",
38 => "0000000000001011",
39 => "0000000000001011",
40 => "0000000000001011",
41 => "0000000000001011",
42 => "0000000000001011",
43 => "0000000000001011",
44 => "0000000000001011",
45 => "0000000000001011",
46 => "0000000000001011",
47 => "0000000000001011",
48 => "0000000000001011",
49 => "0000000000001011",
50 => "0000000000001011",
51 => "0000000000001011",
52 => "0000000000001011",
53 => "0000000000001011",
54 => "0000000000001011",
55 => "0000000000001011",
56 => "0000000000001011",
57 => "0000000000001011",
58 => "0000000000001011",
59 => "0000000000001011",
60 => "0000000000001011",
61 => "0000000000001011",
62 => "0000000000001011",
63 => "0000000000001011",
64 => "0000000000001011",
65 => "0000000000001011",
66 => "0000000000001011",
67 => "0000000000001011",
68 => "0000000000001011",
69 => "0000000000001011",
70 => "0000000000001011",
71 => "0000000000001011",
72 => "0000000000001011",
73 => "0000000000001011",
74 => "0000000000001011",
75 => "0000000000001011",
76 => "0000000000001011",
77 => "0000000000001011",
78 => "0000000000001011",
79 => "0000000000001011",
80 => "0000000000001011",
81 => "0000000000001011",
82 => "0000000000001011",
83 => "0000000000001011",
84 => "0000000000001011",
85 => "0000000000001011",
86 => "0000000000001011",
87 => "0000000000001011",
88 => "0000000000001011",
89 => "0000000000001011",
90 => "0000000000001011",
91 => "0000000000001011",
92 => "0000000000001011",
93 => "0000000000001011",
94 => "0000000000001011",
95 => "0000000000001011",
96 => "0000000000001011",
97 => "0000000000001011",
98 => "0000000000001011",
99 => "0000000000001011",
100 => "0000000000001011",
101 => "0000000000001011",
102 => "0000000000001011",
103 => "0000000000001011",
104 => "0000000000001011",
105 => "0000000000001011",
106 => "0000000000001011",
107 => "0000000000001011",
108 => "0000000000001011",
109 => "0000000000001011",
110 => "0000000000001011",
111 => "0000000000001011",
112 => "0000000000001011",
113 => "0000000000001011",
114 => "0000000000001011",
115 => "0000000000001011",
116 => "0000000000001011",
117 => "0000000000001011",
118 => "0000000000001011",
119 => "0000000000001011",
120 => "0000000000001011",
121 => "0000000000001011",
122 => "0000000000001011",
123 => "0000000000001011",
124 => "0000000000001011",
125 => "0000000000001011",
126 => "0000000000001011",
127 => "0000000000001011",
128 => "0000000000001011",
129 => "0000000000001011",
130 => "0000000000001011",
131 => "0000000000001011",
132 => "0000000000001011",
133 => "0000000000001011",
134 => "0000000000001011",
135 => "0000000000001011",
136 => "0000000000001011",
137 => "0000000000001011",
138 => "0000000000001011",
139 => "0000000000001011",
140 => "0000000000001011",
141 => "0000000000001011",
142 => "0000000000001011",
143 => "0000000000001011",
144 => "0000000000001011",
145 => "0000000000001011",
146 => "0000000000001011",
147 => "0000000000001011",
148 => "0000000000001011",
149 => "0000000000001011",
150 => "0000000000001011",
151 => "0000000000001011",
152 => "0000000000001011",
153 => "0000000000001011",
154 => "0000000000001011",
155 => "0000000000001011",
156 => "0000000000001011",
157 => "0000000000001011",
158 => "0000000000001011",
159 => "0000000000001011",
160 => "0000000000001011",
161 => "0000000000001011",
162 => "0000000000001011",
163 => "0000000000001011",
164 => "0000000000001011",
165 => "0000000000001011",
166 => "0000000000001011",
167 => "0000000000001011",
168 => "0000000000001011",
169 => "0000000000001011",
170 => "0000000000001011",
171 => "0000000000001011",
172 => "0000000000001011",
173 => "0000000000001011",
174 => "0000000000001011",
175 => "0000000000001011",
176 => "0000000000001011",
177 => "0000000000001011",
178 => "0000000000001011",
179 => "0000000000001011",
180 => "0000000000001011",
181 => "0000000000001011",
182 => "0000000000001011",
183 => "0000000000001011",
184 => "0000000000001011",
185 => "0000000000001011",
186 => "0000000000001011",
187 => "0000000000001011",
188 => "0000000000001011",
189 => "0000000000001011",
190 => "0000000000001011",
191 => "0000000000001011",
192 => "0000000000001011",
193 => "0000000000001011",
194 => "0000000000001011",
195 => "0000000000001011",
196 => "0000000000001011",
197 => "0000000000001011",
198 => "0000000000001011",
199 => "0000000000001011",
200 => "0000000000001011",
201 => "0000000000001011",
202 => "0000000000001011",
203 => "0000000000001011",
204 => "0000000000001011",
205 => "0000000000001011",
206 => "0000000000001011",
207 => "0000000000001011",
208 => "0000000000001011",
209 => "0000000000001011",
210 => "0000000000001011",
211 => "0000000000001011",
212 => "0000000000001011",
213 => "0000000000001011",
214 => "0000000000001011",
215 => "0000000000001011",
216 => "0000000000001011",
217 => "0000000000001011",
218 => "0000000000001011",
219 => "0000000000001011",
220 => "0000000000001011",
221 => "0000000000001011",
222 => "0000000000001011",
223 => "0000000000001011",
224 => "0000000000001011",
225 => "0000000000001011",
226 => "0000000000001011",
227 => "0000000000001011",
228 => "0000000000001011",
229 => "0000000000001011",
230 => "0000000000001011",
231 => "0000000000001011",
232 => "0000000000001011",
233 => "0000000000001011",
234 => "0000000000001011",
235 => "0000000000001011",
236 => "0000000000001011",
237 => "0000000000001011",
238 => "0000000000001011",
239 => "0000000000001011",
240 => "0000000000001011",
241 => "0000000000001011",
242 => "0000000000001011",
243 => "0000000000001011",
244 => "0000000000001011",
245 => "0000000000001011",
246 => "0000000000001011",
247 => "0000000000001011",
248 => "0000000000001011",
249 => "0000000000001011",
250 => "0000000000001011",
251 => "0000000000001011",
252 => "0000000000001011",
253 => "0000000000001011",
254 => "0000000000001011",
255 => "0000000000001011",
256 => "0000000000001011",
257 => "0000000000001011",
258 => "0000000000001011",
259 => "0000000000001011",
260 => "0000000000001011",
261 => "0000000000001011",
262 => "0000000000001011",
263 => "0000000000001011",
264 => "0000000000001011",
265 => "0000000000001011",
266 => "0000000000001011",
267 => "0000000000001011",
268 => "0000000000001011",
269 => "0000000000001011",
270 => "0000000000001011",
271 => "0000000000001011",
272 => "0000000000001011",
273 => "0000000000001011",
274 => "0000000000001011",
275 => "0000000000001011",
276 => "0000000000001011",
277 => "0000000000001011",
278 => "0000000000001011",
279 => "0000000000001011",
280 => "0000000000001011",
281 => "0000000000001011",
282 => "0000000000001011",
283 => "0000000000001011",
284 => "0000000000001011",
285 => "0000000000001011",
286 => "0000000000001011",
287 => "0000000000001011",
288 => "0000000000001011",
289 => "0000000000001011",
290 => "0000000000001011",
291 => "0000000000001011",
292 => "0000000000001011",
293 => "0000000000001011",
294 => "0000000000001011",
295 => "0000000000001011",
296 => "0000000000001011",
297 => "0000000000001011",
298 => "0000000000001011",
299 => "0000000000001011",
300 => "0000000000001011",
301 => "0000000000001011",
302 => "0000000000001011",
303 => "0000000000001011",
304 => "0000000000001011",
305 => "0000000000001011",
306 => "0000000000001011",
307 => "0000000000001011",
308 => "0000000000001011",
309 => "0000000000001011",
310 => "0000000000001011",
311 => "0000000000001011",
312 => "0000000000001011",
313 => "0000000000001011",
314 => "0000000000001011",
315 => "0000000000001011",
316 => "0000000000001011",
317 => "0000000000001011",
318 => "0000000000001011",
319 => "0000000000001011",
320 => "0000000000001011",
321 => "0000000000001011",
322 => "0000000000001011",
323 => "0000000000001011",
324 => "0000000000001011",
325 => "0000000000001011",
326 => "0000000000001011",
327 => "0000000000001011",
328 => "0000000000001011",
329 => "0000000000001011",
330 => "0000000000001011",
331 => "0000000000001011",
332 => "0000000000001011",
333 => "0000000000001011",
334 => "0000000000001011",
335 => "0000000000001011",
336 => "0000000000001011",
337 => "0000000000001011",
338 => "0000000000001011",
339 => "0000000000001011",
340 => "0000000000001011",
341 => "0000000000001011",
342 => "0000000000001011",
343 => "0000000000001011",
344 => "0000000000001011",
345 => "0000000000001011",
346 => "0000000000001011",
347 => "0000000000001011",
348 => "0000000000001011",
349 => "0000000000001011",
350 => "0000000000001011",
351 => "0000000000001011",
352 => "0000000000001011",
353 => "0000000000001011",
354 => "0000000000001011",
355 => "0000000000001011",
356 => "0000000000001011",
357 => "0000000000001011",
358 => "0000000000001011",
359 => "0000000000001011",
360 => "0000000000001100",
361 => "0000000000001100",
362 => "0000000000001100",
363 => "0000000000001100",
364 => "0000000000001100",
365 => "0000000000001100",
366 => "0000000000001100",
367 => "0000000000001100",
368 => "0000000000001100",
369 => "0000000000001100",
370 => "0000000000001100",
371 => "0000000000001100",
372 => "0000000000001100",
373 => "0000000000001100",
374 => "0000000000001100",
375 => "0000000000001100",
376 => "0000000000001100",
377 => "0000000000001100",
378 => "0000000000001100",
379 => "0000000000001100",
380 => "0000000000001100",
381 => "0000000000001100",
382 => "0000000000001100",
383 => "0000000000001100",
384 => "0000000000001100",
385 => "0000000000001100",
386 => "0000000000001100",
387 => "0000000000001100",
388 => "0000000000001100",
389 => "0000000000001100",
390 => "0000000000001100",
391 => "0000000000001100",
392 => "0000000000001100",
393 => "0000000000001100",
394 => "0000000000001100",
395 => "0000000000001100",
396 => "0000000000001100",
397 => "0000000000001100",
398 => "0000000000001100",
399 => "0000000000001100",
400 => "0000000000001100",
401 => "0000000000001100",
402 => "0000000000001100",
403 => "0000000000001100",
404 => "0000000000001100",
405 => "0000000000001100",
406 => "0000000000001100",
407 => "0000000000001100",
408 => "0000000000001100",
409 => "0000000000001100",
410 => "0000000000001100",
411 => "0000000000001100",
412 => "0000000000001100",
413 => "0000000000001100",
414 => "0000000000001100",
415 => "0000000000001100",
416 => "0000000000001100",
417 => "0000000000001100",
418 => "0000000000001100",
419 => "0000000000001100",
420 => "0000000000001100",
421 => "0000000000001100",
422 => "0000000000001100",
423 => "0000000000001100",
424 => "0000000000001100",
425 => "0000000000001100",
426 => "0000000000001100",
427 => "0000000000001100",
428 => "0000000000001100",
429 => "0000000000001100",
430 => "0000000000001100",
431 => "0000000000001100",
432 => "0000000000001100",
433 => "0000000000001100",
434 => "0000000000001100",
435 => "0000000000001100",
436 => "0000000000001100",
437 => "0000000000001100",
438 => "0000000000001100",
439 => "0000000000001100",
440 => "0000000000001100",
441 => "0000000000001100",
442 => "0000000000001100",
443 => "0000000000001100",
444 => "0000000000001100",
445 => "0000000000001100",
446 => "0000000000001100",
447 => "0000000000001100",
448 => "0000000000001100",
449 => "0000000000001100",
450 => "0000000000001100",
451 => "0000000000001100",
452 => "0000000000001100",
453 => "0000000000001100",
454 => "0000000000001100",
455 => "0000000000001100",
456 => "0000000000001100",
457 => "0000000000001100",
458 => "0000000000001100",
459 => "0000000000001100",
460 => "0000000000001100",
461 => "0000000000001100",
462 => "0000000000001100",
463 => "0000000000001100",
464 => "0000000000001100",
465 => "0000000000001100",
466 => "0000000000001100",
467 => "0000000000001100",
468 => "0000000000001100",
469 => "0000000000001100",
470 => "0000000000001100",
471 => "0000000000001100",
472 => "0000000000001100",
473 => "0000000000001100",
474 => "0000000000001100",
475 => "0000000000001100",
476 => "0000000000001100",
477 => "0000000000001100",
478 => "0000000000001100",
479 => "0000000000001100",
480 => "0000000000001100",
481 => "0000000000001100",
482 => "0000000000001100",
483 => "0000000000001100",
484 => "0000000000001100",
485 => "0000000000001100",
486 => "0000000000001100",
487 => "0000000000001100",
488 => "0000000000001100",
489 => "0000000000001100",
490 => "0000000000001100",
491 => "0000000000001100",
492 => "0000000000001100",
493 => "0000000000001100",
494 => "0000000000001100",
495 => "0000000000001100",
496 => "0000000000001100",
497 => "0000000000001100",
498 => "0000000000001100",
499 => "0000000000001100",
500 => "0000000000001100",
501 => "0000000000001100",
502 => "0000000000001100",
503 => "0000000000001100",
504 => "0000000000001100",
505 => "0000000000001100",
506 => "0000000000001100",
507 => "0000000000001100",
508 => "0000000000001100",
509 => "0000000000001100",
510 => "0000000000001100",
511 => "0000000000001100",
512 => "0000000000001100",
513 => "0000000000001100",
514 => "0000000000001100",
515 => "0000000000001100",
516 => "0000000000001100",
517 => "0000000000001100",
518 => "0000000000001100",
519 => "0000000000001100",
520 => "0000000000001100",
521 => "0000000000001100",
522 => "0000000000001100",
523 => "0000000000001100",
524 => "0000000000001100",
525 => "0000000000001100",
526 => "0000000000001100",
527 => "0000000000001100",
528 => "0000000000001100",
529 => "0000000000001100",
530 => "0000000000001100",
531 => "0000000000001100",
532 => "0000000000001100",
533 => "0000000000001100",
534 => "0000000000001100",
535 => "0000000000001100",
536 => "0000000000001100",
537 => "0000000000001100",
538 => "0000000000001100",
539 => "0000000000001100",
540 => "0000000000001100",
541 => "0000000000001100",
542 => "0000000000001100",
543 => "0000000000001100",
544 => "0000000000001100",
545 => "0000000000001100",
546 => "0000000000001100",
547 => "0000000000001100",
548 => "0000000000001100",
549 => "0000000000001100",
550 => "0000000000001100",
551 => "0000000000001100",
552 => "0000000000001100",
553 => "0000000000001100",
554 => "0000000000001100",
555 => "0000000000001100",
556 => "0000000000001100",
557 => "0000000000001100",
558 => "0000000000001100",
559 => "0000000000001100",
560 => "0000000000001100",
561 => "0000000000001100",
562 => "0000000000001100",
563 => "0000000000001100",
564 => "0000000000001100",
565 => "0000000000001100",
566 => "0000000000001100",
567 => "0000000000001100",
568 => "0000000000001100",
569 => "0000000000001100",
570 => "0000000000001100",
571 => "0000000000001100",
572 => "0000000000001100",
573 => "0000000000001100",
574 => "0000000000001100",
575 => "0000000000001100",
576 => "0000000000001100",
577 => "0000000000001100",
578 => "0000000000001100",
579 => "0000000000001100",
580 => "0000000000001100",
581 => "0000000000001100",
582 => "0000000000001100",
583 => "0000000000001100",
584 => "0000000000001100",
585 => "0000000000001100",
586 => "0000000000001100",
587 => "0000000000001100",
588 => "0000000000001100",
589 => "0000000000001100",
590 => "0000000000001100",
591 => "0000000000001100",
592 => "0000000000001100",
593 => "0000000000001100",
594 => "0000000000001100",
595 => "0000000000001100",
596 => "0000000000001100",
597 => "0000000000001100",
598 => "0000000000001100",
599 => "0000000000001100",
600 => "0000000000001100",
601 => "0000000000001100",
602 => "0000000000001100",
603 => "0000000000001100",
604 => "0000000000001100",
605 => "0000000000001100",
606 => "0000000000001100",
607 => "0000000000001100",
608 => "0000000000001100",
609 => "0000000000001100",
610 => "0000000000001100",
611 => "0000000000001100",
612 => "0000000000001100",
613 => "0000000000001100",
614 => "0000000000001100",
615 => "0000000000001100",
616 => "0000000000001100",
617 => "0000000000001100",
618 => "0000000000001100",
619 => "0000000000001100",
620 => "0000000000001100",
621 => "0000000000001100",
622 => "0000000000001100",
623 => "0000000000001100",
624 => "0000000000001100",
625 => "0000000000001100",
626 => "0000000000001100",
627 => "0000000000001100",
628 => "0000000000001100",
629 => "0000000000001100",
630 => "0000000000001100",
631 => "0000000000001100",
632 => "0000000000001100",
633 => "0000000000001100",
634 => "0000000000001100",
635 => "0000000000001100",
636 => "0000000000001100",
637 => "0000000000001100",
638 => "0000000000001100",
639 => "0000000000001100",
640 => "0000000000001100",
641 => "0000000000001100",
642 => "0000000000001100",
643 => "0000000000001100",
644 => "0000000000001100",
645 => "0000000000001100",
646 => "0000000000001100",
647 => "0000000000001100",
648 => "0000000000001100",
649 => "0000000000001100",
650 => "0000000000001100",
651 => "0000000000001100",
652 => "0000000000001100",
653 => "0000000000001100",
654 => "0000000000001100",
655 => "0000000000001100",
656 => "0000000000001100",
657 => "0000000000001100",
658 => "0000000000001100",
659 => "0000000000001100",
660 => "0000000000001100",
661 => "0000000000001100",
662 => "0000000000001100",
663 => "0000000000001100",
664 => "0000000000001100",
665 => "0000000000001100",
666 => "0000000000001100",
667 => "0000000000001100",
668 => "0000000000001100",
669 => "0000000000001100",
670 => "0000000000001100",
671 => "0000000000001100",
672 => "0000000000001100",
673 => "0000000000001100",
674 => "0000000000001100",
675 => "0000000000001100",
676 => "0000000000001100",
677 => "0000000000001100",
678 => "0000000000001100",
679 => "0000000000001100",
680 => "0000000000001100",
681 => "0000000000001100",
682 => "0000000000001100",
683 => "0000000000001100",
684 => "0000000000001100",
685 => "0000000000001100",
686 => "0000000000001100",
687 => "0000000000001100",
688 => "0000000000001101",
689 => "0000000000001101",
690 => "0000000000001101",
691 => "0000000000001101",
692 => "0000000000001101",
693 => "0000000000001101",
694 => "0000000000001101",
695 => "0000000000001101",
696 => "0000000000001101",
697 => "0000000000001101",
698 => "0000000000001101",
699 => "0000000000001101",
700 => "0000000000001101",
701 => "0000000000001101",
702 => "0000000000001101",
703 => "0000000000001101",
704 => "0000000000001101",
705 => "0000000000001101",
706 => "0000000000001101",
707 => "0000000000001101",
708 => "0000000000001101",
709 => "0000000000001101",
710 => "0000000000001101",
711 => "0000000000001101",
712 => "0000000000001101",
713 => "0000000000001101",
714 => "0000000000001101",
715 => "0000000000001101",
716 => "0000000000001101",
717 => "0000000000001101",
718 => "0000000000001101",
719 => "0000000000001101",
720 => "0000000000001101",
721 => "0000000000001101",
722 => "0000000000001101",
723 => "0000000000001101",
724 => "0000000000001101",
725 => "0000000000001101",
726 => "0000000000001101",
727 => "0000000000001101",
728 => "0000000000001101",
729 => "0000000000001101",
730 => "0000000000001101",
731 => "0000000000001101",
732 => "0000000000001101",
733 => "0000000000001101",
734 => "0000000000001101",
735 => "0000000000001101",
736 => "0000000000001101",
737 => "0000000000001101",
738 => "0000000000001101",
739 => "0000000000001101",
740 => "0000000000001101",
741 => "0000000000001101",
742 => "0000000000001101",
743 => "0000000000001101",
744 => "0000000000001101",
745 => "0000000000001101",
746 => "0000000000001101",
747 => "0000000000001101",
748 => "0000000000001101",
749 => "0000000000001101",
750 => "0000000000001101",
751 => "0000000000001101",
752 => "0000000000001101",
753 => "0000000000001101",
754 => "0000000000001101",
755 => "0000000000001101",
756 => "0000000000001101",
757 => "0000000000001101",
758 => "0000000000001101",
759 => "0000000000001101",
760 => "0000000000001101",
761 => "0000000000001101",
762 => "0000000000001101",
763 => "0000000000001101",
764 => "0000000000001101",
765 => "0000000000001101",
766 => "0000000000001101",
767 => "0000000000001101",
768 => "0000000000001101",
769 => "0000000000001101",
770 => "0000000000001101",
771 => "0000000000001101",
772 => "0000000000001101",
773 => "0000000000001101",
774 => "0000000000001101",
775 => "0000000000001101",
776 => "0000000000001101",
777 => "0000000000001101",
778 => "0000000000001101",
779 => "0000000000001101",
780 => "0000000000001101",
781 => "0000000000001101",
782 => "0000000000001101",
783 => "0000000000001101",
784 => "0000000000001101",
785 => "0000000000001101",
786 => "0000000000001101",
787 => "0000000000001101",
788 => "0000000000001101",
789 => "0000000000001101",
790 => "0000000000001101",
791 => "0000000000001101",
792 => "0000000000001101",
793 => "0000000000001101",
794 => "0000000000001101",
795 => "0000000000001101",
796 => "0000000000001101",
797 => "0000000000001101",
798 => "0000000000001101",
799 => "0000000000001101",
800 => "0000000000001101",
801 => "0000000000001101",
802 => "0000000000001101",
803 => "0000000000001101",
804 => "0000000000001101",
805 => "0000000000001101",
806 => "0000000000001101",
807 => "0000000000001101",
808 => "0000000000001101",
809 => "0000000000001101",
810 => "0000000000001101",
811 => "0000000000001101",
812 => "0000000000001101",
813 => "0000000000001101",
814 => "0000000000001101",
815 => "0000000000001101",
816 => "0000000000001101",
817 => "0000000000001101",
818 => "0000000000001101",
819 => "0000000000001101",
820 => "0000000000001101",
821 => "0000000000001101",
822 => "0000000000001101",
823 => "0000000000001101",
824 => "0000000000001101",
825 => "0000000000001101",
826 => "0000000000001101",
827 => "0000000000001101",
828 => "0000000000001101",
829 => "0000000000001101",
830 => "0000000000001101",
831 => "0000000000001101",
832 => "0000000000001101",
833 => "0000000000001101",
834 => "0000000000001101",
835 => "0000000000001101",
836 => "0000000000001101",
837 => "0000000000001101",
838 => "0000000000001101",
839 => "0000000000001101",
840 => "0000000000001101",
841 => "0000000000001101",
842 => "0000000000001101",
843 => "0000000000001101",
844 => "0000000000001101",
845 => "0000000000001101",
846 => "0000000000001101",
847 => "0000000000001101",
848 => "0000000000001101",
849 => "0000000000001101",
850 => "0000000000001101",
851 => "0000000000001101",
852 => "0000000000001101",
853 => "0000000000001101",
854 => "0000000000001101",
855 => "0000000000001101",
856 => "0000000000001101",
857 => "0000000000001101",
858 => "0000000000001101",
859 => "0000000000001101",
860 => "0000000000001101",
861 => "0000000000001101",
862 => "0000000000001101",
863 => "0000000000001101",
864 => "0000000000001101",
865 => "0000000000001101",
866 => "0000000000001101",
867 => "0000000000001101",
868 => "0000000000001101",
869 => "0000000000001101",
870 => "0000000000001101",
871 => "0000000000001101",
872 => "0000000000001101",
873 => "0000000000001101",
874 => "0000000000001101",
875 => "0000000000001101",
876 => "0000000000001101",
877 => "0000000000001101",
878 => "0000000000001101",
879 => "0000000000001101",
880 => "0000000000001101",
881 => "0000000000001101",
882 => "0000000000001101",
883 => "0000000000001101",
884 => "0000000000001101",
885 => "0000000000001101",
886 => "0000000000001101",
887 => "0000000000001101",
888 => "0000000000001101",
889 => "0000000000001101",
890 => "0000000000001101",
891 => "0000000000001101",
892 => "0000000000001101",
893 => "0000000000001101",
894 => "0000000000001101",
895 => "0000000000001101",
896 => "0000000000001101",
897 => "0000000000001101",
898 => "0000000000001101",
899 => "0000000000001101",
900 => "0000000000001101",
901 => "0000000000001101",
902 => "0000000000001101",
903 => "0000000000001101",
904 => "0000000000001101",
905 => "0000000000001101",
906 => "0000000000001101",
907 => "0000000000001101",
908 => "0000000000001101",
909 => "0000000000001101",
910 => "0000000000001101",
911 => "0000000000001101",
912 => "0000000000001101",
913 => "0000000000001101",
914 => "0000000000001101",
915 => "0000000000001101",
916 => "0000000000001101",
917 => "0000000000001101",
918 => "0000000000001101",
919 => "0000000000001101",
920 => "0000000000001101",
921 => "0000000000001101",
922 => "0000000000001101",
923 => "0000000000001101",
924 => "0000000000001101",
925 => "0000000000001101",
926 => "0000000000001101",
927 => "0000000000001101",
928 => "0000000000001101",
929 => "0000000000001101",
930 => "0000000000001101",
931 => "0000000000001101",
932 => "0000000000001101",
933 => "0000000000001101",
934 => "0000000000001101",
935 => "0000000000001101",
936 => "0000000000001101",
937 => "0000000000001101",
938 => "0000000000001101",
939 => "0000000000001101",
940 => "0000000000001101",
941 => "0000000000001101",
942 => "0000000000001101",
943 => "0000000000001101",
944 => "0000000000001101",
945 => "0000000000001101",
946 => "0000000000001101",
947 => "0000000000001101",
948 => "0000000000001101",
949 => "0000000000001101",
950 => "0000000000001101",
951 => "0000000000001101",
952 => "0000000000001101",
953 => "0000000000001101",
954 => "0000000000001101",
955 => "0000000000001101",
956 => "0000000000001101",
957 => "0000000000001101",
958 => "0000000000001101",
959 => "0000000000001101",
960 => "0000000000001101",
961 => "0000000000001101",
962 => "0000000000001101",
963 => "0000000000001101",
964 => "0000000000001101",
965 => "0000000000001101",
966 => "0000000000001101",
967 => "0000000000001101",
968 => "0000000000001101",
969 => "0000000000001101",
970 => "0000000000001101",
971 => "0000000000001101",
972 => "0000000000001101",
973 => "0000000000001101",
974 => "0000000000001101",
975 => "0000000000001101",
976 => "0000000000001101",
977 => "0000000000001101",
978 => "0000000000001101",
979 => "0000000000001101",
980 => "0000000000001101",
981 => "0000000000001101",
982 => "0000000000001101",
983 => "0000000000001101",
984 => "0000000000001101",
985 => "0000000000001101",
986 => "0000000000001101",
987 => "0000000000001101",
988 => "0000000000001101",
989 => "0000000000001101",
990 => "0000000000001101",
991 => "0000000000001101",
992 => "0000000000001110",
993 => "0000000000001110",
994 => "0000000000001110",
995 => "0000000000001110",
996 => "0000000000001110",
997 => "0000000000001110",
998 => "0000000000001110",
999 => "0000000000001110",
1000 => "0000000000001110",
1001 => "0000000000001110",
1002 => "0000000000001110",
1003 => "0000000000001110",
1004 => "0000000000001110",
1005 => "0000000000001110",
1006 => "0000000000001110",
1007 => "0000000000001110",
1008 => "0000000000001110",
1009 => "0000000000001110",
1010 => "0000000000001110",
1011 => "0000000000001110",
1012 => "0000000000001110",
1013 => "0000000000001110",
1014 => "0000000000001110",
1015 => "0000000000001110",
1016 => "0000000000001110",
1017 => "0000000000001110",
1018 => "0000000000001110",
1019 => "0000000000001110",
1020 => "0000000000001110",
1021 => "0000000000001110",
1022 => "0000000000001110",
1023 => "0000000000001110",
1024 => "0000000000001110",
1025 => "0000000000001110",
1026 => "0000000000001110",
1027 => "0000000000001110",
1028 => "0000000000001110",
1029 => "0000000000001110",
1030 => "0000000000001110",
1031 => "0000000000001110",
1032 => "0000000000001110",
1033 => "0000000000001110",
1034 => "0000000000001110",
1035 => "0000000000001110",
1036 => "0000000000001110",
1037 => "0000000000001110",
1038 => "0000000000001110",
1039 => "0000000000001110",
1040 => "0000000000001110",
1041 => "0000000000001110",
1042 => "0000000000001110",
1043 => "0000000000001110",
1044 => "0000000000001110",
1045 => "0000000000001110",
1046 => "0000000000001110",
1047 => "0000000000001110",
1048 => "0000000000001110",
1049 => "0000000000001110",
1050 => "0000000000001110",
1051 => "0000000000001110",
1052 => "0000000000001110",
1053 => "0000000000001110",
1054 => "0000000000001110",
1055 => "0000000000001110",
1056 => "0000000000001110",
1057 => "0000000000001110",
1058 => "0000000000001110",
1059 => "0000000000001110",
1060 => "0000000000001110",
1061 => "0000000000001110",
1062 => "0000000000001110",
1063 => "0000000000001110",
1064 => "0000000000001110",
1065 => "0000000000001110",
1066 => "0000000000001110",
1067 => "0000000000001110",
1068 => "0000000000001110",
1069 => "0000000000001110",
1070 => "0000000000001110",
1071 => "0000000000001110",
1072 => "0000000000001110",
1073 => "0000000000001110",
1074 => "0000000000001110",
1075 => "0000000000001110",
1076 => "0000000000001110",
1077 => "0000000000001110",
1078 => "0000000000001110",
1079 => "0000000000001110",
1080 => "0000000000001110",
1081 => "0000000000001110",
1082 => "0000000000001110",
1083 => "0000000000001110",
1084 => "0000000000001110",
1085 => "0000000000001110",
1086 => "0000000000001110",
1087 => "0000000000001110",
1088 => "0000000000001110",
1089 => "0000000000001110",
1090 => "0000000000001110",
1091 => "0000000000001110",
1092 => "0000000000001110",
1093 => "0000000000001110",
1094 => "0000000000001110",
1095 => "0000000000001110",
1096 => "0000000000001110",
1097 => "0000000000001110",
1098 => "0000000000001110",
1099 => "0000000000001110",
1100 => "0000000000001110",
1101 => "0000000000001110",
1102 => "0000000000001110",
1103 => "0000000000001110",
1104 => "0000000000001110",
1105 => "0000000000001110",
1106 => "0000000000001110",
1107 => "0000000000001110",
1108 => "0000000000001110",
1109 => "0000000000001110",
1110 => "0000000000001110",
1111 => "0000000000001110",
1112 => "0000000000001110",
1113 => "0000000000001110",
1114 => "0000000000001110",
1115 => "0000000000001110",
1116 => "0000000000001110",
1117 => "0000000000001110",
1118 => "0000000000001110",
1119 => "0000000000001110",
1120 => "0000000000001110",
1121 => "0000000000001110",
1122 => "0000000000001110",
1123 => "0000000000001110",
1124 => "0000000000001110",
1125 => "0000000000001110",
1126 => "0000000000001110",
1127 => "0000000000001110",
1128 => "0000000000001110",
1129 => "0000000000001110",
1130 => "0000000000001110",
1131 => "0000000000001110",
1132 => "0000000000001110",
1133 => "0000000000001110",
1134 => "0000000000001110",
1135 => "0000000000001110",
1136 => "0000000000001110",
1137 => "0000000000001110",
1138 => "0000000000001110",
1139 => "0000000000001110",
1140 => "0000000000001110",
1141 => "0000000000001110",
1142 => "0000000000001110",
1143 => "0000000000001110",
1144 => "0000000000001110",
1145 => "0000000000001110",
1146 => "0000000000001110",
1147 => "0000000000001110",
1148 => "0000000000001110",
1149 => "0000000000001110",
1150 => "0000000000001110",
1151 => "0000000000001110",
1152 => "0000000000001110",
1153 => "0000000000001110",
1154 => "0000000000001110",
1155 => "0000000000001110",
1156 => "0000000000001110",
1157 => "0000000000001110",
1158 => "0000000000001110",
1159 => "0000000000001110",
1160 => "0000000000001110",
1161 => "0000000000001110",
1162 => "0000000000001110",
1163 => "0000000000001110",
1164 => "0000000000001110",
1165 => "0000000000001110",
1166 => "0000000000001110",
1167 => "0000000000001110",
1168 => "0000000000001110",
1169 => "0000000000001110",
1170 => "0000000000001110",
1171 => "0000000000001110",
1172 => "0000000000001110",
1173 => "0000000000001110",
1174 => "0000000000001110",
1175 => "0000000000001110",
1176 => "0000000000001110",
1177 => "0000000000001110",
1178 => "0000000000001110",
1179 => "0000000000001110",
1180 => "0000000000001110",
1181 => "0000000000001110",
1182 => "0000000000001110",
1183 => "0000000000001110",
1184 => "0000000000001110",
1185 => "0000000000001110",
1186 => "0000000000001110",
1187 => "0000000000001110",
1188 => "0000000000001110",
1189 => "0000000000001110",
1190 => "0000000000001110",
1191 => "0000000000001110",
1192 => "0000000000001110",
1193 => "0000000000001110",
1194 => "0000000000001110",
1195 => "0000000000001110",
1196 => "0000000000001110",
1197 => "0000000000001110",
1198 => "0000000000001110",
1199 => "0000000000001110",
1200 => "0000000000001110",
1201 => "0000000000001110",
1202 => "0000000000001110",
1203 => "0000000000001110",
1204 => "0000000000001110",
1205 => "0000000000001110",
1206 => "0000000000001110",
1207 => "0000000000001110",
1208 => "0000000000001110",
1209 => "0000000000001110",
1210 => "0000000000001110",
1211 => "0000000000001110",
1212 => "0000000000001110",
1213 => "0000000000001110",
1214 => "0000000000001110",
1215 => "0000000000001110",
1216 => "0000000000001110",
1217 => "0000000000001110",
1218 => "0000000000001110",
1219 => "0000000000001110",
1220 => "0000000000001110",
1221 => "0000000000001110",
1222 => "0000000000001110",
1223 => "0000000000001110",
1224 => "0000000000001110",
1225 => "0000000000001110",
1226 => "0000000000001110",
1227 => "0000000000001110",
1228 => "0000000000001110",
1229 => "0000000000001110",
1230 => "0000000000001110",
1231 => "0000000000001110",
1232 => "0000000000001110",
1233 => "0000000000001110",
1234 => "0000000000001110",
1235 => "0000000000001110",
1236 => "0000000000001110",
1237 => "0000000000001110",
1238 => "0000000000001110",
1239 => "0000000000001110",
1240 => "0000000000001110",
1241 => "0000000000001110",
1242 => "0000000000001110",
1243 => "0000000000001110",
1244 => "0000000000001110",
1245 => "0000000000001110",
1246 => "0000000000001110",
1247 => "0000000000001110",
1248 => "0000000000001110",
1249 => "0000000000001110",
1250 => "0000000000001110",
1251 => "0000000000001110",
1252 => "0000000000001110",
1253 => "0000000000001110",
1254 => "0000000000001110",
1255 => "0000000000001110",
1256 => "0000000000001110",
1257 => "0000000000001110",
1258 => "0000000000001110",
1259 => "0000000000001110",
1260 => "0000000000001110",
1261 => "0000000000001110",
1262 => "0000000000001110",
1263 => "0000000000001110",
1264 => "0000000000001110",
1265 => "0000000000001110",
1266 => "0000000000001110",
1267 => "0000000000001110",
1268 => "0000000000001110",
1269 => "0000000000001110",
1270 => "0000000000001110",
1271 => "0000000000001110",
1272 => "0000000000001110",
1273 => "0000000000001110",
1274 => "0000000000001111",
1275 => "0000000000001111",
1276 => "0000000000001111",
1277 => "0000000000001111",
1278 => "0000000000001111",
1279 => "0000000000001111",
1280 => "0000000000001111",
1281 => "0000000000001111",
1282 => "0000000000001111",
1283 => "0000000000001111",
1284 => "0000000000001111",
1285 => "0000000000001111",
1286 => "0000000000001111",
1287 => "0000000000001111",
1288 => "0000000000001111",
1289 => "0000000000001111",
1290 => "0000000000001111",
1291 => "0000000000001111",
1292 => "0000000000001111",
1293 => "0000000000001111",
1294 => "0000000000001111",
1295 => "0000000000001111",
1296 => "0000000000001111",
1297 => "0000000000001111",
1298 => "0000000000001111",
1299 => "0000000000001111",
1300 => "0000000000001111",
1301 => "0000000000001111",
1302 => "0000000000001111",
1303 => "0000000000001111",
1304 => "0000000000001111",
1305 => "0000000000001111",
1306 => "0000000000001111",
1307 => "0000000000001111",
1308 => "0000000000001111",
1309 => "0000000000001111",
1310 => "0000000000001111",
1311 => "0000000000001111",
1312 => "0000000000001111",
1313 => "0000000000001111",
1314 => "0000000000001111",
1315 => "0000000000001111",
1316 => "0000000000001111",
1317 => "0000000000001111",
1318 => "0000000000001111",
1319 => "0000000000001111",
1320 => "0000000000001111",
1321 => "0000000000001111",
1322 => "0000000000001111",
1323 => "0000000000001111",
1324 => "0000000000001111",
1325 => "0000000000001111",
1326 => "0000000000001111",
1327 => "0000000000001111",
1328 => "0000000000001111",
1329 => "0000000000001111",
1330 => "0000000000001111",
1331 => "0000000000001111",
1332 => "0000000000001111",
1333 => "0000000000001111",
1334 => "0000000000001111",
1335 => "0000000000001111",
1336 => "0000000000001111",
1337 => "0000000000001111",
1338 => "0000000000001111",
1339 => "0000000000001111",
1340 => "0000000000001111",
1341 => "0000000000001111",
1342 => "0000000000001111",
1343 => "0000000000001111",
1344 => "0000000000001111",
1345 => "0000000000001111",
1346 => "0000000000001111",
1347 => "0000000000001111",
1348 => "0000000000001111",
1349 => "0000000000001111",
1350 => "0000000000001111",
1351 => "0000000000001111",
1352 => "0000000000001111",
1353 => "0000000000001111",
1354 => "0000000000001111",
1355 => "0000000000001111",
1356 => "0000000000001111",
1357 => "0000000000001111",
1358 => "0000000000001111",
1359 => "0000000000001111",
1360 => "0000000000001111",
1361 => "0000000000001111",
1362 => "0000000000001111",
1363 => "0000000000001111",
1364 => "0000000000001111",
1365 => "0000000000001111",
1366 => "0000000000001111",
1367 => "0000000000001111",
1368 => "0000000000001111",
1369 => "0000000000001111",
1370 => "0000000000001111",
1371 => "0000000000001111",
1372 => "0000000000001111",
1373 => "0000000000001111",
1374 => "0000000000001111",
1375 => "0000000000001111",
1376 => "0000000000001111",
1377 => "0000000000001111",
1378 => "0000000000001111",
1379 => "0000000000001111",
1380 => "0000000000001111",
1381 => "0000000000001111",
1382 => "0000000000001111",
1383 => "0000000000001111",
1384 => "0000000000001111",
1385 => "0000000000001111",
1386 => "0000000000001111",
1387 => "0000000000001111",
1388 => "0000000000001111",
1389 => "0000000000001111",
1390 => "0000000000001111",
1391 => "0000000000001111",
1392 => "0000000000001111",
1393 => "0000000000001111",
1394 => "0000000000001111",
1395 => "0000000000001111",
1396 => "0000000000001111",
1397 => "0000000000001111",
1398 => "0000000000001111",
1399 => "0000000000001111",
1400 => "0000000000001111",
1401 => "0000000000001111",
1402 => "0000000000001111",
1403 => "0000000000001111",
1404 => "0000000000001111",
1405 => "0000000000001111",
1406 => "0000000000001111",
1407 => "0000000000001111",
1408 => "0000000000001111",
1409 => "0000000000001111",
1410 => "0000000000001111",
1411 => "0000000000001111",
1412 => "0000000000001111",
1413 => "0000000000001111",
1414 => "0000000000001111",
1415 => "0000000000001111",
1416 => "0000000000001111",
1417 => "0000000000001111",
1418 => "0000000000001111",
1419 => "0000000000001111",
1420 => "0000000000001111",
1421 => "0000000000001111",
1422 => "0000000000001111",
1423 => "0000000000001111",
1424 => "0000000000001111",
1425 => "0000000000001111",
1426 => "0000000000001111",
1427 => "0000000000001111",
1428 => "0000000000001111",
1429 => "0000000000001111",
1430 => "0000000000001111",
1431 => "0000000000001111",
1432 => "0000000000001111",
1433 => "0000000000001111",
1434 => "0000000000001111",
1435 => "0000000000001111",
1436 => "0000000000001111",
1437 => "0000000000001111",
1438 => "0000000000001111",
1439 => "0000000000001111",
1440 => "0000000000001111",
1441 => "0000000000001111",
1442 => "0000000000001111",
1443 => "0000000000001111",
1444 => "0000000000001111",
1445 => "0000000000001111",
1446 => "0000000000001111",
1447 => "0000000000001111",
1448 => "0000000000001111",
1449 => "0000000000001111",
1450 => "0000000000001111",
1451 => "0000000000001111",
1452 => "0000000000001111",
1453 => "0000000000001111",
1454 => "0000000000001111",
1455 => "0000000000001111",
1456 => "0000000000001111",
1457 => "0000000000001111",
1458 => "0000000000001111",
1459 => "0000000000001111",
1460 => "0000000000001111",
1461 => "0000000000001111",
1462 => "0000000000001111",
1463 => "0000000000001111",
1464 => "0000000000001111",
1465 => "0000000000001111",
1466 => "0000000000001111",
1467 => "0000000000001111",
1468 => "0000000000001111",
1469 => "0000000000001111",
1470 => "0000000000001111",
1471 => "0000000000001111",
1472 => "0000000000001111",
1473 => "0000000000001111",
1474 => "0000000000001111",
1475 => "0000000000001111",
1476 => "0000000000001111",
1477 => "0000000000001111",
1478 => "0000000000001111",
1479 => "0000000000001111",
1480 => "0000000000001111",
1481 => "0000000000001111",
1482 => "0000000000001111",
1483 => "0000000000001111",
1484 => "0000000000001111",
1485 => "0000000000001111",
1486 => "0000000000001111",
1487 => "0000000000001111",
1488 => "0000000000001111",
1489 => "0000000000001111",
1490 => "0000000000001111",
1491 => "0000000000001111",
1492 => "0000000000001111",
1493 => "0000000000001111",
1494 => "0000000000001111",
1495 => "0000000000001111",
1496 => "0000000000001111",
1497 => "0000000000001111",
1498 => "0000000000001111",
1499 => "0000000000001111",
1500 => "0000000000001111",
1501 => "0000000000001111",
1502 => "0000000000001111",
1503 => "0000000000001111",
1504 => "0000000000001111",
1505 => "0000000000001111",
1506 => "0000000000001111",
1507 => "0000000000001111",
1508 => "0000000000001111",
1509 => "0000000000001111",
1510 => "0000000000001111",
1511 => "0000000000001111",
1512 => "0000000000001111",
1513 => "0000000000001111",
1514 => "0000000000001111",
1515 => "0000000000001111",
1516 => "0000000000001111",
1517 => "0000000000001111",
1518 => "0000000000001111",
1519 => "0000000000001111",
1520 => "0000000000001111",
1521 => "0000000000001111",
1522 => "0000000000001111",
1523 => "0000000000001111",
1524 => "0000000000001111",
1525 => "0000000000001111",
1526 => "0000000000001111",
1527 => "0000000000001111",
1528 => "0000000000001111",
1529 => "0000000000001111",
1530 => "0000000000001111",
1531 => "0000000000001111",
1532 => "0000000000001111",
1533 => "0000000000001111",
1534 => "0000000000001111",
1535 => "0000000000001111",
1536 => "0000000000001111",
1537 => "0000000000001111",
1538 => "0000000000001111",
1539 => "0000000000010000",
1540 => "0000000000010000",
1541 => "0000000000010000",
1542 => "0000000000010000",
1543 => "0000000000010000",
1544 => "0000000000010000",
1545 => "0000000000010000",
1546 => "0000000000010000",
1547 => "0000000000010000",
1548 => "0000000000010000",
1549 => "0000000000010000",
1550 => "0000000000010000",
1551 => "0000000000010000",
1552 => "0000000000010000",
1553 => "0000000000010000",
1554 => "0000000000010000",
1555 => "0000000000010000",
1556 => "0000000000010000",
1557 => "0000000000010000",
1558 => "0000000000010000",
1559 => "0000000000010000",
1560 => "0000000000010000",
1561 => "0000000000010000",
1562 => "0000000000010000",
1563 => "0000000000010000",
1564 => "0000000000010000",
1565 => "0000000000010000",
1566 => "0000000000010000",
1567 => "0000000000010000",
1568 => "0000000000010000",
1569 => "0000000000010000",
1570 => "0000000000010000",
1571 => "0000000000010000",
1572 => "0000000000010000",
1573 => "0000000000010000",
1574 => "0000000000010000",
1575 => "0000000000010000",
1576 => "0000000000010000",
1577 => "0000000000010000",
1578 => "0000000000010000",
1579 => "0000000000010000",
1580 => "0000000000010000",
1581 => "0000000000010000",
1582 => "0000000000010000",
1583 => "0000000000010000",
1584 => "0000000000010000",
1585 => "0000000000010000",
1586 => "0000000000010000",
1587 => "0000000000010000",
1588 => "0000000000010000",
1589 => "0000000000010000",
1590 => "0000000000010000",
1591 => "0000000000010000",
1592 => "0000000000010000",
1593 => "0000000000010000",
1594 => "0000000000010000",
1595 => "0000000000010000",
1596 => "0000000000010000",
1597 => "0000000000010000",
1598 => "0000000000010000",
1599 => "0000000000010000",
1600 => "0000000000010000",
1601 => "0000000000010000",
1602 => "0000000000010000",
1603 => "0000000000010000",
1604 => "0000000000010000",
1605 => "0000000000010000",
1606 => "0000000000010000",
1607 => "0000000000010000",
1608 => "0000000000010000",
1609 => "0000000000010000",
1610 => "0000000000010000",
1611 => "0000000000010000",
1612 => "0000000000010000",
1613 => "0000000000010000",
1614 => "0000000000010000",
1615 => "0000000000010000",
1616 => "0000000000010000",
1617 => "0000000000010000",
1618 => "0000000000010000",
1619 => "0000000000010000",
1620 => "0000000000010000",
1621 => "0000000000010000",
1622 => "0000000000010000",
1623 => "0000000000010000",
1624 => "0000000000010000",
1625 => "0000000000010000",
1626 => "0000000000010000",
1627 => "0000000000010000",
1628 => "0000000000010000",
1629 => "0000000000010000",
1630 => "0000000000010000",
1631 => "0000000000010000",
1632 => "0000000000010000",
1633 => "0000000000010000",
1634 => "0000000000010000",
1635 => "0000000000010000",
1636 => "0000000000010000",
1637 => "0000000000010000",
1638 => "0000000000010000",
1639 => "0000000000010000",
1640 => "0000000000010000",
1641 => "0000000000010000",
1642 => "0000000000010000",
1643 => "0000000000010000",
1644 => "0000000000010000",
1645 => "0000000000010000",
1646 => "0000000000010000",
1647 => "0000000000010000",
1648 => "0000000000010000",
1649 => "0000000000010000",
1650 => "0000000000010000",
1651 => "0000000000010000",
1652 => "0000000000010000",
1653 => "0000000000010000",
1654 => "0000000000010000",
1655 => "0000000000010000",
1656 => "0000000000010000",
1657 => "0000000000010000",
1658 => "0000000000010000",
1659 => "0000000000010000",
1660 => "0000000000010000",
1661 => "0000000000010000",
1662 => "0000000000010000",
1663 => "0000000000010000",
1664 => "0000000000010000",
1665 => "0000000000010000",
1666 => "0000000000010000",
1667 => "0000000000010000",
1668 => "0000000000010000",
1669 => "0000000000010000",
1670 => "0000000000010000",
1671 => "0000000000010000",
1672 => "0000000000010000",
1673 => "0000000000010000",
1674 => "0000000000010000",
1675 => "0000000000010000",
1676 => "0000000000010000",
1677 => "0000000000010000",
1678 => "0000000000010000",
1679 => "0000000000010000",
1680 => "0000000000010000",
1681 => "0000000000010000",
1682 => "0000000000010000",
1683 => "0000000000010000",
1684 => "0000000000010000",
1685 => "0000000000010000",
1686 => "0000000000010000",
1687 => "0000000000010000",
1688 => "0000000000010000",
1689 => "0000000000010000",
1690 => "0000000000010000",
1691 => "0000000000010000",
1692 => "0000000000010000",
1693 => "0000000000010000",
1694 => "0000000000010000",
1695 => "0000000000010000",
1696 => "0000000000010000",
1697 => "0000000000010000",
1698 => "0000000000010000",
1699 => "0000000000010000",
1700 => "0000000000010000",
1701 => "0000000000010000",
1702 => "0000000000010000",
1703 => "0000000000010000",
1704 => "0000000000010000",
1705 => "0000000000010000",
1706 => "0000000000010000",
1707 => "0000000000010000",
1708 => "0000000000010000",
1709 => "0000000000010000",
1710 => "0000000000010000",
1711 => "0000000000010000",
1712 => "0000000000010000",
1713 => "0000000000010000",
1714 => "0000000000010000",
1715 => "0000000000010000",
1716 => "0000000000010000",
1717 => "0000000000010000",
1718 => "0000000000010000",
1719 => "0000000000010000",
1720 => "0000000000010000",
1721 => "0000000000010000",
1722 => "0000000000010000",
1723 => "0000000000010000",
1724 => "0000000000010000",
1725 => "0000000000010000",
1726 => "0000000000010000",
1727 => "0000000000010000",
1728 => "0000000000010000",
1729 => "0000000000010000",
1730 => "0000000000010000",
1731 => "0000000000010000",
1732 => "0000000000010000",
1733 => "0000000000010000",
1734 => "0000000000010000",
1735 => "0000000000010000",
1736 => "0000000000010000",
1737 => "0000000000010000",
1738 => "0000000000010000",
1739 => "0000000000010000",
1740 => "0000000000010000",
1741 => "0000000000010000",
1742 => "0000000000010000",
1743 => "0000000000010000",
1744 => "0000000000010000",
1745 => "0000000000010000",
1746 => "0000000000010000",
1747 => "0000000000010000",
1748 => "0000000000010000",
1749 => "0000000000010000",
1750 => "0000000000010000",
1751 => "0000000000010000",
1752 => "0000000000010000",
1753 => "0000000000010000",
1754 => "0000000000010000",
1755 => "0000000000010000",
1756 => "0000000000010000",
1757 => "0000000000010000",
1758 => "0000000000010000",
1759 => "0000000000010000",
1760 => "0000000000010000",
1761 => "0000000000010000",
1762 => "0000000000010000",
1763 => "0000000000010000",
1764 => "0000000000010000",
1765 => "0000000000010000",
1766 => "0000000000010000",
1767 => "0000000000010000",
1768 => "0000000000010000",
1769 => "0000000000010000",
1770 => "0000000000010000",
1771 => "0000000000010000",
1772 => "0000000000010000",
1773 => "0000000000010000",
1774 => "0000000000010000",
1775 => "0000000000010000",
1776 => "0000000000010000",
1777 => "0000000000010000",
1778 => "0000000000010000",
1779 => "0000000000010000",
1780 => "0000000000010000",
1781 => "0000000000010000",
1782 => "0000000000010000",
1783 => "0000000000010000",
1784 => "0000000000010000",
1785 => "0000000000010000",
1786 => "0000000000010000",
1787 => "0000000000010001",
1788 => "0000000000010001",
1789 => "0000000000010001",
1790 => "0000000000010001",
1791 => "0000000000010001",
1792 => "0000000000010001",
1793 => "0000000000010001",
1794 => "0000000000010001",
1795 => "0000000000010001",
1796 => "0000000000010001",
1797 => "0000000000010001",
1798 => "0000000000010001",
1799 => "0000000000010001",
1800 => "0000000000010001",
1801 => "0000000000010001",
1802 => "0000000000010001",
1803 => "0000000000010001",
1804 => "0000000000010001",
1805 => "0000000000010001",
1806 => "0000000000010001",
1807 => "0000000000010001",
1808 => "0000000000010001",
1809 => "0000000000010001",
1810 => "0000000000010001",
1811 => "0000000000010001",
1812 => "0000000000010001",
1813 => "0000000000010001",
1814 => "0000000000010001",
1815 => "0000000000010001",
1816 => "0000000000010001",
1817 => "0000000000010001",
1818 => "0000000000010001",
1819 => "0000000000010001",
1820 => "0000000000010001",
1821 => "0000000000010001",
1822 => "0000000000010001",
1823 => "0000000000010001",
1824 => "0000000000010001",
1825 => "0000000000010001",
1826 => "0000000000010001",
1827 => "0000000000010001",
1828 => "0000000000010001",
1829 => "0000000000010001",
1830 => "0000000000010001",
1831 => "0000000000010001",
1832 => "0000000000010001",
1833 => "0000000000010001",
1834 => "0000000000010001",
1835 => "0000000000010001",
1836 => "0000000000010001",
1837 => "0000000000010001",
1838 => "0000000000010001",
1839 => "0000000000010001",
1840 => "0000000000010001",
1841 => "0000000000010001",
1842 => "0000000000010001",
1843 => "0000000000010001",
1844 => "0000000000010001",
1845 => "0000000000010001",
1846 => "0000000000010001",
1847 => "0000000000010001",
1848 => "0000000000010001",
1849 => "0000000000010001",
1850 => "0000000000010001",
1851 => "0000000000010001",
1852 => "0000000000010001",
1853 => "0000000000010001",
1854 => "0000000000010001",
1855 => "0000000000010001",
1856 => "0000000000010001",
1857 => "0000000000010001",
1858 => "0000000000010001",
1859 => "0000000000010001",
1860 => "0000000000010001",
1861 => "0000000000010001",
1862 => "0000000000010001",
1863 => "0000000000010001",
1864 => "0000000000010001",
1865 => "0000000000010001",
1866 => "0000000000010001",
1867 => "0000000000010001",
1868 => "0000000000010001",
1869 => "0000000000010001",
1870 => "0000000000010001",
1871 => "0000000000010001",
1872 => "0000000000010001",
1873 => "0000000000010001",
1874 => "0000000000010001",
1875 => "0000000000010001",
1876 => "0000000000010001",
1877 => "0000000000010001",
1878 => "0000000000010001",
1879 => "0000000000010001",
1880 => "0000000000010001",
1881 => "0000000000010001",
1882 => "0000000000010001",
1883 => "0000000000010001",
1884 => "0000000000010001",
1885 => "0000000000010001",
1886 => "0000000000010001",
1887 => "0000000000010001",
1888 => "0000000000010001",
1889 => "0000000000010001",
1890 => "0000000000010001",
1891 => "0000000000010001",
1892 => "0000000000010001",
1893 => "0000000000010001",
1894 => "0000000000010001",
1895 => "0000000000010001",
1896 => "0000000000010001",
1897 => "0000000000010001",
1898 => "0000000000010001",
1899 => "0000000000010001",
1900 => "0000000000010001",
1901 => "0000000000010001",
1902 => "0000000000010001",
1903 => "0000000000010001",
1904 => "0000000000010001",
1905 => "0000000000010001",
1906 => "0000000000010001",
1907 => "0000000000010001",
1908 => "0000000000010001",
1909 => "0000000000010001",
1910 => "0000000000010001",
1911 => "0000000000010001",
1912 => "0000000000010001",
1913 => "0000000000010001",
1914 => "0000000000010001",
1915 => "0000000000010001",
1916 => "0000000000010001",
1917 => "0000000000010001",
1918 => "0000000000010001",
1919 => "0000000000010001",
1920 => "0000000000010001",
1921 => "0000000000010001",
1922 => "0000000000010001",
1923 => "0000000000010001",
1924 => "0000000000010001",
1925 => "0000000000010001",
1926 => "0000000000010001",
1927 => "0000000000010001",
1928 => "0000000000010001",
1929 => "0000000000010001",
1930 => "0000000000010001",
1931 => "0000000000010001",
1932 => "0000000000010001",
1933 => "0000000000010001",
1934 => "0000000000010001",
1935 => "0000000000010001",
1936 => "0000000000010001",
1937 => "0000000000010001",
1938 => "0000000000010001",
1939 => "0000000000010001",
1940 => "0000000000010001",
1941 => "0000000000010001",
1942 => "0000000000010001",
1943 => "0000000000010001",
1944 => "0000000000010001",
1945 => "0000000000010001",
1946 => "0000000000010001",
1947 => "0000000000010001",
1948 => "0000000000010001",
1949 => "0000000000010001",
1950 => "0000000000010001",
1951 => "0000000000010001",
1952 => "0000000000010001",
1953 => "0000000000010001",
1954 => "0000000000010001",
1955 => "0000000000010001",
1956 => "0000000000010001",
1957 => "0000000000010001",
1958 => "0000000000010001",
1959 => "0000000000010001",
1960 => "0000000000010001",
1961 => "0000000000010001",
1962 => "0000000000010001",
1963 => "0000000000010001",
1964 => "0000000000010001",
1965 => "0000000000010001",
1966 => "0000000000010001",
1967 => "0000000000010001",
1968 => "0000000000010001",
1969 => "0000000000010001",
1970 => "0000000000010001",
1971 => "0000000000010001",
1972 => "0000000000010001",
1973 => "0000000000010001",
1974 => "0000000000010001",
1975 => "0000000000010001",
1976 => "0000000000010001",
1977 => "0000000000010001",
1978 => "0000000000010001",
1979 => "0000000000010001",
1980 => "0000000000010001",
1981 => "0000000000010001",
1982 => "0000000000010001",
1983 => "0000000000010001",
1984 => "0000000000010001",
1985 => "0000000000010001",
1986 => "0000000000010001",
1987 => "0000000000010001",
1988 => "0000000000010001",
1989 => "0000000000010001",
1990 => "0000000000010001",
1991 => "0000000000010001",
1992 => "0000000000010001",
1993 => "0000000000010001",
1994 => "0000000000010001",
1995 => "0000000000010001",
1996 => "0000000000010001",
1997 => "0000000000010001",
1998 => "0000000000010001",
1999 => "0000000000010001",
2000 => "0000000000010001",
2001 => "0000000000010001",
2002 => "0000000000010001",
2003 => "0000000000010001",
2004 => "0000000000010001",
2005 => "0000000000010001",
2006 => "0000000000010001",
2007 => "0000000000010001",
2008 => "0000000000010001",
2009 => "0000000000010001",
2010 => "0000000000010001",
2011 => "0000000000010001",
2012 => "0000000000010001",
2013 => "0000000000010001",
2014 => "0000000000010001",
2015 => "0000000000010001",
2016 => "0000000000010001",
2017 => "0000000000010001",
2018 => "0000000000010001",
2019 => "0000000000010001",
2020 => "0000000000010001",
2021 => "0000000000010010",
2022 => "0000000000010010",
2023 => "0000000000010010",
2024 => "0000000000010010",
2025 => "0000000000010010",
2026 => "0000000000010010",
2027 => "0000000000010010",
2028 => "0000000000010010",
2029 => "0000000000010010",
2030 => "0000000000010010",
2031 => "0000000000010010",
2032 => "0000000000010010",
2033 => "0000000000010010",
2034 => "0000000000010010",
2035 => "0000000000010010",
2036 => "0000000000010010",
2037 => "0000000000010010",
2038 => "0000000000010010",
2039 => "0000000000010010",
2040 => "0000000000010010",
2041 => "0000000000010010",
2042 => "0000000000010010",
2043 => "0000000000010010",
2044 => "0000000000010010",
2045 => "0000000000010010",
2046 => "0000000000010010",
2047 => "0000000000010010",
2048 => "0000000000010010",
2049 => "0000000000010010",
2050 => "0000000000010010",
2051 => "0000000000010010",
2052 => "0000000000010010",
2053 => "0000000000010010",
2054 => "0000000000010010",
2055 => "0000000000010010",
2056 => "0000000000010010",
2057 => "0000000000010010",
2058 => "0000000000010010",
2059 => "0000000000010010",
2060 => "0000000000010010",
2061 => "0000000000010010",
2062 => "0000000000010010",
2063 => "0000000000010010",
2064 => "0000000000010010",
2065 => "0000000000010010",
2066 => "0000000000010010",
2067 => "0000000000010010",
2068 => "0000000000010010",
2069 => "0000000000010010",
2070 => "0000000000010010",
2071 => "0000000000010010",
2072 => "0000000000010010",
2073 => "0000000000010010",
2074 => "0000000000010010",
2075 => "0000000000010010",
2076 => "0000000000010010",
2077 => "0000000000010010",
2078 => "0000000000010010",
2079 => "0000000000010010",
2080 => "0000000000010010",
2081 => "0000000000010010",
2082 => "0000000000010010",
2083 => "0000000000010010",
2084 => "0000000000010010",
2085 => "0000000000010010",
2086 => "0000000000010010",
2087 => "0000000000010010",
2088 => "0000000000010010",
2089 => "0000000000010010",
2090 => "0000000000010010",
2091 => "0000000000010010",
2092 => "0000000000010010",
2093 => "0000000000010010",
2094 => "0000000000010010",
2095 => "0000000000010010",
2096 => "0000000000010010",
2097 => "0000000000010010",
2098 => "0000000000010010",
2099 => "0000000000010010",
2100 => "0000000000010010",
2101 => "0000000000010010",
2102 => "0000000000010010",
2103 => "0000000000010010",
2104 => "0000000000010010",
2105 => "0000000000010010",
2106 => "0000000000010010",
2107 => "0000000000010010",
2108 => "0000000000010010",
2109 => "0000000000010010",
2110 => "0000000000010010",
2111 => "0000000000010010",
2112 => "0000000000010010",
2113 => "0000000000010010",
2114 => "0000000000010010",
2115 => "0000000000010010",
2116 => "0000000000010010",
2117 => "0000000000010010",
2118 => "0000000000010010",
2119 => "0000000000010010",
2120 => "0000000000010010",
2121 => "0000000000010010",
2122 => "0000000000010010",
2123 => "0000000000010010",
2124 => "0000000000010010",
2125 => "0000000000010010",
2126 => "0000000000010010",
2127 => "0000000000010010",
2128 => "0000000000010010",
2129 => "0000000000010010",
2130 => "0000000000010010",
2131 => "0000000000010010",
2132 => "0000000000010010",
2133 => "0000000000010010",
2134 => "0000000000010010",
2135 => "0000000000010010",
2136 => "0000000000010010",
2137 => "0000000000010010",
2138 => "0000000000010010",
2139 => "0000000000010010",
2140 => "0000000000010010",
2141 => "0000000000010010",
2142 => "0000000000010010",
2143 => "0000000000010010",
2144 => "0000000000010010",
2145 => "0000000000010010",
2146 => "0000000000010010",
2147 => "0000000000010010",
2148 => "0000000000010010",
2149 => "0000000000010010",
2150 => "0000000000010010",
2151 => "0000000000010010",
2152 => "0000000000010010",
2153 => "0000000000010010",
2154 => "0000000000010010",
2155 => "0000000000010010",
2156 => "0000000000010010",
2157 => "0000000000010010",
2158 => "0000000000010010",
2159 => "0000000000010010",
2160 => "0000000000010010",
2161 => "0000000000010010",
2162 => "0000000000010010",
2163 => "0000000000010010",
2164 => "0000000000010010",
2165 => "0000000000010010",
2166 => "0000000000010010",
2167 => "0000000000010010",
2168 => "0000000000010010",
2169 => "0000000000010010",
2170 => "0000000000010010",
2171 => "0000000000010010",
2172 => "0000000000010010",
2173 => "0000000000010010",
2174 => "0000000000010010",
2175 => "0000000000010010",
2176 => "0000000000010010",
2177 => "0000000000010010",
2178 => "0000000000010010",
2179 => "0000000000010010",
2180 => "0000000000010010",
2181 => "0000000000010010",
2182 => "0000000000010010",
2183 => "0000000000010010",
2184 => "0000000000010010",
2185 => "0000000000010010",
2186 => "0000000000010010",
2187 => "0000000000010010",
2188 => "0000000000010010",
2189 => "0000000000010010",
2190 => "0000000000010010",
2191 => "0000000000010010",
2192 => "0000000000010010",
2193 => "0000000000010010",
2194 => "0000000000010010",
2195 => "0000000000010010",
2196 => "0000000000010010",
2197 => "0000000000010010",
2198 => "0000000000010010",
2199 => "0000000000010010",
2200 => "0000000000010010",
2201 => "0000000000010010",
2202 => "0000000000010010",
2203 => "0000000000010010",
2204 => "0000000000010010",
2205 => "0000000000010010",
2206 => "0000000000010010",
2207 => "0000000000010010",
2208 => "0000000000010010",
2209 => "0000000000010010",
2210 => "0000000000010010",
2211 => "0000000000010010",
2212 => "0000000000010010",
2213 => "0000000000010010",
2214 => "0000000000010010",
2215 => "0000000000010010",
2216 => "0000000000010010",
2217 => "0000000000010010",
2218 => "0000000000010010",
2219 => "0000000000010010",
2220 => "0000000000010010",
2221 => "0000000000010010",
2222 => "0000000000010010",
2223 => "0000000000010010",
2224 => "0000000000010010",
2225 => "0000000000010010",
2226 => "0000000000010010",
2227 => "0000000000010010",
2228 => "0000000000010010",
2229 => "0000000000010010",
2230 => "0000000000010010",
2231 => "0000000000010010",
2232 => "0000000000010010",
2233 => "0000000000010010",
2234 => "0000000000010010",
2235 => "0000000000010010",
2236 => "0000000000010010",
2237 => "0000000000010010",
2238 => "0000000000010010",
2239 => "0000000000010010",
2240 => "0000000000010010",
2241 => "0000000000010010",
2242 => "0000000000010010",
2243 => "0000000000010011",
2244 => "0000000000010011",
2245 => "0000000000010011",
2246 => "0000000000010011",
2247 => "0000000000010011",
2248 => "0000000000010011",
2249 => "0000000000010011",
2250 => "0000000000010011",
2251 => "0000000000010011",
2252 => "0000000000010011",
2253 => "0000000000010011",
2254 => "0000000000010011",
2255 => "0000000000010011",
2256 => "0000000000010011",
2257 => "0000000000010011",
2258 => "0000000000010011",
2259 => "0000000000010011",
2260 => "0000000000010011",
2261 => "0000000000010011",
2262 => "0000000000010011",
2263 => "0000000000010011",
2264 => "0000000000010011",
2265 => "0000000000010011",
2266 => "0000000000010011",
2267 => "0000000000010011",
2268 => "0000000000010011",
2269 => "0000000000010011",
2270 => "0000000000010011",
2271 => "0000000000010011",
2272 => "0000000000010011",
2273 => "0000000000010011",
2274 => "0000000000010011",
2275 => "0000000000010011",
2276 => "0000000000010011",
2277 => "0000000000010011",
2278 => "0000000000010011",
2279 => "0000000000010011",
2280 => "0000000000010011",
2281 => "0000000000010011",
2282 => "0000000000010011",
2283 => "0000000000010011",
2284 => "0000000000010011",
2285 => "0000000000010011",
2286 => "0000000000010011",
2287 => "0000000000010011",
2288 => "0000000000010011",
2289 => "0000000000010011",
2290 => "0000000000010011",
2291 => "0000000000010011",
2292 => "0000000000010011",
2293 => "0000000000010011",
2294 => "0000000000010011",
2295 => "0000000000010011",
2296 => "0000000000010011",
2297 => "0000000000010011",
2298 => "0000000000010011",
2299 => "0000000000010011",
2300 => "0000000000010011",
2301 => "0000000000010011",
2302 => "0000000000010011",
2303 => "0000000000010011",
2304 => "0000000000010011",
2305 => "0000000000010011",
2306 => "0000000000010011",
2307 => "0000000000010011",
2308 => "0000000000010011",
2309 => "0000000000010011",
2310 => "0000000000010011",
2311 => "0000000000010011",
2312 => "0000000000010011",
2313 => "0000000000010011",
2314 => "0000000000010011",
2315 => "0000000000010011",
2316 => "0000000000010011",
2317 => "0000000000010011",
2318 => "0000000000010011",
2319 => "0000000000010011",
2320 => "0000000000010011",
2321 => "0000000000010011",
2322 => "0000000000010011",
2323 => "0000000000010011",
2324 => "0000000000010011",
2325 => "0000000000010011",
2326 => "0000000000010011",
2327 => "0000000000010011",
2328 => "0000000000010011",
2329 => "0000000000010011",
2330 => "0000000000010011",
2331 => "0000000000010011",
2332 => "0000000000010011",
2333 => "0000000000010011",
2334 => "0000000000010011",
2335 => "0000000000010011",
2336 => "0000000000010011",
2337 => "0000000000010011",
2338 => "0000000000010011",
2339 => "0000000000010011",
2340 => "0000000000010011",
2341 => "0000000000010011",
2342 => "0000000000010011",
2343 => "0000000000010011",
2344 => "0000000000010011",
2345 => "0000000000010011",
2346 => "0000000000010011",
2347 => "0000000000010011",
2348 => "0000000000010011",
2349 => "0000000000010011",
2350 => "0000000000010011",
2351 => "0000000000010011",
2352 => "0000000000010011",
2353 => "0000000000010011",
2354 => "0000000000010011",
2355 => "0000000000010011",
2356 => "0000000000010011",
2357 => "0000000000010011",
2358 => "0000000000010011",
2359 => "0000000000010011",
2360 => "0000000000010011",
2361 => "0000000000010011",
2362 => "0000000000010011",
2363 => "0000000000010011",
2364 => "0000000000010011",
2365 => "0000000000010011",
2366 => "0000000000010011",
2367 => "0000000000010011",
2368 => "0000000000010011",
2369 => "0000000000010011",
2370 => "0000000000010011",
2371 => "0000000000010011",
2372 => "0000000000010011",
2373 => "0000000000010011",
2374 => "0000000000010011",
2375 => "0000000000010011",
2376 => "0000000000010011",
2377 => "0000000000010011",
2378 => "0000000000010011",
2379 => "0000000000010011",
2380 => "0000000000010011",
2381 => "0000000000010011",
2382 => "0000000000010011",
2383 => "0000000000010011",
2384 => "0000000000010011",
2385 => "0000000000010011",
2386 => "0000000000010011",
2387 => "0000000000010011",
2388 => "0000000000010011",
2389 => "0000000000010011",
2390 => "0000000000010011",
2391 => "0000000000010011",
2392 => "0000000000010011",
2393 => "0000000000010011",
2394 => "0000000000010011",
2395 => "0000000000010011",
2396 => "0000000000010011",
2397 => "0000000000010011",
2398 => "0000000000010011",
2399 => "0000000000010011",
2400 => "0000000000010011",
2401 => "0000000000010011",
2402 => "0000000000010011",
2403 => "0000000000010011",
2404 => "0000000000010011",
2405 => "0000000000010011",
2406 => "0000000000010011",
2407 => "0000000000010011",
2408 => "0000000000010011",
2409 => "0000000000010011",
2410 => "0000000000010011",
2411 => "0000000000010011",
2412 => "0000000000010011",
2413 => "0000000000010011",
2414 => "0000000000010011",
2415 => "0000000000010011",
2416 => "0000000000010011",
2417 => "0000000000010011",
2418 => "0000000000010011",
2419 => "0000000000010011",
2420 => "0000000000010011",
2421 => "0000000000010011",
2422 => "0000000000010011",
2423 => "0000000000010011",
2424 => "0000000000010011",
2425 => "0000000000010011",
2426 => "0000000000010011",
2427 => "0000000000010011",
2428 => "0000000000010011",
2429 => "0000000000010011",
2430 => "0000000000010011",
2431 => "0000000000010011",
2432 => "0000000000010011",
2433 => "0000000000010011",
2434 => "0000000000010011",
2435 => "0000000000010011",
2436 => "0000000000010011",
2437 => "0000000000010011",
2438 => "0000000000010011",
2439 => "0000000000010011",
2440 => "0000000000010011",
2441 => "0000000000010011",
2442 => "0000000000010011",
2443 => "0000000000010011",
2444 => "0000000000010011",
2445 => "0000000000010011",
2446 => "0000000000010011",
2447 => "0000000000010011",
2448 => "0000000000010011",
2449 => "0000000000010011",
2450 => "0000000000010011",
2451 => "0000000000010011",
2452 => "0000000000010011",
2453 => "0000000000010100",
2454 => "0000000000010100",
2455 => "0000000000010100",
2456 => "0000000000010100",
2457 => "0000000000010100",
2458 => "0000000000010100",
2459 => "0000000000010100",
2460 => "0000000000010100",
2461 => "0000000000010100",
2462 => "0000000000010100",
2463 => "0000000000010100",
2464 => "0000000000010100",
2465 => "0000000000010100",
2466 => "0000000000010100",
2467 => "0000000000010100",
2468 => "0000000000010100",
2469 => "0000000000010100",
2470 => "0000000000010100",
2471 => "0000000000010100",
2472 => "0000000000010100",
2473 => "0000000000010100",
2474 => "0000000000010100",
2475 => "0000000000010100",
2476 => "0000000000010100",
2477 => "0000000000010100",
2478 => "0000000000010100",
2479 => "0000000000010100",
2480 => "0000000000010100",
2481 => "0000000000010100",
2482 => "0000000000010100",
2483 => "0000000000010100",
2484 => "0000000000010100",
2485 => "0000000000010100",
2486 => "0000000000010100",
2487 => "0000000000010100",
2488 => "0000000000010100",
2489 => "0000000000010100",
2490 => "0000000000010100",
2491 => "0000000000010100",
2492 => "0000000000010100",
2493 => "0000000000010100",
2494 => "0000000000010100",
2495 => "0000000000010100",
2496 => "0000000000010100",
2497 => "0000000000010100",
2498 => "0000000000010100",
2499 => "0000000000010100",
2500 => "0000000000010100",
2501 => "0000000000010100",
2502 => "0000000000010100",
2503 => "0000000000010100",
2504 => "0000000000010100",
2505 => "0000000000010100",
2506 => "0000000000010100",
2507 => "0000000000010100",
2508 => "0000000000010100",
2509 => "0000000000010100",
2510 => "0000000000010100",
2511 => "0000000000010100",
2512 => "0000000000010100",
2513 => "0000000000010100",
2514 => "0000000000010100",
2515 => "0000000000010100",
2516 => "0000000000010100",
2517 => "0000000000010100",
2518 => "0000000000010100",
2519 => "0000000000010100",
2520 => "0000000000010100",
2521 => "0000000000010100",
2522 => "0000000000010100",
2523 => "0000000000010100",
2524 => "0000000000010100",
2525 => "0000000000010100",
2526 => "0000000000010100",
2527 => "0000000000010100",
2528 => "0000000000010100",
2529 => "0000000000010100",
2530 => "0000000000010100",
2531 => "0000000000010100",
2532 => "0000000000010100",
2533 => "0000000000010100",
2534 => "0000000000010100",
2535 => "0000000000010100",
2536 => "0000000000010100",
2537 => "0000000000010100",
2538 => "0000000000010100",
2539 => "0000000000010100",
2540 => "0000000000010100",
2541 => "0000000000010100",
2542 => "0000000000010100",
2543 => "0000000000010100",
2544 => "0000000000010100",
2545 => "0000000000010100",
2546 => "0000000000010100",
2547 => "0000000000010100",
2548 => "0000000000010100",
2549 => "0000000000010100",
2550 => "0000000000010100",
2551 => "0000000000010100",
2552 => "0000000000010100",
2553 => "0000000000010100",
2554 => "0000000000010100",
2555 => "0000000000010100",
2556 => "0000000000010100",
2557 => "0000000000010100",
2558 => "0000000000010100",
2559 => "0000000000010100",
2560 => "0000000000010100",
2561 => "0000000000010100",
2562 => "0000000000010100",
2563 => "0000000000010100",
2564 => "0000000000010100",
2565 => "0000000000010100",
2566 => "0000000000010100",
2567 => "0000000000010100",
2568 => "0000000000010100",
2569 => "0000000000010100",
2570 => "0000000000010100",
2571 => "0000000000010100",
2572 => "0000000000010100",
2573 => "0000000000010100",
2574 => "0000000000010100",
2575 => "0000000000010100",
2576 => "0000000000010100",
2577 => "0000000000010100",
2578 => "0000000000010100",
2579 => "0000000000010100",
2580 => "0000000000010100",
2581 => "0000000000010100",
2582 => "0000000000010100",
2583 => "0000000000010100",
2584 => "0000000000010100",
2585 => "0000000000010100",
2586 => "0000000000010100",
2587 => "0000000000010100",
2588 => "0000000000010100",
2589 => "0000000000010100",
2590 => "0000000000010100",
2591 => "0000000000010100",
2592 => "0000000000010100",
2593 => "0000000000010100",
2594 => "0000000000010100",
2595 => "0000000000010100",
2596 => "0000000000010100",
2597 => "0000000000010100",
2598 => "0000000000010100",
2599 => "0000000000010100",
2600 => "0000000000010100",
2601 => "0000000000010100",
2602 => "0000000000010100",
2603 => "0000000000010100",
2604 => "0000000000010100",
2605 => "0000000000010100",
2606 => "0000000000010100",
2607 => "0000000000010100",
2608 => "0000000000010100",
2609 => "0000000000010100",
2610 => "0000000000010100",
2611 => "0000000000010100",
2612 => "0000000000010100",
2613 => "0000000000010100",
2614 => "0000000000010100",
2615 => "0000000000010100",
2616 => "0000000000010100",
2617 => "0000000000010100",
2618 => "0000000000010100",
2619 => "0000000000010100",
2620 => "0000000000010100",
2621 => "0000000000010100",
2622 => "0000000000010100",
2623 => "0000000000010100",
2624 => "0000000000010100",
2625 => "0000000000010100",
2626 => "0000000000010100",
2627 => "0000000000010100",
2628 => "0000000000010100",
2629 => "0000000000010100",
2630 => "0000000000010100",
2631 => "0000000000010100",
2632 => "0000000000010100",
2633 => "0000000000010100",
2634 => "0000000000010100",
2635 => "0000000000010100",
2636 => "0000000000010100",
2637 => "0000000000010100",
2638 => "0000000000010100",
2639 => "0000000000010100",
2640 => "0000000000010100",
2641 => "0000000000010100",
2642 => "0000000000010100",
2643 => "0000000000010100",
2644 => "0000000000010100",
2645 => "0000000000010100",
2646 => "0000000000010100",
2647 => "0000000000010100",
2648 => "0000000000010100",
2649 => "0000000000010100",
2650 => "0000000000010100",
2651 => "0000000000010100",
2652 => "0000000000010100",
2653 => "0000000000010101",
2654 => "0000000000010101",
2655 => "0000000000010101",
2656 => "0000000000010101",
2657 => "0000000000010101",
2658 => "0000000000010101",
2659 => "0000000000010101",
2660 => "0000000000010101",
2661 => "0000000000010101",
2662 => "0000000000010101",
2663 => "0000000000010101",
2664 => "0000000000010101",
2665 => "0000000000010101",
2666 => "0000000000010101",
2667 => "0000000000010101",
2668 => "0000000000010101",
2669 => "0000000000010101",
2670 => "0000000000010101",
2671 => "0000000000010101",
2672 => "0000000000010101",
2673 => "0000000000010101",
2674 => "0000000000010101",
2675 => "0000000000010101",
2676 => "0000000000010101",
2677 => "0000000000010101",
2678 => "0000000000010101",
2679 => "0000000000010101",
2680 => "0000000000010101",
2681 => "0000000000010101",
2682 => "0000000000010101",
2683 => "0000000000010101",
2684 => "0000000000010101",
2685 => "0000000000010101",
2686 => "0000000000010101",
2687 => "0000000000010101",
2688 => "0000000000010101",
2689 => "0000000000010101",
2690 => "0000000000010101",
2691 => "0000000000010101",
2692 => "0000000000010101",
2693 => "0000000000010101",
2694 => "0000000000010101",
2695 => "0000000000010101",
2696 => "0000000000010101",
2697 => "0000000000010101",
2698 => "0000000000010101",
2699 => "0000000000010101",
2700 => "0000000000010101",
2701 => "0000000000010101",
2702 => "0000000000010101",
2703 => "0000000000010101",
2704 => "0000000000010101",
2705 => "0000000000010101",
2706 => "0000000000010101",
2707 => "0000000000010101",
2708 => "0000000000010101",
2709 => "0000000000010101",
2710 => "0000000000010101",
2711 => "0000000000010101",
2712 => "0000000000010101",
2713 => "0000000000010101",
2714 => "0000000000010101",
2715 => "0000000000010101",
2716 => "0000000000010101",
2717 => "0000000000010101",
2718 => "0000000000010101",
2719 => "0000000000010101",
2720 => "0000000000010101",
2721 => "0000000000010101",
2722 => "0000000000010101",
2723 => "0000000000010101",
2724 => "0000000000010101",
2725 => "0000000000010101",
2726 => "0000000000010101",
2727 => "0000000000010101",
2728 => "0000000000010101",
2729 => "0000000000010101",
2730 => "0000000000010101",
2731 => "0000000000010101",
2732 => "0000000000010101",
2733 => "0000000000010101",
2734 => "0000000000010101",
2735 => "0000000000010101",
2736 => "0000000000010101",
2737 => "0000000000010101",
2738 => "0000000000010101",
2739 => "0000000000010101",
2740 => "0000000000010101",
2741 => "0000000000010101",
2742 => "0000000000010101",
2743 => "0000000000010101",
2744 => "0000000000010101",
2745 => "0000000000010101",
2746 => "0000000000010101",
2747 => "0000000000010101",
2748 => "0000000000010101",
2749 => "0000000000010101",
2750 => "0000000000010101",
2751 => "0000000000010101",
2752 => "0000000000010101",
2753 => "0000000000010101",
2754 => "0000000000010101",
2755 => "0000000000010101",
2756 => "0000000000010101",
2757 => "0000000000010101",
2758 => "0000000000010101",
2759 => "0000000000010101",
2760 => "0000000000010101",
2761 => "0000000000010101",
2762 => "0000000000010101",
2763 => "0000000000010101",
2764 => "0000000000010101",
2765 => "0000000000010101",
2766 => "0000000000010101",
2767 => "0000000000010101",
2768 => "0000000000010101",
2769 => "0000000000010101",
2770 => "0000000000010101",
2771 => "0000000000010101",
2772 => "0000000000010101",
2773 => "0000000000010101",
2774 => "0000000000010101",
2775 => "0000000000010101",
2776 => "0000000000010101",
2777 => "0000000000010101",
2778 => "0000000000010101",
2779 => "0000000000010101",
2780 => "0000000000010101",
2781 => "0000000000010101",
2782 => "0000000000010101",
2783 => "0000000000010101",
2784 => "0000000000010101",
2785 => "0000000000010101",
2786 => "0000000000010101",
2787 => "0000000000010101",
2788 => "0000000000010101",
2789 => "0000000000010101",
2790 => "0000000000010101",
2791 => "0000000000010101",
2792 => "0000000000010101",
2793 => "0000000000010101",
2794 => "0000000000010101",
2795 => "0000000000010101",
2796 => "0000000000010101",
2797 => "0000000000010101",
2798 => "0000000000010101",
2799 => "0000000000010101",
2800 => "0000000000010101",
2801 => "0000000000010101",
2802 => "0000000000010101",
2803 => "0000000000010101",
2804 => "0000000000010101",
2805 => "0000000000010101",
2806 => "0000000000010101",
2807 => "0000000000010101",
2808 => "0000000000010101",
2809 => "0000000000010101",
2810 => "0000000000010101",
2811 => "0000000000010101",
2812 => "0000000000010101",
2813 => "0000000000010101",
2814 => "0000000000010101",
2815 => "0000000000010101",
2816 => "0000000000010101",
2817 => "0000000000010101",
2818 => "0000000000010101",
2819 => "0000000000010101",
2820 => "0000000000010101",
2821 => "0000000000010101",
2822 => "0000000000010101",
2823 => "0000000000010101",
2824 => "0000000000010101",
2825 => "0000000000010101",
2826 => "0000000000010101",
2827 => "0000000000010101",
2828 => "0000000000010101",
2829 => "0000000000010101",
2830 => "0000000000010101",
2831 => "0000000000010101",
2832 => "0000000000010101",
2833 => "0000000000010101",
2834 => "0000000000010101",
2835 => "0000000000010101",
2836 => "0000000000010101",
2837 => "0000000000010101",
2838 => "0000000000010101",
2839 => "0000000000010101",
2840 => "0000000000010101",
2841 => "0000000000010101",
2842 => "0000000000010101",
2843 => "0000000000010101",
2844 => "0000000000010110",
2845 => "0000000000010110",
2846 => "0000000000010110",
2847 => "0000000000010110",
2848 => "0000000000010110",
2849 => "0000000000010110",
2850 => "0000000000010110",
2851 => "0000000000010110",
2852 => "0000000000010110",
2853 => "0000000000010110",
2854 => "0000000000010110",
2855 => "0000000000010110",
2856 => "0000000000010110",
2857 => "0000000000010110",
2858 => "0000000000010110",
2859 => "0000000000010110",
2860 => "0000000000010110",
2861 => "0000000000010110",
2862 => "0000000000010110",
2863 => "0000000000010110",
2864 => "0000000000010110",
2865 => "0000000000010110",
2866 => "0000000000010110",
2867 => "0000000000010110",
2868 => "0000000000010110",
2869 => "0000000000010110",
2870 => "0000000000010110",
2871 => "0000000000010110",
2872 => "0000000000010110",
2873 => "0000000000010110",
2874 => "0000000000010110",
2875 => "0000000000010110",
2876 => "0000000000010110",
2877 => "0000000000010110",
2878 => "0000000000010110",
2879 => "0000000000010110",
2880 => "0000000000010110",
2881 => "0000000000010110",
2882 => "0000000000010110",
2883 => "0000000000010110",
2884 => "0000000000010110",
2885 => "0000000000010110",
2886 => "0000000000010110",
2887 => "0000000000010110",
2888 => "0000000000010110",
2889 => "0000000000010110",
2890 => "0000000000010110",
2891 => "0000000000010110",
2892 => "0000000000010110",
2893 => "0000000000010110",
2894 => "0000000000010110",
2895 => "0000000000010110",
2896 => "0000000000010110",
2897 => "0000000000010110",
2898 => "0000000000010110",
2899 => "0000000000010110",
2900 => "0000000000010110",
2901 => "0000000000010110",
2902 => "0000000000010110",
2903 => "0000000000010110",
2904 => "0000000000010110",
2905 => "0000000000010110",
2906 => "0000000000010110",
2907 => "0000000000010110",
2908 => "0000000000010110",
2909 => "0000000000010110",
2910 => "0000000000010110",
2911 => "0000000000010110",
2912 => "0000000000010110",
2913 => "0000000000010110",
2914 => "0000000000010110",
2915 => "0000000000010110",
2916 => "0000000000010110",
2917 => "0000000000010110",
2918 => "0000000000010110",
2919 => "0000000000010110",
2920 => "0000000000010110",
2921 => "0000000000010110",
2922 => "0000000000010110",
2923 => "0000000000010110",
2924 => "0000000000010110",
2925 => "0000000000010110",
2926 => "0000000000010110",
2927 => "0000000000010110",
2928 => "0000000000010110",
2929 => "0000000000010110",
2930 => "0000000000010110",
2931 => "0000000000010110",
2932 => "0000000000010110",
2933 => "0000000000010110",
2934 => "0000000000010110",
2935 => "0000000000010110",
2936 => "0000000000010110",
2937 => "0000000000010110",
2938 => "0000000000010110",
2939 => "0000000000010110",
2940 => "0000000000010110",
2941 => "0000000000010110",
2942 => "0000000000010110",
2943 => "0000000000010110",
2944 => "0000000000010110",
2945 => "0000000000010110",
2946 => "0000000000010110",
2947 => "0000000000010110",
2948 => "0000000000010110",
2949 => "0000000000010110",
2950 => "0000000000010110",
2951 => "0000000000010110",
2952 => "0000000000010110",
2953 => "0000000000010110",
2954 => "0000000000010110",
2955 => "0000000000010110",
2956 => "0000000000010110",
2957 => "0000000000010110",
2958 => "0000000000010110",
2959 => "0000000000010110",
2960 => "0000000000010110",
2961 => "0000000000010110",
2962 => "0000000000010110",
2963 => "0000000000010110",
2964 => "0000000000010110",
2965 => "0000000000010110",
2966 => "0000000000010110",
2967 => "0000000000010110",
2968 => "0000000000010110",
2969 => "0000000000010110",
2970 => "0000000000010110",
2971 => "0000000000010110",
2972 => "0000000000010110",
2973 => "0000000000010110",
2974 => "0000000000010110",
2975 => "0000000000010110",
2976 => "0000000000010110",
2977 => "0000000000010110",
2978 => "0000000000010110",
2979 => "0000000000010110",
2980 => "0000000000010110",
2981 => "0000000000010110",
2982 => "0000000000010110",
2983 => "0000000000010110",
2984 => "0000000000010110",
2985 => "0000000000010110",
2986 => "0000000000010110",
2987 => "0000000000010110",
2988 => "0000000000010110",
2989 => "0000000000010110",
2990 => "0000000000010110",
2991 => "0000000000010110",
2992 => "0000000000010110",
2993 => "0000000000010110",
2994 => "0000000000010110",
2995 => "0000000000010110",
2996 => "0000000000010110",
2997 => "0000000000010110",
2998 => "0000000000010110",
2999 => "0000000000010110",
3000 => "0000000000010110",
3001 => "0000000000010110",
3002 => "0000000000010110",
3003 => "0000000000010110",
3004 => "0000000000010110",
3005 => "0000000000010110",
3006 => "0000000000010110",
3007 => "0000000000010110",
3008 => "0000000000010110",
3009 => "0000000000010110",
3010 => "0000000000010110",
3011 => "0000000000010110",
3012 => "0000000000010110",
3013 => "0000000000010110",
3014 => "0000000000010110",
3015 => "0000000000010110",
3016 => "0000000000010110",
3017 => "0000000000010110",
3018 => "0000000000010110",
3019 => "0000000000010110",
3020 => "0000000000010110",
3021 => "0000000000010110",
3022 => "0000000000010110",
3023 => "0000000000010110",
3024 => "0000000000010110",
3025 => "0000000000010110",
3026 => "0000000000010111",
3027 => "0000000000010111",
3028 => "0000000000010111",
3029 => "0000000000010111",
3030 => "0000000000010111",
3031 => "0000000000010111",
3032 => "0000000000010111",
3033 => "0000000000010111",
3034 => "0000000000010111",
3035 => "0000000000010111",
3036 => "0000000000010111",
3037 => "0000000000010111",
3038 => "0000000000010111",
3039 => "0000000000010111",
3040 => "0000000000010111",
3041 => "0000000000010111",
3042 => "0000000000010111",
3043 => "0000000000010111",
3044 => "0000000000010111",
3045 => "0000000000010111",
3046 => "0000000000010111",
3047 => "0000000000010111",
3048 => "0000000000010111",
3049 => "0000000000010111",
3050 => "0000000000010111",
3051 => "0000000000010111",
3052 => "0000000000010111",
3053 => "0000000000010111",
3054 => "0000000000010111",
3055 => "0000000000010111",
3056 => "0000000000010111",
3057 => "0000000000010111",
3058 => "0000000000010111",
3059 => "0000000000010111",
3060 => "0000000000010111",
3061 => "0000000000010111",
3062 => "0000000000010111",
3063 => "0000000000010111",
3064 => "0000000000010111",
3065 => "0000000000010111",
3066 => "0000000000010111",
3067 => "0000000000010111",
3068 => "0000000000010111",
3069 => "0000000000010111",
3070 => "0000000000010111",
3071 => "0000000000010111",
3072 => "0000000000010111",
3073 => "0000000000010111",
3074 => "0000000000010111",
3075 => "0000000000010111",
3076 => "0000000000010111",
3077 => "0000000000010111",
3078 => "0000000000010111",
3079 => "0000000000010111",
3080 => "0000000000010111",
3081 => "0000000000010111",
3082 => "0000000000010111",
3083 => "0000000000010111",
3084 => "0000000000010111",
3085 => "0000000000010111",
3086 => "0000000000010111",
3087 => "0000000000010111",
3088 => "0000000000010111",
3089 => "0000000000010111",
3090 => "0000000000010111",
3091 => "0000000000010111",
3092 => "0000000000010111",
3093 => "0000000000010111",
3094 => "0000000000010111",
3095 => "0000000000010111",
3096 => "0000000000010111",
3097 => "0000000000010111",
3098 => "0000000000010111",
3099 => "0000000000010111",
3100 => "0000000000010111",
3101 => "0000000000010111",
3102 => "0000000000010111",
3103 => "0000000000010111",
3104 => "0000000000010111",
3105 => "0000000000010111",
3106 => "0000000000010111",
3107 => "0000000000010111",
3108 => "0000000000010111",
3109 => "0000000000010111",
3110 => "0000000000010111",
3111 => "0000000000010111",
3112 => "0000000000010111",
3113 => "0000000000010111",
3114 => "0000000000010111",
3115 => "0000000000010111",
3116 => "0000000000010111",
3117 => "0000000000010111",
3118 => "0000000000010111",
3119 => "0000000000010111",
3120 => "0000000000010111",
3121 => "0000000000010111",
3122 => "0000000000010111",
3123 => "0000000000010111",
3124 => "0000000000010111",
3125 => "0000000000010111",
3126 => "0000000000010111",
3127 => "0000000000010111",
3128 => "0000000000010111",
3129 => "0000000000010111",
3130 => "0000000000010111",
3131 => "0000000000010111",
3132 => "0000000000010111",
3133 => "0000000000010111",
3134 => "0000000000010111",
3135 => "0000000000010111",
3136 => "0000000000010111",
3137 => "0000000000010111",
3138 => "0000000000010111",
3139 => "0000000000010111",
3140 => "0000000000010111",
3141 => "0000000000010111",
3142 => "0000000000010111",
3143 => "0000000000010111",
3144 => "0000000000010111",
3145 => "0000000000010111",
3146 => "0000000000010111",
3147 => "0000000000010111",
3148 => "0000000000010111",
3149 => "0000000000010111",
3150 => "0000000000010111",
3151 => "0000000000010111",
3152 => "0000000000010111",
3153 => "0000000000010111",
3154 => "0000000000010111",
3155 => "0000000000010111",
3156 => "0000000000010111",
3157 => "0000000000010111",
3158 => "0000000000010111",
3159 => "0000000000010111",
3160 => "0000000000010111",
3161 => "0000000000010111",
3162 => "0000000000010111",
3163 => "0000000000010111",
3164 => "0000000000010111",
3165 => "0000000000010111",
3166 => "0000000000010111",
3167 => "0000000000010111",
3168 => "0000000000010111",
3169 => "0000000000010111",
3170 => "0000000000010111",
3171 => "0000000000010111",
3172 => "0000000000010111",
3173 => "0000000000010111",
3174 => "0000000000010111",
3175 => "0000000000010111",
3176 => "0000000000010111",
3177 => "0000000000010111",
3178 => "0000000000010111",
3179 => "0000000000010111",
3180 => "0000000000010111",
3181 => "0000000000010111",
3182 => "0000000000010111",
3183 => "0000000000010111",
3184 => "0000000000010111",
3185 => "0000000000010111",
3186 => "0000000000010111",
3187 => "0000000000010111",
3188 => "0000000000010111",
3189 => "0000000000010111",
3190 => "0000000000010111",
3191 => "0000000000010111",
3192 => "0000000000010111",
3193 => "0000000000010111",
3194 => "0000000000010111",
3195 => "0000000000010111",
3196 => "0000000000010111",
3197 => "0000000000010111",
3198 => "0000000000010111",
3199 => "0000000000010111",
3200 => "0000000000011000",
3201 => "0000000000011000",
3202 => "0000000000011000",
3203 => "0000000000011000",
3204 => "0000000000011000",
3205 => "0000000000011000",
3206 => "0000000000011000",
3207 => "0000000000011000",
3208 => "0000000000011000",
3209 => "0000000000011000",
3210 => "0000000000011000",
3211 => "0000000000011000",
3212 => "0000000000011000",
3213 => "0000000000011000",
3214 => "0000000000011000",
3215 => "0000000000011000",
3216 => "0000000000011000",
3217 => "0000000000011000",
3218 => "0000000000011000",
3219 => "0000000000011000",
3220 => "0000000000011000",
3221 => "0000000000011000",
3222 => "0000000000011000",
3223 => "0000000000011000",
3224 => "0000000000011000",
3225 => "0000000000011000",
3226 => "0000000000011000",
3227 => "0000000000011000",
3228 => "0000000000011000",
3229 => "0000000000011000",
3230 => "0000000000011000",
3231 => "0000000000011000",
3232 => "0000000000011000",
3233 => "0000000000011000",
3234 => "0000000000011000",
3235 => "0000000000011000",
3236 => "0000000000011000",
3237 => "0000000000011000",
3238 => "0000000000011000",
3239 => "0000000000011000",
3240 => "0000000000011000",
3241 => "0000000000011000",
3242 => "0000000000011000",
3243 => "0000000000011000",
3244 => "0000000000011000",
3245 => "0000000000011000",
3246 => "0000000000011000",
3247 => "0000000000011000",
3248 => "0000000000011000",
3249 => "0000000000011000",
3250 => "0000000000011000",
3251 => "0000000000011000",
3252 => "0000000000011000",
3253 => "0000000000011000",
3254 => "0000000000011000",
3255 => "0000000000011000",
3256 => "0000000000011000",
3257 => "0000000000011000",
3258 => "0000000000011000",
3259 => "0000000000011000",
3260 => "0000000000011000",
3261 => "0000000000011000",
3262 => "0000000000011000",
3263 => "0000000000011000",
3264 => "0000000000011000",
3265 => "0000000000011000",
3266 => "0000000000011000",
3267 => "0000000000011000",
3268 => "0000000000011000",
3269 => "0000000000011000",
3270 => "0000000000011000",
3271 => "0000000000011000",
3272 => "0000000000011000",
3273 => "0000000000011000",
3274 => "0000000000011000",
3275 => "0000000000011000",
3276 => "0000000000011000",
3277 => "0000000000011000",
3278 => "0000000000011000",
3279 => "0000000000011000",
3280 => "0000000000011000",
3281 => "0000000000011000",
3282 => "0000000000011000",
3283 => "0000000000011000",
3284 => "0000000000011000",
3285 => "0000000000011000",
3286 => "0000000000011000",
3287 => "0000000000011000",
3288 => "0000000000011000",
3289 => "0000000000011000",
3290 => "0000000000011000",
3291 => "0000000000011000",
3292 => "0000000000011000",
3293 => "0000000000011000",
3294 => "0000000000011000",
3295 => "0000000000011000",
3296 => "0000000000011000",
3297 => "0000000000011000",
3298 => "0000000000011000",
3299 => "0000000000011000",
3300 => "0000000000011000",
3301 => "0000000000011000",
3302 => "0000000000011000",
3303 => "0000000000011000",
3304 => "0000000000011000",
3305 => "0000000000011000",
3306 => "0000000000011000",
3307 => "0000000000011000",
3308 => "0000000000011000",
3309 => "0000000000011000",
3310 => "0000000000011000",
3311 => "0000000000011000",
3312 => "0000000000011000",
3313 => "0000000000011000",
3314 => "0000000000011000",
3315 => "0000000000011000",
3316 => "0000000000011000",
3317 => "0000000000011000",
3318 => "0000000000011000",
3319 => "0000000000011000",
3320 => "0000000000011000",
3321 => "0000000000011000",
3322 => "0000000000011000",
3323 => "0000000000011000",
3324 => "0000000000011000",
3325 => "0000000000011000",
3326 => "0000000000011000",
3327 => "0000000000011000",
3328 => "0000000000011000",
3329 => "0000000000011000",
3330 => "0000000000011000",
3331 => "0000000000011000",
3332 => "0000000000011000",
3333 => "0000000000011000",
3334 => "0000000000011000",
3335 => "0000000000011000",
3336 => "0000000000011000",
3337 => "0000000000011000",
3338 => "0000000000011000",
3339 => "0000000000011000",
3340 => "0000000000011000",
3341 => "0000000000011000",
3342 => "0000000000011000",
3343 => "0000000000011000",
3344 => "0000000000011000",
3345 => "0000000000011000",
3346 => "0000000000011000",
3347 => "0000000000011000",
3348 => "0000000000011000",
3349 => "0000000000011000",
3350 => "0000000000011000",
3351 => "0000000000011000",
3352 => "0000000000011000",
3353 => "0000000000011000",
3354 => "0000000000011000",
3355 => "0000000000011000",
3356 => "0000000000011000",
3357 => "0000000000011000",
3358 => "0000000000011000",
3359 => "0000000000011000",
3360 => "0000000000011000",
3361 => "0000000000011000",
3362 => "0000000000011000",
3363 => "0000000000011000",
3364 => "0000000000011000",
3365 => "0000000000011000",
3366 => "0000000000011000",
3367 => "0000000000011000",
3368 => "0000000000011001",
3369 => "0000000000011001",
3370 => "0000000000011001",
3371 => "0000000000011001",
3372 => "0000000000011001",
3373 => "0000000000011001",
3374 => "0000000000011001",
3375 => "0000000000011001",
3376 => "0000000000011001",
3377 => "0000000000011001",
3378 => "0000000000011001",
3379 => "0000000000011001",
3380 => "0000000000011001",
3381 => "0000000000011001",
3382 => "0000000000011001",
3383 => "0000000000011001",
3384 => "0000000000011001",
3385 => "0000000000011001",
3386 => "0000000000011001",
3387 => "0000000000011001",
3388 => "0000000000011001",
3389 => "0000000000011001",
3390 => "0000000000011001",
3391 => "0000000000011001",
3392 => "0000000000011001",
3393 => "0000000000011001",
3394 => "0000000000011001",
3395 => "0000000000011001",
3396 => "0000000000011001",
3397 => "0000000000011001",
3398 => "0000000000011001",
3399 => "0000000000011001",
3400 => "0000000000011001",
3401 => "0000000000011001",
3402 => "0000000000011001",
3403 => "0000000000011001",
3404 => "0000000000011001",
3405 => "0000000000011001",
3406 => "0000000000011001",
3407 => "0000000000011001",
3408 => "0000000000011001",
3409 => "0000000000011001",
3410 => "0000000000011001",
3411 => "0000000000011001",
3412 => "0000000000011001",
3413 => "0000000000011001",
3414 => "0000000000011001",
3415 => "0000000000011001",
3416 => "0000000000011001",
3417 => "0000000000011001",
3418 => "0000000000011001",
3419 => "0000000000011001",
3420 => "0000000000011001",
3421 => "0000000000011001",
3422 => "0000000000011001",
3423 => "0000000000011001",
3424 => "0000000000011001",
3425 => "0000000000011001",
3426 => "0000000000011001",
3427 => "0000000000011001",
3428 => "0000000000011001",
3429 => "0000000000011001",
3430 => "0000000000011001",
3431 => "0000000000011001",
3432 => "0000000000011001",
3433 => "0000000000011001",
3434 => "0000000000011001",
3435 => "0000000000011001",
3436 => "0000000000011001",
3437 => "0000000000011001",
3438 => "0000000000011001",
3439 => "0000000000011001",
3440 => "0000000000011001",
3441 => "0000000000011001",
3442 => "0000000000011001",
3443 => "0000000000011001",
3444 => "0000000000011001",
3445 => "0000000000011001",
3446 => "0000000000011001",
3447 => "0000000000011001",
3448 => "0000000000011001",
3449 => "0000000000011001",
3450 => "0000000000011001",
3451 => "0000000000011001",
3452 => "0000000000011001",
3453 => "0000000000011001",
3454 => "0000000000011001",
3455 => "0000000000011001",
3456 => "0000000000011001",
3457 => "0000000000011001",
3458 => "0000000000011001",
3459 => "0000000000011001",
3460 => "0000000000011001",
3461 => "0000000000011001",
3462 => "0000000000011001",
3463 => "0000000000011001",
3464 => "0000000000011001",
3465 => "0000000000011001",
3466 => "0000000000011001",
3467 => "0000000000011001",
3468 => "0000000000011001",
3469 => "0000000000011001",
3470 => "0000000000011001",
3471 => "0000000000011001",
3472 => "0000000000011001",
3473 => "0000000000011001",
3474 => "0000000000011001",
3475 => "0000000000011001",
3476 => "0000000000011001",
3477 => "0000000000011001",
3478 => "0000000000011001",
3479 => "0000000000011001",
3480 => "0000000000011001",
3481 => "0000000000011001",
3482 => "0000000000011001",
3483 => "0000000000011001",
3484 => "0000000000011001",
3485 => "0000000000011001",
3486 => "0000000000011001",
3487 => "0000000000011001",
3488 => "0000000000011001",
3489 => "0000000000011001",
3490 => "0000000000011001",
3491 => "0000000000011001",
3492 => "0000000000011001",
3493 => "0000000000011001",
3494 => "0000000000011001",
3495 => "0000000000011001",
3496 => "0000000000011001",
3497 => "0000000000011001",
3498 => "0000000000011001",
3499 => "0000000000011001",
3500 => "0000000000011001",
3501 => "0000000000011001",
3502 => "0000000000011001",
3503 => "0000000000011001",
3504 => "0000000000011001",
3505 => "0000000000011001",
3506 => "0000000000011001",
3507 => "0000000000011001",
3508 => "0000000000011001",
3509 => "0000000000011001",
3510 => "0000000000011001",
3511 => "0000000000011001",
3512 => "0000000000011001",
3513 => "0000000000011001",
3514 => "0000000000011001",
3515 => "0000000000011001",
3516 => "0000000000011001",
3517 => "0000000000011001",
3518 => "0000000000011001",
3519 => "0000000000011001",
3520 => "0000000000011001",
3521 => "0000000000011001",
3522 => "0000000000011001",
3523 => "0000000000011001",
3524 => "0000000000011001",
3525 => "0000000000011001",
3526 => "0000000000011001",
3527 => "0000000000011001",
3528 => "0000000000011001",
3529 => "0000000000011010",
3530 => "0000000000011010",
3531 => "0000000000011010",
3532 => "0000000000011010",
3533 => "0000000000011010",
3534 => "0000000000011010",
3535 => "0000000000011010",
3536 => "0000000000011010",
3537 => "0000000000011010",
3538 => "0000000000011010",
3539 => "0000000000011010",
3540 => "0000000000011010",
3541 => "0000000000011010",
3542 => "0000000000011010",
3543 => "0000000000011010",
3544 => "0000000000011010",
3545 => "0000000000011010",
3546 => "0000000000011010",
3547 => "0000000000011010",
3548 => "0000000000011010",
3549 => "0000000000011010",
3550 => "0000000000011010",
3551 => "0000000000011010",
3552 => "0000000000011010",
3553 => "0000000000011010",
3554 => "0000000000011010",
3555 => "0000000000011010",
3556 => "0000000000011010",
3557 => "0000000000011010",
3558 => "0000000000011010",
3559 => "0000000000011010",
3560 => "0000000000011010",
3561 => "0000000000011010",
3562 => "0000000000011010",
3563 => "0000000000011010",
3564 => "0000000000011010",
3565 => "0000000000011010",
3566 => "0000000000011010",
3567 => "0000000000011010",
3568 => "0000000000011010",
3569 => "0000000000011010",
3570 => "0000000000011010",
3571 => "0000000000011010",
3572 => "0000000000011010",
3573 => "0000000000011010",
3574 => "0000000000011010",
3575 => "0000000000011010",
3576 => "0000000000011010",
3577 => "0000000000011010",
3578 => "0000000000011010",
3579 => "0000000000011010",
3580 => "0000000000011010",
3581 => "0000000000011010",
3582 => "0000000000011010",
3583 => "0000000000011010",
3584 => "0000000000011010",
3585 => "0000000000011010",
3586 => "0000000000011010",
3587 => "0000000000011010",
3588 => "0000000000011010",
3589 => "0000000000011010",
3590 => "0000000000011010",
3591 => "0000000000011010",
3592 => "0000000000011010",
3593 => "0000000000011010",
3594 => "0000000000011010",
3595 => "0000000000011010",
3596 => "0000000000011010",
3597 => "0000000000011010",
3598 => "0000000000011010",
3599 => "0000000000011010",
3600 => "0000000000011010",
3601 => "0000000000011010",
3602 => "0000000000011010",
3603 => "0000000000011010",
3604 => "0000000000011010",
3605 => "0000000000011010",
3606 => "0000000000011010",
3607 => "0000000000011010",
3608 => "0000000000011010",
3609 => "0000000000011010",
3610 => "0000000000011010",
3611 => "0000000000011010",
3612 => "0000000000011010",
3613 => "0000000000011010",
3614 => "0000000000011010",
3615 => "0000000000011010",
3616 => "0000000000011010",
3617 => "0000000000011010",
3618 => "0000000000011010",
3619 => "0000000000011010",
3620 => "0000000000011010",
3621 => "0000000000011010",
3622 => "0000000000011010",
3623 => "0000000000011010",
3624 => "0000000000011010",
3625 => "0000000000011010",
3626 => "0000000000011010",
3627 => "0000000000011010",
3628 => "0000000000011010",
3629 => "0000000000011010",
3630 => "0000000000011010",
3631 => "0000000000011010",
3632 => "0000000000011010",
3633 => "0000000000011010",
3634 => "0000000000011010",
3635 => "0000000000011010",
3636 => "0000000000011010",
3637 => "0000000000011010",
3638 => "0000000000011010",
3639 => "0000000000011010",
3640 => "0000000000011010",
3641 => "0000000000011010",
3642 => "0000000000011010",
3643 => "0000000000011010",
3644 => "0000000000011010",
3645 => "0000000000011010",
3646 => "0000000000011010",
3647 => "0000000000011010",
3648 => "0000000000011010",
3649 => "0000000000011010",
3650 => "0000000000011010",
3651 => "0000000000011010",
3652 => "0000000000011010",
3653 => "0000000000011010",
3654 => "0000000000011010",
3655 => "0000000000011010",
3656 => "0000000000011010",
3657 => "0000000000011010",
3658 => "0000000000011010",
3659 => "0000000000011010",
3660 => "0000000000011010",
3661 => "0000000000011010",
3662 => "0000000000011010",
3663 => "0000000000011010",
3664 => "0000000000011010",
3665 => "0000000000011010",
3666 => "0000000000011010",
3667 => "0000000000011010",
3668 => "0000000000011010",
3669 => "0000000000011010",
3670 => "0000000000011010",
3671 => "0000000000011010",
3672 => "0000000000011010",
3673 => "0000000000011010",
3674 => "0000000000011010",
3675 => "0000000000011010",
3676 => "0000000000011010",
3677 => "0000000000011010",
3678 => "0000000000011010",
3679 => "0000000000011010",
3680 => "0000000000011010",
3681 => "0000000000011010",
3682 => "0000000000011010",
3683 => "0000000000011011",
3684 => "0000000000011011",
3685 => "0000000000011011",
3686 => "0000000000011011",
3687 => "0000000000011011",
3688 => "0000000000011011",
3689 => "0000000000011011",
3690 => "0000000000011011",
3691 => "0000000000011011",
3692 => "0000000000011011",
3693 => "0000000000011011",
3694 => "0000000000011011",
3695 => "0000000000011011",
3696 => "0000000000011011",
3697 => "0000000000011011",
3698 => "0000000000011011",
3699 => "0000000000011011",
3700 => "0000000000011011",
3701 => "0000000000011011",
3702 => "0000000000011011",
3703 => "0000000000011011",
3704 => "0000000000011011",
3705 => "0000000000011011",
3706 => "0000000000011011",
3707 => "0000000000011011",
3708 => "0000000000011011",
3709 => "0000000000011011",
3710 => "0000000000011011",
3711 => "0000000000011011",
3712 => "0000000000011011",
3713 => "0000000000011011",
3714 => "0000000000011011",
3715 => "0000000000011011",
3716 => "0000000000011011",
3717 => "0000000000011011",
3718 => "0000000000011011",
3719 => "0000000000011011",
3720 => "0000000000011011",
3721 => "0000000000011011",
3722 => "0000000000011011",
3723 => "0000000000011011",
3724 => "0000000000011011",
3725 => "0000000000011011",
3726 => "0000000000011011",
3727 => "0000000000011011",
3728 => "0000000000011011",
3729 => "0000000000011011",
3730 => "0000000000011011",
3731 => "0000000000011011",
3732 => "0000000000011011",
3733 => "0000000000011011",
3734 => "0000000000011011",
3735 => "0000000000011011",
3736 => "0000000000011011",
3737 => "0000000000011011",
3738 => "0000000000011011",
3739 => "0000000000011011",
3740 => "0000000000011011",
3741 => "0000000000011011",
3742 => "0000000000011011",
3743 => "0000000000011011",
3744 => "0000000000011011",
3745 => "0000000000011011",
3746 => "0000000000011011",
3747 => "0000000000011011",
3748 => "0000000000011011",
3749 => "0000000000011011",
3750 => "0000000000011011",
3751 => "0000000000011011",
3752 => "0000000000011011",
3753 => "0000000000011011",
3754 => "0000000000011011",
3755 => "0000000000011011",
3756 => "0000000000011011",
3757 => "0000000000011011",
3758 => "0000000000011011",
3759 => "0000000000011011",
3760 => "0000000000011011",
3761 => "0000000000011011",
3762 => "0000000000011011",
3763 => "0000000000011011",
3764 => "0000000000011011",
3765 => "0000000000011011",
3766 => "0000000000011011",
3767 => "0000000000011011",
3768 => "0000000000011011",
3769 => "0000000000011011",
3770 => "0000000000011011",
3771 => "0000000000011011",
3772 => "0000000000011011",
3773 => "0000000000011011",
3774 => "0000000000011011",
3775 => "0000000000011011",
3776 => "0000000000011011",
3777 => "0000000000011011",
3778 => "0000000000011011",
3779 => "0000000000011011",
3780 => "0000000000011011",
3781 => "0000000000011011",
3782 => "0000000000011011",
3783 => "0000000000011011",
3784 => "0000000000011011",
3785 => "0000000000011011",
3786 => "0000000000011011",
3787 => "0000000000011011",
3788 => "0000000000011011",
3789 => "0000000000011011",
3790 => "0000000000011011",
3791 => "0000000000011011",
3792 => "0000000000011011",
3793 => "0000000000011011",
3794 => "0000000000011011",
3795 => "0000000000011011",
3796 => "0000000000011011",
3797 => "0000000000011011",
3798 => "0000000000011011",
3799 => "0000000000011011",
3800 => "0000000000011011",
3801 => "0000000000011011",
3802 => "0000000000011011",
3803 => "0000000000011011",
3804 => "0000000000011011",
3805 => "0000000000011011",
3806 => "0000000000011011",
3807 => "0000000000011011",
3808 => "0000000000011011",
3809 => "0000000000011011",
3810 => "0000000000011011",
3811 => "0000000000011011",
3812 => "0000000000011011",
3813 => "0000000000011011",
3814 => "0000000000011011",
3815 => "0000000000011011",
3816 => "0000000000011011",
3817 => "0000000000011011",
3818 => "0000000000011011",
3819 => "0000000000011011",
3820 => "0000000000011011",
3821 => "0000000000011011",
3822 => "0000000000011011",
3823 => "0000000000011011",
3824 => "0000000000011011",
3825 => "0000000000011011",
3826 => "0000000000011011",
3827 => "0000000000011011",
3828 => "0000000000011011",
3829 => "0000000000011011",
3830 => "0000000000011011",
3831 => "0000000000011011",
3832 => "0000000000011011",
3833 => "0000000000011100",
3834 => "0000000000011100",
3835 => "0000000000011100",
3836 => "0000000000011100",
3837 => "0000000000011100",
3838 => "0000000000011100",
3839 => "0000000000011100",
3840 => "0000000000011100",
3841 => "0000000000011100",
3842 => "0000000000011100",
3843 => "0000000000011100",
3844 => "0000000000011100",
3845 => "0000000000011100",
3846 => "0000000000011100",
3847 => "0000000000011100",
3848 => "0000000000011100",
3849 => "0000000000011100",
3850 => "0000000000011100",
3851 => "0000000000011100",
3852 => "0000000000011100",
3853 => "0000000000011100",
3854 => "0000000000011100",
3855 => "0000000000011100",
3856 => "0000000000011100",
3857 => "0000000000011100",
3858 => "0000000000011100",
3859 => "0000000000011100",
3860 => "0000000000011100",
3861 => "0000000000011100",
3862 => "0000000000011100",
3863 => "0000000000011100",
3864 => "0000000000011100",
3865 => "0000000000011100",
3866 => "0000000000011100",
3867 => "0000000000011100",
3868 => "0000000000011100",
3869 => "0000000000011100",
3870 => "0000000000011100",
3871 => "0000000000011100",
3872 => "0000000000011100",
3873 => "0000000000011100",
3874 => "0000000000011100",
3875 => "0000000000011100",
3876 => "0000000000011100",
3877 => "0000000000011100",
3878 => "0000000000011100",
3879 => "0000000000011100",
3880 => "0000000000011100",
3881 => "0000000000011100",
3882 => "0000000000011100",
3883 => "0000000000011100",
3884 => "0000000000011100",
3885 => "0000000000011100",
3886 => "0000000000011100",
3887 => "0000000000011100",
3888 => "0000000000011100",
3889 => "0000000000011100",
3890 => "0000000000011100",
3891 => "0000000000011100",
3892 => "0000000000011100",
3893 => "0000000000011100",
3894 => "0000000000011100",
3895 => "0000000000011100",
3896 => "0000000000011100",
3897 => "0000000000011100",
3898 => "0000000000011100",
3899 => "0000000000011100",
3900 => "0000000000011100",
3901 => "0000000000011100",
3902 => "0000000000011100",
3903 => "0000000000011100",
3904 => "0000000000011100",
3905 => "0000000000011100",
3906 => "0000000000011100",
3907 => "0000000000011100",
3908 => "0000000000011100",
3909 => "0000000000011100",
3910 => "0000000000011100",
3911 => "0000000000011100",
3912 => "0000000000011100",
3913 => "0000000000011100",
3914 => "0000000000011100",
3915 => "0000000000011100",
3916 => "0000000000011100",
3917 => "0000000000011100",
3918 => "0000000000011100",
3919 => "0000000000011100",
3920 => "0000000000011100",
3921 => "0000000000011100",
3922 => "0000000000011100",
3923 => "0000000000011100",
3924 => "0000000000011100",
3925 => "0000000000011100",
3926 => "0000000000011100",
3927 => "0000000000011100",
3928 => "0000000000011100",
3929 => "0000000000011100",
3930 => "0000000000011100",
3931 => "0000000000011100",
3932 => "0000000000011100",
3933 => "0000000000011100",
3934 => "0000000000011100",
3935 => "0000000000011100",
3936 => "0000000000011100",
3937 => "0000000000011100",
3938 => "0000000000011100",
3939 => "0000000000011100",
3940 => "0000000000011100",
3941 => "0000000000011100",
3942 => "0000000000011100",
3943 => "0000000000011100",
3944 => "0000000000011100",
3945 => "0000000000011100",
3946 => "0000000000011100",
3947 => "0000000000011100",
3948 => "0000000000011100",
3949 => "0000000000011100",
3950 => "0000000000011100",
3951 => "0000000000011100",
3952 => "0000000000011100",
3953 => "0000000000011100",
3954 => "0000000000011100",
3955 => "0000000000011100",
3956 => "0000000000011100",
3957 => "0000000000011100",
3958 => "0000000000011100",
3959 => "0000000000011100",
3960 => "0000000000011100",
3961 => "0000000000011100",
3962 => "0000000000011100",
3963 => "0000000000011100",
3964 => "0000000000011100",
3965 => "0000000000011100",
3966 => "0000000000011100",
3967 => "0000000000011100",
3968 => "0000000000011100",
3969 => "0000000000011100",
3970 => "0000000000011100",
3971 => "0000000000011100",
3972 => "0000000000011100",
3973 => "0000000000011100",
3974 => "0000000000011100",
3975 => "0000000000011100",
3976 => "0000000000011101",
3977 => "0000000000011101",
3978 => "0000000000011101",
3979 => "0000000000011101",
3980 => "0000000000011101",
3981 => "0000000000011101",
3982 => "0000000000011101",
3983 => "0000000000011101",
3984 => "0000000000011101",
3985 => "0000000000011101",
3986 => "0000000000011101",
3987 => "0000000000011101",
3988 => "0000000000011101",
3989 => "0000000000011101",
3990 => "0000000000011101",
3991 => "0000000000011101",
3992 => "0000000000011101",
3993 => "0000000000011101",
3994 => "0000000000011101",
3995 => "0000000000011101",
3996 => "0000000000011101",
3997 => "0000000000011101",
3998 => "0000000000011101",
3999 => "0000000000011101",
4000 => "0000000000011101",
4001 => "0000000000011101",
4002 => "0000000000011101",
4003 => "0000000000011101",
4004 => "0000000000011101",
4005 => "0000000000011101",
4006 => "0000000000011101",
4007 => "0000000000011101",
4008 => "0000000000011101",
4009 => "0000000000011101",
4010 => "0000000000011101",
4011 => "0000000000011101",
4012 => "0000000000011101",
4013 => "0000000000011101",
4014 => "0000000000011101",
4015 => "0000000000011101",
4016 => "0000000000011101",
4017 => "0000000000011101",
4018 => "0000000000011101",
4019 => "0000000000011101",
4020 => "0000000000011101",
4021 => "0000000000011101",
4022 => "0000000000011101",
4023 => "0000000000011101",
4024 => "0000000000011101",
4025 => "0000000000011101",
4026 => "0000000000011101",
4027 => "0000000000011101",
4028 => "0000000000011101",
4029 => "0000000000011101",
4030 => "0000000000011101",
4031 => "0000000000011101",
4032 => "0000000000011101",
4033 => "0000000000011101",
4034 => "0000000000011101",
4035 => "0000000000011101",
4036 => "0000000000011101",
4037 => "0000000000011101",
4038 => "0000000000011101",
4039 => "0000000000011101",
4040 => "0000000000011101",
4041 => "0000000000011101",
4042 => "0000000000011101",
4043 => "0000000000011101",
4044 => "0000000000011101",
4045 => "0000000000011101",
4046 => "0000000000011101",
4047 => "0000000000011101",
4048 => "0000000000011101",
4049 => "0000000000011101",
4050 => "0000000000011101",
4051 => "0000000000011101",
4052 => "0000000000011101",
4053 => "0000000000011101",
4054 => "0000000000011101",
4055 => "0000000000011101",
4056 => "0000000000011101",
4057 => "0000000000011101",
4058 => "0000000000011101",
4059 => "0000000000011101",
4060 => "0000000000011101",
4061 => "0000000000011101",
4062 => "0000000000011101",
4063 => "0000000000011101",
4064 => "0000000000011101",
4065 => "0000000000011101",
4066 => "0000000000011101",
4067 => "0000000000011101",
4068 => "0000000000011101",
4069 => "0000000000011101",
4070 => "0000000000011101",
4071 => "0000000000011101",
4072 => "0000000000011101",
4073 => "0000000000011101",
4074 => "0000000000011101",
4075 => "0000000000011101",
4076 => "0000000000011101",
4077 => "0000000000011101",
4078 => "0000000000011101",
4079 => "0000000000011101",
4080 => "0000000000011101",
4081 => "0000000000011101",
4082 => "0000000000011101",
4083 => "0000000000011101",
4084 => "0000000000011101",
4085 => "0000000000011101",
4086 => "0000000000011101",
4087 => "0000000000011101",
4088 => "0000000000011101",
4089 => "0000000000011101",
4090 => "0000000000011101",
4091 => "0000000000011101",
4092 => "0000000000011101",
4093 => "0000000000011101",
4094 => "0000000000011101",
4095 => "0000000000011101",
4096 => "0000000000011101",
4097 => "0000000000011101",
4098 => "0000000000011101",
4099 => "0000000000011101",
4100 => "0000000000011101",
4101 => "0000000000011101",
4102 => "0000000000011101",
4103 => "0000000000011101",
4104 => "0000000000011101",
4105 => "0000000000011101",
4106 => "0000000000011101",
4107 => "0000000000011101",
4108 => "0000000000011101",
4109 => "0000000000011101",
4110 => "0000000000011101",
4111 => "0000000000011101",
4112 => "0000000000011101",
4113 => "0000000000011101",
4114 => "0000000000011101",
4115 => "0000000000011110",
4116 => "0000000000011110",
4117 => "0000000000011110",
4118 => "0000000000011110",
4119 => "0000000000011110",
4120 => "0000000000011110",
4121 => "0000000000011110",
4122 => "0000000000011110",
4123 => "0000000000011110",
4124 => "0000000000011110",
4125 => "0000000000011110",
4126 => "0000000000011110",
4127 => "0000000000011110",
4128 => "0000000000011110",
4129 => "0000000000011110",
4130 => "0000000000011110",
4131 => "0000000000011110",
4132 => "0000000000011110",
4133 => "0000000000011110",
4134 => "0000000000011110",
4135 => "0000000000011110",
4136 => "0000000000011110",
4137 => "0000000000011110",
4138 => "0000000000011110",
4139 => "0000000000011110",
4140 => "0000000000011110",
4141 => "0000000000011110",
4142 => "0000000000011110",
4143 => "0000000000011110",
4144 => "0000000000011110",
4145 => "0000000000011110",
4146 => "0000000000011110",
4147 => "0000000000011110",
4148 => "0000000000011110",
4149 => "0000000000011110",
4150 => "0000000000011110",
4151 => "0000000000011110",
4152 => "0000000000011110",
4153 => "0000000000011110",
4154 => "0000000000011110",
4155 => "0000000000011110",
4156 => "0000000000011110",
4157 => "0000000000011110",
4158 => "0000000000011110",
4159 => "0000000000011110",
4160 => "0000000000011110",
4161 => "0000000000011110",
4162 => "0000000000011110",
4163 => "0000000000011110",
4164 => "0000000000011110",
4165 => "0000000000011110",
4166 => "0000000000011110",
4167 => "0000000000011110",
4168 => "0000000000011110",
4169 => "0000000000011110",
4170 => "0000000000011110",
4171 => "0000000000011110",
4172 => "0000000000011110",
4173 => "0000000000011110",
4174 => "0000000000011110",
4175 => "0000000000011110",
4176 => "0000000000011110",
4177 => "0000000000011110",
4178 => "0000000000011110",
4179 => "0000000000011110",
4180 => "0000000000011110",
4181 => "0000000000011110",
4182 => "0000000000011110",
4183 => "0000000000011110",
4184 => "0000000000011110",
4185 => "0000000000011110",
4186 => "0000000000011110",
4187 => "0000000000011110",
4188 => "0000000000011110",
4189 => "0000000000011110",
4190 => "0000000000011110",
4191 => "0000000000011110",
4192 => "0000000000011110",
4193 => "0000000000011110",
4194 => "0000000000011110",
4195 => "0000000000011110",
4196 => "0000000000011110",
4197 => "0000000000011110",
4198 => "0000000000011110",
4199 => "0000000000011110",
4200 => "0000000000011110",
4201 => "0000000000011110",
4202 => "0000000000011110",
4203 => "0000000000011110",
4204 => "0000000000011110",
4205 => "0000000000011110",
4206 => "0000000000011110",
4207 => "0000000000011110",
4208 => "0000000000011110",
4209 => "0000000000011110",
4210 => "0000000000011110",
4211 => "0000000000011110",
4212 => "0000000000011110",
4213 => "0000000000011110",
4214 => "0000000000011110",
4215 => "0000000000011110",
4216 => "0000000000011110",
4217 => "0000000000011110",
4218 => "0000000000011110",
4219 => "0000000000011110",
4220 => "0000000000011110",
4221 => "0000000000011110",
4222 => "0000000000011110",
4223 => "0000000000011110",
4224 => "0000000000011110",
4225 => "0000000000011110",
4226 => "0000000000011110",
4227 => "0000000000011110",
4228 => "0000000000011110",
4229 => "0000000000011110",
4230 => "0000000000011110",
4231 => "0000000000011110",
4232 => "0000000000011110",
4233 => "0000000000011110",
4234 => "0000000000011110",
4235 => "0000000000011110",
4236 => "0000000000011110",
4237 => "0000000000011110",
4238 => "0000000000011110",
4239 => "0000000000011110",
4240 => "0000000000011110",
4241 => "0000000000011110",
4242 => "0000000000011110",
4243 => "0000000000011110",
4244 => "0000000000011110",
4245 => "0000000000011110",
4246 => "0000000000011110",
4247 => "0000000000011110",
4248 => "0000000000011110",
4249 => "0000000000011110",
4250 => "0000000000011111",
4251 => "0000000000011111",
4252 => "0000000000011111",
4253 => "0000000000011111",
4254 => "0000000000011111",
4255 => "0000000000011111",
4256 => "0000000000011111",
4257 => "0000000000011111",
4258 => "0000000000011111",
4259 => "0000000000011111",
4260 => "0000000000011111",
4261 => "0000000000011111",
4262 => "0000000000011111",
4263 => "0000000000011111",
4264 => "0000000000011111",
4265 => "0000000000011111",
4266 => "0000000000011111",
4267 => "0000000000011111",
4268 => "0000000000011111",
4269 => "0000000000011111",
4270 => "0000000000011111",
4271 => "0000000000011111",
4272 => "0000000000011111",
4273 => "0000000000011111",
4274 => "0000000000011111",
4275 => "0000000000011111",
4276 => "0000000000011111",
4277 => "0000000000011111",
4278 => "0000000000011111",
4279 => "0000000000011111",
4280 => "0000000000011111",
4281 => "0000000000011111",
4282 => "0000000000011111",
4283 => "0000000000011111",
4284 => "0000000000011111",
4285 => "0000000000011111",
4286 => "0000000000011111",
4287 => "0000000000011111",
4288 => "0000000000011111",
4289 => "0000000000011111",
4290 => "0000000000011111",
4291 => "0000000000011111",
4292 => "0000000000011111",
4293 => "0000000000011111",
4294 => "0000000000011111",
4295 => "0000000000011111",
4296 => "0000000000011111",
4297 => "0000000000011111",
4298 => "0000000000011111",
4299 => "0000000000011111",
4300 => "0000000000011111",
4301 => "0000000000011111",
4302 => "0000000000011111",
4303 => "0000000000011111",
4304 => "0000000000011111",
4305 => "0000000000011111",
4306 => "0000000000011111",
4307 => "0000000000011111",
4308 => "0000000000011111",
4309 => "0000000000011111",
4310 => "0000000000011111",
4311 => "0000000000011111",
4312 => "0000000000011111",
4313 => "0000000000011111",
4314 => "0000000000011111",
4315 => "0000000000011111",
4316 => "0000000000011111",
4317 => "0000000000011111",
4318 => "0000000000011111",
4319 => "0000000000011111",
4320 => "0000000000011111",
4321 => "0000000000011111",
4322 => "0000000000011111",
4323 => "0000000000011111",
4324 => "0000000000011111",
4325 => "0000000000011111",
4326 => "0000000000011111",
4327 => "0000000000011111",
4328 => "0000000000011111",
4329 => "0000000000011111",
4330 => "0000000000011111",
4331 => "0000000000011111",
4332 => "0000000000011111",
4333 => "0000000000011111",
4334 => "0000000000011111",
4335 => "0000000000011111",
4336 => "0000000000011111",
4337 => "0000000000011111",
4338 => "0000000000011111",
4339 => "0000000000011111",
4340 => "0000000000011111",
4341 => "0000000000011111",
4342 => "0000000000011111",
4343 => "0000000000011111",
4344 => "0000000000011111",
4345 => "0000000000011111",
4346 => "0000000000011111",
4347 => "0000000000011111",
4348 => "0000000000011111",
4349 => "0000000000011111",
4350 => "0000000000011111",
4351 => "0000000000011111",
4352 => "0000000000011111",
4353 => "0000000000011111",
4354 => "0000000000011111",
4355 => "0000000000011111",
4356 => "0000000000011111",
4357 => "0000000000011111",
4358 => "0000000000011111",
4359 => "0000000000011111",
4360 => "0000000000011111",
4361 => "0000000000011111",
4362 => "0000000000011111",
4363 => "0000000000011111",
4364 => "0000000000011111",
4365 => "0000000000011111",
4366 => "0000000000011111",
4367 => "0000000000011111",
4368 => "0000000000011111",
4369 => "0000000000011111",
4370 => "0000000000011111",
4371 => "0000000000011111",
4372 => "0000000000011111",
4373 => "0000000000011111",
4374 => "0000000000011111",
4375 => "0000000000011111",
4376 => "0000000000011111",
4377 => "0000000000011111",
4378 => "0000000000011111",
4379 => "0000000000011111",
4380 => "0000000000100000",
4381 => "0000000000100000",
4382 => "0000000000100000",
4383 => "0000000000100000",
4384 => "0000000000100000",
4385 => "0000000000100000",
4386 => "0000000000100000",
4387 => "0000000000100000",
4388 => "0000000000100000",
4389 => "0000000000100000",
4390 => "0000000000100000",
4391 => "0000000000100000",
4392 => "0000000000100000",
4393 => "0000000000100000",
4394 => "0000000000100000",
4395 => "0000000000100000",
4396 => "0000000000100000",
4397 => "0000000000100000",
4398 => "0000000000100000",
4399 => "0000000000100000",
4400 => "0000000000100000",
4401 => "0000000000100000",
4402 => "0000000000100000",
4403 => "0000000000100000",
4404 => "0000000000100000",
4405 => "0000000000100000",
4406 => "0000000000100000",
4407 => "0000000000100000",
4408 => "0000000000100000",
4409 => "0000000000100000",
4410 => "0000000000100000",
4411 => "0000000000100000",
4412 => "0000000000100000",
4413 => "0000000000100000",
4414 => "0000000000100000",
4415 => "0000000000100000",
4416 => "0000000000100000",
4417 => "0000000000100000",
4418 => "0000000000100000",
4419 => "0000000000100000",
4420 => "0000000000100000",
4421 => "0000000000100000",
4422 => "0000000000100000",
4423 => "0000000000100000",
4424 => "0000000000100000",
4425 => "0000000000100000",
4426 => "0000000000100000",
4427 => "0000000000100000",
4428 => "0000000000100000",
4429 => "0000000000100000",
4430 => "0000000000100000",
4431 => "0000000000100000",
4432 => "0000000000100000",
4433 => "0000000000100000",
4434 => "0000000000100000",
4435 => "0000000000100000",
4436 => "0000000000100000",
4437 => "0000000000100000",
4438 => "0000000000100000",
4439 => "0000000000100000",
4440 => "0000000000100000",
4441 => "0000000000100000",
4442 => "0000000000100000",
4443 => "0000000000100000",
4444 => "0000000000100000",
4445 => "0000000000100000",
4446 => "0000000000100000",
4447 => "0000000000100000",
4448 => "0000000000100000",
4449 => "0000000000100000",
4450 => "0000000000100000",
4451 => "0000000000100000",
4452 => "0000000000100000",
4453 => "0000000000100000",
4454 => "0000000000100000",
4455 => "0000000000100000",
4456 => "0000000000100000",
4457 => "0000000000100000",
4458 => "0000000000100000",
4459 => "0000000000100000",
4460 => "0000000000100000",
4461 => "0000000000100000",
4462 => "0000000000100000",
4463 => "0000000000100000",
4464 => "0000000000100000",
4465 => "0000000000100000",
4466 => "0000000000100000",
4467 => "0000000000100000",
4468 => "0000000000100000",
4469 => "0000000000100000",
4470 => "0000000000100000",
4471 => "0000000000100000",
4472 => "0000000000100000",
4473 => "0000000000100000",
4474 => "0000000000100000",
4475 => "0000000000100000",
4476 => "0000000000100000",
4477 => "0000000000100000",
4478 => "0000000000100000",
4479 => "0000000000100000",
4480 => "0000000000100000",
4481 => "0000000000100000",
4482 => "0000000000100000",
4483 => "0000000000100000",
4484 => "0000000000100000",
4485 => "0000000000100000",
4486 => "0000000000100000",
4487 => "0000000000100000",
4488 => "0000000000100000",
4489 => "0000000000100000",
4490 => "0000000000100000",
4491 => "0000000000100000",
4492 => "0000000000100000",
4493 => "0000000000100000",
4494 => "0000000000100000",
4495 => "0000000000100000",
4496 => "0000000000100000",
4497 => "0000000000100000",
4498 => "0000000000100000",
4499 => "0000000000100000",
4500 => "0000000000100000",
4501 => "0000000000100000",
4502 => "0000000000100000",
4503 => "0000000000100000",
4504 => "0000000000100000",
4505 => "0000000000100001",
4506 => "0000000000100001",
4507 => "0000000000100001",
4508 => "0000000000100001",
4509 => "0000000000100001",
4510 => "0000000000100001",
4511 => "0000000000100001",
4512 => "0000000000100001",
4513 => "0000000000100001",
4514 => "0000000000100001",
4515 => "0000000000100001",
4516 => "0000000000100001",
4517 => "0000000000100001",
4518 => "0000000000100001",
4519 => "0000000000100001",
4520 => "0000000000100001",
4521 => "0000000000100001",
4522 => "0000000000100001",
4523 => "0000000000100001",
4524 => "0000000000100001",
4525 => "0000000000100001",
4526 => "0000000000100001",
4527 => "0000000000100001",
4528 => "0000000000100001",
4529 => "0000000000100001",
4530 => "0000000000100001",
4531 => "0000000000100001",
4532 => "0000000000100001",
4533 => "0000000000100001",
4534 => "0000000000100001",
4535 => "0000000000100001",
4536 => "0000000000100001",
4537 => "0000000000100001",
4538 => "0000000000100001",
4539 => "0000000000100001",
4540 => "0000000000100001",
4541 => "0000000000100001",
4542 => "0000000000100001",
4543 => "0000000000100001",
4544 => "0000000000100001",
4545 => "0000000000100001",
4546 => "0000000000100001",
4547 => "0000000000100001",
4548 => "0000000000100001",
4549 => "0000000000100001",
4550 => "0000000000100001",
4551 => "0000000000100001",
4552 => "0000000000100001",
4553 => "0000000000100001",
4554 => "0000000000100001",
4555 => "0000000000100001",
4556 => "0000000000100001",
4557 => "0000000000100001",
4558 => "0000000000100001",
4559 => "0000000000100001",
4560 => "0000000000100001",
4561 => "0000000000100001",
4562 => "0000000000100001",
4563 => "0000000000100001",
4564 => "0000000000100001",
4565 => "0000000000100001",
4566 => "0000000000100001",
4567 => "0000000000100001",
4568 => "0000000000100001",
4569 => "0000000000100001",
4570 => "0000000000100001",
4571 => "0000000000100001",
4572 => "0000000000100001",
4573 => "0000000000100001",
4574 => "0000000000100001",
4575 => "0000000000100001",
4576 => "0000000000100001",
4577 => "0000000000100001",
4578 => "0000000000100001",
4579 => "0000000000100001",
4580 => "0000000000100001",
4581 => "0000000000100001",
4582 => "0000000000100001",
4583 => "0000000000100001",
4584 => "0000000000100001",
4585 => "0000000000100001",
4586 => "0000000000100001",
4587 => "0000000000100001",
4588 => "0000000000100001",
4589 => "0000000000100001",
4590 => "0000000000100001",
4591 => "0000000000100001",
4592 => "0000000000100001",
4593 => "0000000000100001",
4594 => "0000000000100001",
4595 => "0000000000100001",
4596 => "0000000000100001",
4597 => "0000000000100001",
4598 => "0000000000100001",
4599 => "0000000000100001",
4600 => "0000000000100001",
4601 => "0000000000100001",
4602 => "0000000000100001",
4603 => "0000000000100001",
4604 => "0000000000100001",
4605 => "0000000000100001",
4606 => "0000000000100001",
4607 => "0000000000100001",
4608 => "0000000000100001",
4609 => "0000000000100001",
4610 => "0000000000100001",
4611 => "0000000000100001",
4612 => "0000000000100001",
4613 => "0000000000100001",
4614 => "0000000000100001",
4615 => "0000000000100001",
4616 => "0000000000100001",
4617 => "0000000000100001",
4618 => "0000000000100001",
4619 => "0000000000100001",
4620 => "0000000000100001",
4621 => "0000000000100001",
4622 => "0000000000100001",
4623 => "0000000000100001",
4624 => "0000000000100001",
4625 => "0000000000100001",
4626 => "0000000000100001",
4627 => "0000000000100001",
4628 => "0000000000100010",
4629 => "0000000000100010",
4630 => "0000000000100010",
4631 => "0000000000100010",
4632 => "0000000000100010",
4633 => "0000000000100010",
4634 => "0000000000100010",
4635 => "0000000000100010",
4636 => "0000000000100010",
4637 => "0000000000100010",
4638 => "0000000000100010",
4639 => "0000000000100010",
4640 => "0000000000100010",
4641 => "0000000000100010",
4642 => "0000000000100010",
4643 => "0000000000100010",
4644 => "0000000000100010",
4645 => "0000000000100010",
4646 => "0000000000100010",
4647 => "0000000000100010",
4648 => "0000000000100010",
4649 => "0000000000100010",
4650 => "0000000000100010",
4651 => "0000000000100010",
4652 => "0000000000100010",
4653 => "0000000000100010",
4654 => "0000000000100010",
4655 => "0000000000100010",
4656 => "0000000000100010",
4657 => "0000000000100010",
4658 => "0000000000100010",
4659 => "0000000000100010",
4660 => "0000000000100010",
4661 => "0000000000100010",
4662 => "0000000000100010",
4663 => "0000000000100010",
4664 => "0000000000100010",
4665 => "0000000000100010",
4666 => "0000000000100010",
4667 => "0000000000100010",
4668 => "0000000000100010",
4669 => "0000000000100010",
4670 => "0000000000100010",
4671 => "0000000000100010",
4672 => "0000000000100010",
4673 => "0000000000100010",
4674 => "0000000000100010",
4675 => "0000000000100010",
4676 => "0000000000100010",
4677 => "0000000000100010",
4678 => "0000000000100010",
4679 => "0000000000100010",
4680 => "0000000000100010",
4681 => "0000000000100010",
4682 => "0000000000100010",
4683 => "0000000000100010",
4684 => "0000000000100010",
4685 => "0000000000100010",
4686 => "0000000000100010",
4687 => "0000000000100010",
4688 => "0000000000100010",
4689 => "0000000000100010",
4690 => "0000000000100010",
4691 => "0000000000100010",
4692 => "0000000000100010",
4693 => "0000000000100010",
4694 => "0000000000100010",
4695 => "0000000000100010",
4696 => "0000000000100010",
4697 => "0000000000100010",
4698 => "0000000000100010",
4699 => "0000000000100010",
4700 => "0000000000100010",
4701 => "0000000000100010",
4702 => "0000000000100010",
4703 => "0000000000100010",
4704 => "0000000000100010",
4705 => "0000000000100010",
4706 => "0000000000100010",
4707 => "0000000000100010",
4708 => "0000000000100010",
4709 => "0000000000100010",
4710 => "0000000000100010",
4711 => "0000000000100010",
4712 => "0000000000100010",
4713 => "0000000000100010",
4714 => "0000000000100010",
4715 => "0000000000100010",
4716 => "0000000000100010",
4717 => "0000000000100010",
4718 => "0000000000100010",
4719 => "0000000000100010",
4720 => "0000000000100010",
4721 => "0000000000100010",
4722 => "0000000000100010",
4723 => "0000000000100010",
4724 => "0000000000100010",
4725 => "0000000000100010",
4726 => "0000000000100010",
4727 => "0000000000100010",
4728 => "0000000000100010",
4729 => "0000000000100010",
4730 => "0000000000100010",
4731 => "0000000000100010",
4732 => "0000000000100010",
4733 => "0000000000100010",
4734 => "0000000000100010",
4735 => "0000000000100010",
4736 => "0000000000100010",
4737 => "0000000000100010",
4738 => "0000000000100010",
4739 => "0000000000100010",
4740 => "0000000000100010",
4741 => "0000000000100010",
4742 => "0000000000100010",
4743 => "0000000000100010",
4744 => "0000000000100010",
4745 => "0000000000100010",
4746 => "0000000000100010",
4747 => "0000000000100011",
4748 => "0000000000100011",
4749 => "0000000000100011",
4750 => "0000000000100011",
4751 => "0000000000100011",
4752 => "0000000000100011",
4753 => "0000000000100011",
4754 => "0000000000100011",
4755 => "0000000000100011",
4756 => "0000000000100011",
4757 => "0000000000100011",
4758 => "0000000000100011",
4759 => "0000000000100011",
4760 => "0000000000100011",
4761 => "0000000000100011",
4762 => "0000000000100011",
4763 => "0000000000100011",
4764 => "0000000000100011",
4765 => "0000000000100011",
4766 => "0000000000100011",
4767 => "0000000000100011",
4768 => "0000000000100011",
4769 => "0000000000100011",
4770 => "0000000000100011",
4771 => "0000000000100011",
4772 => "0000000000100011",
4773 => "0000000000100011",
4774 => "0000000000100011",
4775 => "0000000000100011",
4776 => "0000000000100011",
4777 => "0000000000100011",
4778 => "0000000000100011",
4779 => "0000000000100011",
4780 => "0000000000100011",
4781 => "0000000000100011",
4782 => "0000000000100011",
4783 => "0000000000100011",
4784 => "0000000000100011",
4785 => "0000000000100011",
4786 => "0000000000100011",
4787 => "0000000000100011",
4788 => "0000000000100011",
4789 => "0000000000100011",
4790 => "0000000000100011",
4791 => "0000000000100011",
4792 => "0000000000100011",
4793 => "0000000000100011",
4794 => "0000000000100011",
4795 => "0000000000100011",
4796 => "0000000000100011",
4797 => "0000000000100011",
4798 => "0000000000100011",
4799 => "0000000000100011",
4800 => "0000000000100011",
4801 => "0000000000100011",
4802 => "0000000000100011",
4803 => "0000000000100011",
4804 => "0000000000100011",
4805 => "0000000000100011",
4806 => "0000000000100011",
4807 => "0000000000100011",
4808 => "0000000000100011",
4809 => "0000000000100011",
4810 => "0000000000100011",
4811 => "0000000000100011",
4812 => "0000000000100011",
4813 => "0000000000100011",
4814 => "0000000000100011",
4815 => "0000000000100011",
4816 => "0000000000100011",
4817 => "0000000000100011",
4818 => "0000000000100011",
4819 => "0000000000100011",
4820 => "0000000000100011",
4821 => "0000000000100011",
4822 => "0000000000100011",
4823 => "0000000000100011",
4824 => "0000000000100011",
4825 => "0000000000100011",
4826 => "0000000000100011",
4827 => "0000000000100011",
4828 => "0000000000100011",
4829 => "0000000000100011",
4830 => "0000000000100011",
4831 => "0000000000100011",
4832 => "0000000000100011",
4833 => "0000000000100011",
4834 => "0000000000100011",
4835 => "0000000000100011",
4836 => "0000000000100011",
4837 => "0000000000100011",
4838 => "0000000000100011",
4839 => "0000000000100011",
4840 => "0000000000100011",
4841 => "0000000000100011",
4842 => "0000000000100011",
4843 => "0000000000100011",
4844 => "0000000000100011",
4845 => "0000000000100011",
4846 => "0000000000100011",
4847 => "0000000000100011",
4848 => "0000000000100011",
4849 => "0000000000100011",
4850 => "0000000000100011",
4851 => "0000000000100011",
4852 => "0000000000100011",
4853 => "0000000000100011",
4854 => "0000000000100011",
4855 => "0000000000100011",
4856 => "0000000000100011",
4857 => "0000000000100011",
4858 => "0000000000100011",
4859 => "0000000000100011",
4860 => "0000000000100011",
4861 => "0000000000100011",
4862 => "0000000000100100",
4863 => "0000000000100100",
4864 => "0000000000100100",
4865 => "0000000000100100",
4866 => "0000000000100100",
4867 => "0000000000100100",
4868 => "0000000000100100",
4869 => "0000000000100100",
4870 => "0000000000100100",
4871 => "0000000000100100",
4872 => "0000000000100100",
4873 => "0000000000100100",
4874 => "0000000000100100",
4875 => "0000000000100100",
4876 => "0000000000100100",
4877 => "0000000000100100",
4878 => "0000000000100100",
4879 => "0000000000100100",
4880 => "0000000000100100",
4881 => "0000000000100100",
4882 => "0000000000100100",
4883 => "0000000000100100",
4884 => "0000000000100100",
4885 => "0000000000100100",
4886 => "0000000000100100",
4887 => "0000000000100100",
4888 => "0000000000100100",
4889 => "0000000000100100",
4890 => "0000000000100100",
4891 => "0000000000100100",
4892 => "0000000000100100",
4893 => "0000000000100100",
4894 => "0000000000100100",
4895 => "0000000000100100",
4896 => "0000000000100100",
4897 => "0000000000100100",
4898 => "0000000000100100",
4899 => "0000000000100100",
4900 => "0000000000100100",
4901 => "0000000000100100",
4902 => "0000000000100100",
4903 => "0000000000100100",
4904 => "0000000000100100",
4905 => "0000000000100100",
4906 => "0000000000100100",
4907 => "0000000000100100",
4908 => "0000000000100100",
4909 => "0000000000100100",
4910 => "0000000000100100",
4911 => "0000000000100100",
4912 => "0000000000100100",
4913 => "0000000000100100",
4914 => "0000000000100100",
4915 => "0000000000100100",
4916 => "0000000000100100",
4917 => "0000000000100100",
4918 => "0000000000100100",
4919 => "0000000000100100",
4920 => "0000000000100100",
4921 => "0000000000100100",
4922 => "0000000000100100",
4923 => "0000000000100100",
4924 => "0000000000100100",
4925 => "0000000000100100",
4926 => "0000000000100100",
4927 => "0000000000100100",
4928 => "0000000000100100",
4929 => "0000000000100100",
4930 => "0000000000100100",
4931 => "0000000000100100",
4932 => "0000000000100100",
4933 => "0000000000100100",
4934 => "0000000000100100",
4935 => "0000000000100100",
4936 => "0000000000100100",
4937 => "0000000000100100",
4938 => "0000000000100100",
4939 => "0000000000100100",
4940 => "0000000000100100",
4941 => "0000000000100100",
4942 => "0000000000100100",
4943 => "0000000000100100",
4944 => "0000000000100100",
4945 => "0000000000100100",
4946 => "0000000000100100",
4947 => "0000000000100100",
4948 => "0000000000100100",
4949 => "0000000000100100",
4950 => "0000000000100100",
4951 => "0000000000100100",
4952 => "0000000000100100",
4953 => "0000000000100100",
4954 => "0000000000100100",
4955 => "0000000000100100",
4956 => "0000000000100100",
4957 => "0000000000100100",
4958 => "0000000000100100",
4959 => "0000000000100100",
4960 => "0000000000100100",
4961 => "0000000000100100",
4962 => "0000000000100100",
4963 => "0000000000100100",
4964 => "0000000000100100",
4965 => "0000000000100100",
4966 => "0000000000100100",
4967 => "0000000000100100",
4968 => "0000000000100100",
4969 => "0000000000100100",
4970 => "0000000000100100",
4971 => "0000000000100100",
4972 => "0000000000100100",
4973 => "0000000000100100",
4974 => "0000000000100100",
4975 => "0000000000100101",
4976 => "0000000000100101",
4977 => "0000000000100101",
4978 => "0000000000100101",
4979 => "0000000000100101",
4980 => "0000000000100101",
4981 => "0000000000100101",
4982 => "0000000000100101",
4983 => "0000000000100101",
4984 => "0000000000100101",
4985 => "0000000000100101",
4986 => "0000000000100101",
4987 => "0000000000100101",
4988 => "0000000000100101",
4989 => "0000000000100101",
4990 => "0000000000100101",
4991 => "0000000000100101",
4992 => "0000000000100101",
4993 => "0000000000100101",
4994 => "0000000000100101",
4995 => "0000000000100101",
4996 => "0000000000100101",
4997 => "0000000000100101",
4998 => "0000000000100101",
4999 => "0000000000100101",
5000 => "0000000000100101",
5001 => "0000000000100101",
5002 => "0000000000100101",
5003 => "0000000000100101",
5004 => "0000000000100101",
5005 => "0000000000100101",
5006 => "0000000000100101",
5007 => "0000000000100101",
5008 => "0000000000100101",
5009 => "0000000000100101",
5010 => "0000000000100101",
5011 => "0000000000100101",
5012 => "0000000000100101",
5013 => "0000000000100101",
5014 => "0000000000100101",
5015 => "0000000000100101",
5016 => "0000000000100101",
5017 => "0000000000100101",
5018 => "0000000000100101",
5019 => "0000000000100101",
5020 => "0000000000100101",
5021 => "0000000000100101",
5022 => "0000000000100101",
5023 => "0000000000100101",
5024 => "0000000000100101",
5025 => "0000000000100101",
5026 => "0000000000100101",
5027 => "0000000000100101",
5028 => "0000000000100101",
5029 => "0000000000100101",
5030 => "0000000000100101",
5031 => "0000000000100101",
5032 => "0000000000100101",
5033 => "0000000000100101",
5034 => "0000000000100101",
5035 => "0000000000100101",
5036 => "0000000000100101",
5037 => "0000000000100101",
5038 => "0000000000100101",
5039 => "0000000000100101",
5040 => "0000000000100101",
5041 => "0000000000100101",
5042 => "0000000000100101",
5043 => "0000000000100101",
5044 => "0000000000100101",
5045 => "0000000000100101",
5046 => "0000000000100101",
5047 => "0000000000100101",
5048 => "0000000000100101",
5049 => "0000000000100101",
5050 => "0000000000100101",
5051 => "0000000000100101",
5052 => "0000000000100101",
5053 => "0000000000100101",
5054 => "0000000000100101",
5055 => "0000000000100101",
5056 => "0000000000100101",
5057 => "0000000000100101",
5058 => "0000000000100101",
5059 => "0000000000100101",
5060 => "0000000000100101",
5061 => "0000000000100101",
5062 => "0000000000100101",
5063 => "0000000000100101",
5064 => "0000000000100101",
5065 => "0000000000100101",
5066 => "0000000000100101",
5067 => "0000000000100101",
5068 => "0000000000100101",
5069 => "0000000000100101",
5070 => "0000000000100101",
5071 => "0000000000100101",
5072 => "0000000000100101",
5073 => "0000000000100101",
5074 => "0000000000100101",
5075 => "0000000000100101",
5076 => "0000000000100101",
5077 => "0000000000100101",
5078 => "0000000000100101",
5079 => "0000000000100101",
5080 => "0000000000100101",
5081 => "0000000000100101",
5082 => "0000000000100101",
5083 => "0000000000100101",
5084 => "0000000000100110",
5085 => "0000000000100110",
5086 => "0000000000100110",
5087 => "0000000000100110",
5088 => "0000000000100110",
5089 => "0000000000100110",
5090 => "0000000000100110",
5091 => "0000000000100110",
5092 => "0000000000100110",
5093 => "0000000000100110",
5094 => "0000000000100110",
5095 => "0000000000100110",
5096 => "0000000000100110",
5097 => "0000000000100110",
5098 => "0000000000100110",
5099 => "0000000000100110",
5100 => "0000000000100110",
5101 => "0000000000100110",
5102 => "0000000000100110",
5103 => "0000000000100110",
5104 => "0000000000100110",
5105 => "0000000000100110",
5106 => "0000000000100110",
5107 => "0000000000100110",
5108 => "0000000000100110",
5109 => "0000000000100110",
5110 => "0000000000100110",
5111 => "0000000000100110",
5112 => "0000000000100110",
5113 => "0000000000100110",
5114 => "0000000000100110",
5115 => "0000000000100110",
5116 => "0000000000100110",
5117 => "0000000000100110",
5118 => "0000000000100110",
5119 => "0000000000100110",
5120 => "0000000000100110",
5121 => "0000000000100110",
5122 => "0000000000100110",
5123 => "0000000000100110",
5124 => "0000000000100110",
5125 => "0000000000100110",
5126 => "0000000000100110",
5127 => "0000000000100110",
5128 => "0000000000100110",
5129 => "0000000000100110",
5130 => "0000000000100110",
5131 => "0000000000100110",
5132 => "0000000000100110",
5133 => "0000000000100110",
5134 => "0000000000100110",
5135 => "0000000000100110",
5136 => "0000000000100110",
5137 => "0000000000100110",
5138 => "0000000000100110",
5139 => "0000000000100110",
5140 => "0000000000100110",
5141 => "0000000000100110",
5142 => "0000000000100110",
5143 => "0000000000100110",
5144 => "0000000000100110",
5145 => "0000000000100110",
5146 => "0000000000100110",
5147 => "0000000000100110",
5148 => "0000000000100110",
5149 => "0000000000100110",
5150 => "0000000000100110",
5151 => "0000000000100110",
5152 => "0000000000100110",
5153 => "0000000000100110",
5154 => "0000000000100110",
5155 => "0000000000100110",
5156 => "0000000000100110",
5157 => "0000000000100110",
5158 => "0000000000100110",
5159 => "0000000000100110",
5160 => "0000000000100110",
5161 => "0000000000100110",
5162 => "0000000000100110",
5163 => "0000000000100110",
5164 => "0000000000100110",
5165 => "0000000000100110",
5166 => "0000000000100110",
5167 => "0000000000100110",
5168 => "0000000000100110",
5169 => "0000000000100110",
5170 => "0000000000100110",
5171 => "0000000000100110",
5172 => "0000000000100110",
5173 => "0000000000100110",
5174 => "0000000000100110",
5175 => "0000000000100110",
5176 => "0000000000100110",
5177 => "0000000000100110",
5178 => "0000000000100110",
5179 => "0000000000100110",
5180 => "0000000000100110",
5181 => "0000000000100110",
5182 => "0000000000100110",
5183 => "0000000000100110",
5184 => "0000000000100110",
5185 => "0000000000100110",
5186 => "0000000000100110",
5187 => "0000000000100110",
5188 => "0000000000100110",
5189 => "0000000000100110",
5190 => "0000000000100110",
5191 => "0000000000100111",
5192 => "0000000000100111",
5193 => "0000000000100111",
5194 => "0000000000100111",
5195 => "0000000000100111",
5196 => "0000000000100111",
5197 => "0000000000100111",
5198 => "0000000000100111",
5199 => "0000000000100111",
5200 => "0000000000100111",
5201 => "0000000000100111",
5202 => "0000000000100111",
5203 => "0000000000100111",
5204 => "0000000000100111",
5205 => "0000000000100111",
5206 => "0000000000100111",
5207 => "0000000000100111",
5208 => "0000000000100111",
5209 => "0000000000100111",
5210 => "0000000000100111",
5211 => "0000000000100111",
5212 => "0000000000100111",
5213 => "0000000000100111",
5214 => "0000000000100111",
5215 => "0000000000100111",
5216 => "0000000000100111",
5217 => "0000000000100111",
5218 => "0000000000100111",
5219 => "0000000000100111",
5220 => "0000000000100111",
5221 => "0000000000100111",
5222 => "0000000000100111",
5223 => "0000000000100111",
5224 => "0000000000100111",
5225 => "0000000000100111",
5226 => "0000000000100111",
5227 => "0000000000100111",
5228 => "0000000000100111",
5229 => "0000000000100111",
5230 => "0000000000100111",
5231 => "0000000000100111",
5232 => "0000000000100111",
5233 => "0000000000100111",
5234 => "0000000000100111",
5235 => "0000000000100111",
5236 => "0000000000100111",
5237 => "0000000000100111",
5238 => "0000000000100111",
5239 => "0000000000100111",
5240 => "0000000000100111",
5241 => "0000000000100111",
5242 => "0000000000100111",
5243 => "0000000000100111",
5244 => "0000000000100111",
5245 => "0000000000100111",
5246 => "0000000000100111",
5247 => "0000000000100111",
5248 => "0000000000100111",
5249 => "0000000000100111",
5250 => "0000000000100111",
5251 => "0000000000100111",
5252 => "0000000000100111",
5253 => "0000000000100111",
5254 => "0000000000100111",
5255 => "0000000000100111",
5256 => "0000000000100111",
5257 => "0000000000100111",
5258 => "0000000000100111",
5259 => "0000000000100111",
5260 => "0000000000100111",
5261 => "0000000000100111",
5262 => "0000000000100111",
5263 => "0000000000100111",
5264 => "0000000000100111",
5265 => "0000000000100111",
5266 => "0000000000100111",
5267 => "0000000000100111",
5268 => "0000000000100111",
5269 => "0000000000100111",
5270 => "0000000000100111",
5271 => "0000000000100111",
5272 => "0000000000100111",
5273 => "0000000000100111",
5274 => "0000000000100111",
5275 => "0000000000100111",
5276 => "0000000000100111",
5277 => "0000000000100111",
5278 => "0000000000100111",
5279 => "0000000000100111",
5280 => "0000000000100111",
5281 => "0000000000100111",
5282 => "0000000000100111",
5283 => "0000000000100111",
5284 => "0000000000100111",
5285 => "0000000000100111",
5286 => "0000000000100111",
5287 => "0000000000100111",
5288 => "0000000000100111",
5289 => "0000000000100111",
5290 => "0000000000100111",
5291 => "0000000000100111",
5292 => "0000000000100111",
5293 => "0000000000100111",
5294 => "0000000000100111",
5295 => "0000000000101000",
5296 => "0000000000101000",
5297 => "0000000000101000",
5298 => "0000000000101000",
5299 => "0000000000101000",
5300 => "0000000000101000",
5301 => "0000000000101000",
5302 => "0000000000101000",
5303 => "0000000000101000",
5304 => "0000000000101000",
5305 => "0000000000101000",
5306 => "0000000000101000",
5307 => "0000000000101000",
5308 => "0000000000101000",
5309 => "0000000000101000",
5310 => "0000000000101000",
5311 => "0000000000101000",
5312 => "0000000000101000",
5313 => "0000000000101000",
5314 => "0000000000101000",
5315 => "0000000000101000",
5316 => "0000000000101000",
5317 => "0000000000101000",
5318 => "0000000000101000",
5319 => "0000000000101000",
5320 => "0000000000101000",
5321 => "0000000000101000",
5322 => "0000000000101000",
5323 => "0000000000101000",
5324 => "0000000000101000",
5325 => "0000000000101000",
5326 => "0000000000101000",
5327 => "0000000000101000",
5328 => "0000000000101000",
5329 => "0000000000101000",
5330 => "0000000000101000",
5331 => "0000000000101000",
5332 => "0000000000101000",
5333 => "0000000000101000",
5334 => "0000000000101000",
5335 => "0000000000101000",
5336 => "0000000000101000",
5337 => "0000000000101000",
5338 => "0000000000101000",
5339 => "0000000000101000",
5340 => "0000000000101000",
5341 => "0000000000101000",
5342 => "0000000000101000",
5343 => "0000000000101000",
5344 => "0000000000101000",
5345 => "0000000000101000",
5346 => "0000000000101000",
5347 => "0000000000101000",
5348 => "0000000000101000",
5349 => "0000000000101000",
5350 => "0000000000101000",
5351 => "0000000000101000",
5352 => "0000000000101000",
5353 => "0000000000101000",
5354 => "0000000000101000",
5355 => "0000000000101000",
5356 => "0000000000101000",
5357 => "0000000000101000",
5358 => "0000000000101000",
5359 => "0000000000101000",
5360 => "0000000000101000",
5361 => "0000000000101000",
5362 => "0000000000101000",
5363 => "0000000000101000",
5364 => "0000000000101000",
5365 => "0000000000101000",
5366 => "0000000000101000",
5367 => "0000000000101000",
5368 => "0000000000101000",
5369 => "0000000000101000",
5370 => "0000000000101000",
5371 => "0000000000101000",
5372 => "0000000000101000",
5373 => "0000000000101000",
5374 => "0000000000101000",
5375 => "0000000000101000",
5376 => "0000000000101000",
5377 => "0000000000101000",
5378 => "0000000000101000",
5379 => "0000000000101000",
5380 => "0000000000101000",
5381 => "0000000000101000",
5382 => "0000000000101000",
5383 => "0000000000101000",
5384 => "0000000000101000",
5385 => "0000000000101000",
5386 => "0000000000101000",
5387 => "0000000000101000",
5388 => "0000000000101000",
5389 => "0000000000101000",
5390 => "0000000000101000",
5391 => "0000000000101000",
5392 => "0000000000101000",
5393 => "0000000000101000",
5394 => "0000000000101000",
5395 => "0000000000101000",
5396 => "0000000000101001",
5397 => "0000000000101001",
5398 => "0000000000101001",
5399 => "0000000000101001",
5400 => "0000000000101001",
5401 => "0000000000101001",
5402 => "0000000000101001",
5403 => "0000000000101001",
5404 => "0000000000101001",
5405 => "0000000000101001",
5406 => "0000000000101001",
5407 => "0000000000101001",
5408 => "0000000000101001",
5409 => "0000000000101001",
5410 => "0000000000101001",
5411 => "0000000000101001",
5412 => "0000000000101001",
5413 => "0000000000101001",
5414 => "0000000000101001",
5415 => "0000000000101001",
5416 => "0000000000101001",
5417 => "0000000000101001",
5418 => "0000000000101001",
5419 => "0000000000101001",
5420 => "0000000000101001",
5421 => "0000000000101001",
5422 => "0000000000101001",
5423 => "0000000000101001",
5424 => "0000000000101001",
5425 => "0000000000101001",
5426 => "0000000000101001",
5427 => "0000000000101001",
5428 => "0000000000101001",
5429 => "0000000000101001",
5430 => "0000000000101001",
5431 => "0000000000101001",
5432 => "0000000000101001",
5433 => "0000000000101001",
5434 => "0000000000101001",
5435 => "0000000000101001",
5436 => "0000000000101001",
5437 => "0000000000101001",
5438 => "0000000000101001",
5439 => "0000000000101001",
5440 => "0000000000101001",
5441 => "0000000000101001",
5442 => "0000000000101001",
5443 => "0000000000101001",
5444 => "0000000000101001",
5445 => "0000000000101001",
5446 => "0000000000101001",
5447 => "0000000000101001",
5448 => "0000000000101001",
5449 => "0000000000101001",
5450 => "0000000000101001",
5451 => "0000000000101001",
5452 => "0000000000101001",
5453 => "0000000000101001",
5454 => "0000000000101001",
5455 => "0000000000101001",
5456 => "0000000000101001",
5457 => "0000000000101001",
5458 => "0000000000101001",
5459 => "0000000000101001",
5460 => "0000000000101001",
5461 => "0000000000101001",
5462 => "0000000000101001",
5463 => "0000000000101001",
5464 => "0000000000101001",
5465 => "0000000000101001",
5466 => "0000000000101001",
5467 => "0000000000101001",
5468 => "0000000000101001",
5469 => "0000000000101001",
5470 => "0000000000101001",
5471 => "0000000000101001",
5472 => "0000000000101001",
5473 => "0000000000101001",
5474 => "0000000000101001",
5475 => "0000000000101001",
5476 => "0000000000101001",
5477 => "0000000000101001",
5478 => "0000000000101001",
5479 => "0000000000101001",
5480 => "0000000000101001",
5481 => "0000000000101001",
5482 => "0000000000101001",
5483 => "0000000000101001",
5484 => "0000000000101001",
5485 => "0000000000101001",
5486 => "0000000000101001",
5487 => "0000000000101001",
5488 => "0000000000101001",
5489 => "0000000000101001",
5490 => "0000000000101001",
5491 => "0000000000101001",
5492 => "0000000000101001",
5493 => "0000000000101001",
5494 => "0000000000101001",
5495 => "0000000000101010",
5496 => "0000000000101010",
5497 => "0000000000101010",
5498 => "0000000000101010",
5499 => "0000000000101010",
5500 => "0000000000101010",
5501 => "0000000000101010",
5502 => "0000000000101010",
5503 => "0000000000101010",
5504 => "0000000000101010",
5505 => "0000000000101010",
5506 => "0000000000101010",
5507 => "0000000000101010",
5508 => "0000000000101010",
5509 => "0000000000101010",
5510 => "0000000000101010",
5511 => "0000000000101010",
5512 => "0000000000101010",
5513 => "0000000000101010",
5514 => "0000000000101010",
5515 => "0000000000101010",
5516 => "0000000000101010",
5517 => "0000000000101010",
5518 => "0000000000101010",
5519 => "0000000000101010",
5520 => "0000000000101010",
5521 => "0000000000101010",
5522 => "0000000000101010",
5523 => "0000000000101010",
5524 => "0000000000101010",
5525 => "0000000000101010",
5526 => "0000000000101010",
5527 => "0000000000101010",
5528 => "0000000000101010",
5529 => "0000000000101010",
5530 => "0000000000101010",
5531 => "0000000000101010",
5532 => "0000000000101010",
5533 => "0000000000101010",
5534 => "0000000000101010",
5535 => "0000000000101010",
5536 => "0000000000101010",
5537 => "0000000000101010",
5538 => "0000000000101010",
5539 => "0000000000101010",
5540 => "0000000000101010",
5541 => "0000000000101010",
5542 => "0000000000101010",
5543 => "0000000000101010",
5544 => "0000000000101010",
5545 => "0000000000101010",
5546 => "0000000000101010",
5547 => "0000000000101010",
5548 => "0000000000101010",
5549 => "0000000000101010",
5550 => "0000000000101010",
5551 => "0000000000101010",
5552 => "0000000000101010",
5553 => "0000000000101010",
5554 => "0000000000101010",
5555 => "0000000000101010",
5556 => "0000000000101010",
5557 => "0000000000101010",
5558 => "0000000000101010",
5559 => "0000000000101010",
5560 => "0000000000101010",
5561 => "0000000000101010",
5562 => "0000000000101010",
5563 => "0000000000101010",
5564 => "0000000000101010",
5565 => "0000000000101010",
5566 => "0000000000101010",
5567 => "0000000000101010",
5568 => "0000000000101010",
5569 => "0000000000101010",
5570 => "0000000000101010",
5571 => "0000000000101010",
5572 => "0000000000101010",
5573 => "0000000000101010",
5574 => "0000000000101010",
5575 => "0000000000101010",
5576 => "0000000000101010",
5577 => "0000000000101010",
5578 => "0000000000101010",
5579 => "0000000000101010",
5580 => "0000000000101010",
5581 => "0000000000101010",
5582 => "0000000000101010",
5583 => "0000000000101010",
5584 => "0000000000101010",
5585 => "0000000000101010",
5586 => "0000000000101010",
5587 => "0000000000101010",
5588 => "0000000000101010",
5589 => "0000000000101010",
5590 => "0000000000101010",
5591 => "0000000000101011",
5592 => "0000000000101011",
5593 => "0000000000101011",
5594 => "0000000000101011",
5595 => "0000000000101011",
5596 => "0000000000101011",
5597 => "0000000000101011",
5598 => "0000000000101011",
5599 => "0000000000101011",
5600 => "0000000000101011",
5601 => "0000000000101011",
5602 => "0000000000101011",
5603 => "0000000000101011",
5604 => "0000000000101011",
5605 => "0000000000101011",
5606 => "0000000000101011",
5607 => "0000000000101011",
5608 => "0000000000101011",
5609 => "0000000000101011",
5610 => "0000000000101011",
5611 => "0000000000101011",
5612 => "0000000000101011",
5613 => "0000000000101011",
5614 => "0000000000101011",
5615 => "0000000000101011",
5616 => "0000000000101011",
5617 => "0000000000101011",
5618 => "0000000000101011",
5619 => "0000000000101011",
5620 => "0000000000101011",
5621 => "0000000000101011",
5622 => "0000000000101011",
5623 => "0000000000101011",
5624 => "0000000000101011",
5625 => "0000000000101011",
5626 => "0000000000101011",
5627 => "0000000000101011",
5628 => "0000000000101011",
5629 => "0000000000101011",
5630 => "0000000000101011",
5631 => "0000000000101011",
5632 => "0000000000101011",
5633 => "0000000000101011",
5634 => "0000000000101011",
5635 => "0000000000101011",
5636 => "0000000000101011",
5637 => "0000000000101011",
5638 => "0000000000101011",
5639 => "0000000000101011",
5640 => "0000000000101011",
5641 => "0000000000101011",
5642 => "0000000000101011",
5643 => "0000000000101011",
5644 => "0000000000101011",
5645 => "0000000000101011",
5646 => "0000000000101011",
5647 => "0000000000101011",
5648 => "0000000000101011",
5649 => "0000000000101011",
5650 => "0000000000101011",
5651 => "0000000000101011",
5652 => "0000000000101011",
5653 => "0000000000101011",
5654 => "0000000000101011",
5655 => "0000000000101011",
5656 => "0000000000101011",
5657 => "0000000000101011",
5658 => "0000000000101011",
5659 => "0000000000101011",
5660 => "0000000000101011",
5661 => "0000000000101011",
5662 => "0000000000101011",
5663 => "0000000000101011",
5664 => "0000000000101011",
5665 => "0000000000101011",
5666 => "0000000000101011",
5667 => "0000000000101011",
5668 => "0000000000101011",
5669 => "0000000000101011",
5670 => "0000000000101011",
5671 => "0000000000101011",
5672 => "0000000000101011",
5673 => "0000000000101011",
5674 => "0000000000101011",
5675 => "0000000000101011",
5676 => "0000000000101011",
5677 => "0000000000101011",
5678 => "0000000000101011",
5679 => "0000000000101011",
5680 => "0000000000101011",
5681 => "0000000000101011",
5682 => "0000000000101011",
5683 => "0000000000101011",
5684 => "0000000000101011",
5685 => "0000000000101011",
5686 => "0000000000101100",
5687 => "0000000000101100",
5688 => "0000000000101100",
5689 => "0000000000101100",
5690 => "0000000000101100",
5691 => "0000000000101100",
5692 => "0000000000101100",
5693 => "0000000000101100",
5694 => "0000000000101100",
5695 => "0000000000101100",
5696 => "0000000000101100",
5697 => "0000000000101100",
5698 => "0000000000101100",
5699 => "0000000000101100",
5700 => "0000000000101100",
5701 => "0000000000101100",
5702 => "0000000000101100",
5703 => "0000000000101100",
5704 => "0000000000101100",
5705 => "0000000000101100",
5706 => "0000000000101100",
5707 => "0000000000101100",
5708 => "0000000000101100",
5709 => "0000000000101100",
5710 => "0000000000101100",
5711 => "0000000000101100",
5712 => "0000000000101100",
5713 => "0000000000101100",
5714 => "0000000000101100",
5715 => "0000000000101100",
5716 => "0000000000101100",
5717 => "0000000000101100",
5718 => "0000000000101100",
5719 => "0000000000101100",
5720 => "0000000000101100",
5721 => "0000000000101100",
5722 => "0000000000101100",
5723 => "0000000000101100",
5724 => "0000000000101100",
5725 => "0000000000101100",
5726 => "0000000000101100",
5727 => "0000000000101100",
5728 => "0000000000101100",
5729 => "0000000000101100",
5730 => "0000000000101100",
5731 => "0000000000101100",
5732 => "0000000000101100",
5733 => "0000000000101100",
5734 => "0000000000101100",
5735 => "0000000000101100",
5736 => "0000000000101100",
5737 => "0000000000101100",
5738 => "0000000000101100",
5739 => "0000000000101100",
5740 => "0000000000101100",
5741 => "0000000000101100",
5742 => "0000000000101100",
5743 => "0000000000101100",
5744 => "0000000000101100",
5745 => "0000000000101100",
5746 => "0000000000101100",
5747 => "0000000000101100",
5748 => "0000000000101100",
5749 => "0000000000101100",
5750 => "0000000000101100",
5751 => "0000000000101100",
5752 => "0000000000101100",
5753 => "0000000000101100",
5754 => "0000000000101100",
5755 => "0000000000101100",
5756 => "0000000000101100",
5757 => "0000000000101100",
5758 => "0000000000101100",
5759 => "0000000000101100",
5760 => "0000000000101100",
5761 => "0000000000101100",
5762 => "0000000000101100",
5763 => "0000000000101100",
5764 => "0000000000101100",
5765 => "0000000000101100",
5766 => "0000000000101100",
5767 => "0000000000101100",
5768 => "0000000000101100",
5769 => "0000000000101100",
5770 => "0000000000101100",
5771 => "0000000000101100",
5772 => "0000000000101100",
5773 => "0000000000101100",
5774 => "0000000000101100",
5775 => "0000000000101100",
5776 => "0000000000101100",
5777 => "0000000000101100",
5778 => "0000000000101101",
5779 => "0000000000101101",
5780 => "0000000000101101",
5781 => "0000000000101101",
5782 => "0000000000101101",
5783 => "0000000000101101",
5784 => "0000000000101101",
5785 => "0000000000101101",
5786 => "0000000000101101",
5787 => "0000000000101101",
5788 => "0000000000101101",
5789 => "0000000000101101",
5790 => "0000000000101101",
5791 => "0000000000101101",
5792 => "0000000000101101",
5793 => "0000000000101101",
5794 => "0000000000101101",
5795 => "0000000000101101",
5796 => "0000000000101101",
5797 => "0000000000101101",
5798 => "0000000000101101",
5799 => "0000000000101101",
5800 => "0000000000101101",
5801 => "0000000000101101",
5802 => "0000000000101101",
5803 => "0000000000101101",
5804 => "0000000000101101",
5805 => "0000000000101101",
5806 => "0000000000101101",
5807 => "0000000000101101",
5808 => "0000000000101101",
5809 => "0000000000101101",
5810 => "0000000000101101",
5811 => "0000000000101101",
5812 => "0000000000101101",
5813 => "0000000000101101",
5814 => "0000000000101101",
5815 => "0000000000101101",
5816 => "0000000000101101",
5817 => "0000000000101101",
5818 => "0000000000101101",
5819 => "0000000000101101",
5820 => "0000000000101101",
5821 => "0000000000101101",
5822 => "0000000000101101",
5823 => "0000000000101101",
5824 => "0000000000101101",
5825 => "0000000000101101",
5826 => "0000000000101101",
5827 => "0000000000101101",
5828 => "0000000000101101",
5829 => "0000000000101101",
5830 => "0000000000101101",
5831 => "0000000000101101",
5832 => "0000000000101101",
5833 => "0000000000101101",
5834 => "0000000000101101",
5835 => "0000000000101101",
5836 => "0000000000101101",
5837 => "0000000000101101",
5838 => "0000000000101101",
5839 => "0000000000101101",
5840 => "0000000000101101",
5841 => "0000000000101101",
5842 => "0000000000101101",
5843 => "0000000000101101",
5844 => "0000000000101101",
5845 => "0000000000101101",
5846 => "0000000000101101",
5847 => "0000000000101101",
5848 => "0000000000101101",
5849 => "0000000000101101",
5850 => "0000000000101101",
5851 => "0000000000101101",
5852 => "0000000000101101",
5853 => "0000000000101101",
5854 => "0000000000101101",
5855 => "0000000000101101",
5856 => "0000000000101101",
5857 => "0000000000101101",
5858 => "0000000000101101",
5859 => "0000000000101101",
5860 => "0000000000101101",
5861 => "0000000000101101",
5862 => "0000000000101101",
5863 => "0000000000101101",
5864 => "0000000000101101",
5865 => "0000000000101101",
5866 => "0000000000101101",
5867 => "0000000000101101",
5868 => "0000000000101110",
5869 => "0000000000101110",
5870 => "0000000000101110",
5871 => "0000000000101110",
5872 => "0000000000101110",
5873 => "0000000000101110",
5874 => "0000000000101110",
5875 => "0000000000101110",
5876 => "0000000000101110",
5877 => "0000000000101110",
5878 => "0000000000101110",
5879 => "0000000000101110",
5880 => "0000000000101110",
5881 => "0000000000101110",
5882 => "0000000000101110",
5883 => "0000000000101110",
5884 => "0000000000101110",
5885 => "0000000000101110",
5886 => "0000000000101110",
5887 => "0000000000101110",
5888 => "0000000000101110",
5889 => "0000000000101110",
5890 => "0000000000101110",
5891 => "0000000000101110",
5892 => "0000000000101110",
5893 => "0000000000101110",
5894 => "0000000000101110",
5895 => "0000000000101110",
5896 => "0000000000101110",
5897 => "0000000000101110",
5898 => "0000000000101110",
5899 => "0000000000101110",
5900 => "0000000000101110",
5901 => "0000000000101110",
5902 => "0000000000101110",
5903 => "0000000000101110",
5904 => "0000000000101110",
5905 => "0000000000101110",
5906 => "0000000000101110",
5907 => "0000000000101110",
5908 => "0000000000101110",
5909 => "0000000000101110",
5910 => "0000000000101110",
5911 => "0000000000101110",
5912 => "0000000000101110",
5913 => "0000000000101110",
5914 => "0000000000101110",
5915 => "0000000000101110",
5916 => "0000000000101110",
5917 => "0000000000101110",
5918 => "0000000000101110",
5919 => "0000000000101110",
5920 => "0000000000101110",
5921 => "0000000000101110",
5922 => "0000000000101110",
5923 => "0000000000101110",
5924 => "0000000000101110",
5925 => "0000000000101110",
5926 => "0000000000101110",
5927 => "0000000000101110",
5928 => "0000000000101110",
5929 => "0000000000101110",
5930 => "0000000000101110",
5931 => "0000000000101110",
5932 => "0000000000101110",
5933 => "0000000000101110",
5934 => "0000000000101110",
5935 => "0000000000101110",
5936 => "0000000000101110",
5937 => "0000000000101110",
5938 => "0000000000101110",
5939 => "0000000000101110",
5940 => "0000000000101110",
5941 => "0000000000101110",
5942 => "0000000000101110",
5943 => "0000000000101110",
5944 => "0000000000101110",
5945 => "0000000000101110",
5946 => "0000000000101110",
5947 => "0000000000101110",
5948 => "0000000000101110",
5949 => "0000000000101110",
5950 => "0000000000101110",
5951 => "0000000000101110",
5952 => "0000000000101110",
5953 => "0000000000101110",
5954 => "0000000000101110",
5955 => "0000000000101110",
5956 => "0000000000101111",
5957 => "0000000000101111",
5958 => "0000000000101111",
5959 => "0000000000101111",
5960 => "0000000000101111",
5961 => "0000000000101111",
5962 => "0000000000101111",
5963 => "0000000000101111",
5964 => "0000000000101111",
5965 => "0000000000101111",
5966 => "0000000000101111",
5967 => "0000000000101111",
5968 => "0000000000101111",
5969 => "0000000000101111",
5970 => "0000000000101111",
5971 => "0000000000101111",
5972 => "0000000000101111",
5973 => "0000000000101111",
5974 => "0000000000101111",
5975 => "0000000000101111",
5976 => "0000000000101111",
5977 => "0000000000101111",
5978 => "0000000000101111",
5979 => "0000000000101111",
5980 => "0000000000101111",
5981 => "0000000000101111",
5982 => "0000000000101111",
5983 => "0000000000101111",
5984 => "0000000000101111",
5985 => "0000000000101111",
5986 => "0000000000101111",
5987 => "0000000000101111",
5988 => "0000000000101111",
5989 => "0000000000101111",
5990 => "0000000000101111",
5991 => "0000000000101111",
5992 => "0000000000101111",
5993 => "0000000000101111",
5994 => "0000000000101111",
5995 => "0000000000101111",
5996 => "0000000000101111",
5997 => "0000000000101111",
5998 => "0000000000101111",
5999 => "0000000000101111",
6000 => "0000000000101111",
6001 => "0000000000101111",
6002 => "0000000000101111",
6003 => "0000000000101111",
6004 => "0000000000101111",
6005 => "0000000000101111",
6006 => "0000000000101111",
6007 => "0000000000101111",
6008 => "0000000000101111",
6009 => "0000000000101111",
6010 => "0000000000101111",
6011 => "0000000000101111",
6012 => "0000000000101111",
6013 => "0000000000101111",
6014 => "0000000000101111",
6015 => "0000000000101111",
6016 => "0000000000101111",
6017 => "0000000000101111",
6018 => "0000000000101111",
6019 => "0000000000101111",
6020 => "0000000000101111",
6021 => "0000000000101111",
6022 => "0000000000101111",
6023 => "0000000000101111",
6024 => "0000000000101111",
6025 => "0000000000101111",
6026 => "0000000000101111",
6027 => "0000000000101111",
6028 => "0000000000101111",
6029 => "0000000000101111",
6030 => "0000000000101111",
6031 => "0000000000101111",
6032 => "0000000000101111",
6033 => "0000000000101111",
6034 => "0000000000101111",
6035 => "0000000000101111",
6036 => "0000000000101111",
6037 => "0000000000101111",
6038 => "0000000000101111",
6039 => "0000000000101111",
6040 => "0000000000101111",
6041 => "0000000000101111",
6042 => "0000000000101111",
6043 => "0000000000110000",
6044 => "0000000000110000",
6045 => "0000000000110000",
6046 => "0000000000110000",
6047 => "0000000000110000",
6048 => "0000000000110000",
6049 => "0000000000110000",
6050 => "0000000000110000",
6051 => "0000000000110000",
6052 => "0000000000110000",
6053 => "0000000000110000",
6054 => "0000000000110000",
6055 => "0000000000110000",
6056 => "0000000000110000",
6057 => "0000000000110000",
6058 => "0000000000110000",
6059 => "0000000000110000",
6060 => "0000000000110000",
6061 => "0000000000110000",
6062 => "0000000000110000",
6063 => "0000000000110000",
6064 => "0000000000110000",
6065 => "0000000000110000",
6066 => "0000000000110000",
6067 => "0000000000110000",
6068 => "0000000000110000",
6069 => "0000000000110000",
6070 => "0000000000110000",
6071 => "0000000000110000",
6072 => "0000000000110000",
6073 => "0000000000110000",
6074 => "0000000000110000",
6075 => "0000000000110000",
6076 => "0000000000110000",
6077 => "0000000000110000",
6078 => "0000000000110000",
6079 => "0000000000110000",
6080 => "0000000000110000",
6081 => "0000000000110000",
6082 => "0000000000110000",
6083 => "0000000000110000",
6084 => "0000000000110000",
6085 => "0000000000110000",
6086 => "0000000000110000",
6087 => "0000000000110000",
6088 => "0000000000110000",
6089 => "0000000000110000",
6090 => "0000000000110000",
6091 => "0000000000110000",
6092 => "0000000000110000",
6093 => "0000000000110000",
6094 => "0000000000110000",
6095 => "0000000000110000",
6096 => "0000000000110000",
6097 => "0000000000110000",
6098 => "0000000000110000",
6099 => "0000000000110000",
6100 => "0000000000110000",
6101 => "0000000000110000",
6102 => "0000000000110000",
6103 => "0000000000110000",
6104 => "0000000000110000",
6105 => "0000000000110000",
6106 => "0000000000110000",
6107 => "0000000000110000",
6108 => "0000000000110000",
6109 => "0000000000110000",
6110 => "0000000000110000",
6111 => "0000000000110000",
6112 => "0000000000110000",
6113 => "0000000000110000",
6114 => "0000000000110000",
6115 => "0000000000110000",
6116 => "0000000000110000",
6117 => "0000000000110000",
6118 => "0000000000110000",
6119 => "0000000000110000",
6120 => "0000000000110000",
6121 => "0000000000110000",
6122 => "0000000000110000",
6123 => "0000000000110000",
6124 => "0000000000110000",
6125 => "0000000000110000",
6126 => "0000000000110000",
6127 => "0000000000110001",
6128 => "0000000000110001",
6129 => "0000000000110001",
6130 => "0000000000110001",
6131 => "0000000000110001",
6132 => "0000000000110001",
6133 => "0000000000110001",
6134 => "0000000000110001",
6135 => "0000000000110001",
6136 => "0000000000110001",
6137 => "0000000000110001",
6138 => "0000000000110001",
6139 => "0000000000110001",
6140 => "0000000000110001",
6141 => "0000000000110001",
6142 => "0000000000110001",
6143 => "0000000000110001",
6144 => "0000000000110001",
6145 => "0000000000110001",
6146 => "0000000000110001",
6147 => "0000000000110001",
6148 => "0000000000110001",
6149 => "0000000000110001",
6150 => "0000000000110001",
6151 => "0000000000110001",
6152 => "0000000000110001",
6153 => "0000000000110001",
6154 => "0000000000110001",
6155 => "0000000000110001",
6156 => "0000000000110001",
6157 => "0000000000110001",
6158 => "0000000000110001",
6159 => "0000000000110001",
6160 => "0000000000110001",
6161 => "0000000000110001",
6162 => "0000000000110001",
6163 => "0000000000110001",
6164 => "0000000000110001",
6165 => "0000000000110001",
6166 => "0000000000110001",
6167 => "0000000000110001",
6168 => "0000000000110001",
6169 => "0000000000110001",
6170 => "0000000000110001",
6171 => "0000000000110001",
6172 => "0000000000110001",
6173 => "0000000000110001",
6174 => "0000000000110001",
6175 => "0000000000110001",
6176 => "0000000000110001",
6177 => "0000000000110001",
6178 => "0000000000110001",
6179 => "0000000000110001",
6180 => "0000000000110001",
6181 => "0000000000110001",
6182 => "0000000000110001",
6183 => "0000000000110001",
6184 => "0000000000110001",
6185 => "0000000000110001",
6186 => "0000000000110001",
6187 => "0000000000110001",
6188 => "0000000000110001",
6189 => "0000000000110001",
6190 => "0000000000110001",
6191 => "0000000000110001",
6192 => "0000000000110001",
6193 => "0000000000110001",
6194 => "0000000000110001",
6195 => "0000000000110001",
6196 => "0000000000110001",
6197 => "0000000000110001",
6198 => "0000000000110001",
6199 => "0000000000110001",
6200 => "0000000000110001",
6201 => "0000000000110001",
6202 => "0000000000110001",
6203 => "0000000000110001",
6204 => "0000000000110001",
6205 => "0000000000110001",
6206 => "0000000000110001",
6207 => "0000000000110001",
6208 => "0000000000110001",
6209 => "0000000000110001",
6210 => "0000000000110010",
6211 => "0000000000110010",
6212 => "0000000000110010",
6213 => "0000000000110010",
6214 => "0000000000110010",
6215 => "0000000000110010",
6216 => "0000000000110010",
6217 => "0000000000110010",
6218 => "0000000000110010",
6219 => "0000000000110010",
6220 => "0000000000110010",
6221 => "0000000000110010",
6222 => "0000000000110010",
6223 => "0000000000110010",
6224 => "0000000000110010",
6225 => "0000000000110010",
6226 => "0000000000110010",
6227 => "0000000000110010",
6228 => "0000000000110010",
6229 => "0000000000110010",
6230 => "0000000000110010",
6231 => "0000000000110010",
6232 => "0000000000110010",
6233 => "0000000000110010",
6234 => "0000000000110010",
6235 => "0000000000110010",
6236 => "0000000000110010",
6237 => "0000000000110010",
6238 => "0000000000110010",
6239 => "0000000000110010",
6240 => "0000000000110010",
6241 => "0000000000110010",
6242 => "0000000000110010",
6243 => "0000000000110010",
6244 => "0000000000110010",
6245 => "0000000000110010",
6246 => "0000000000110010",
6247 => "0000000000110010",
6248 => "0000000000110010",
6249 => "0000000000110010",
6250 => "0000000000110010",
6251 => "0000000000110010",
6252 => "0000000000110010",
6253 => "0000000000110010",
6254 => "0000000000110010",
6255 => "0000000000110010",
6256 => "0000000000110010",
6257 => "0000000000110010",
6258 => "0000000000110010",
6259 => "0000000000110010",
6260 => "0000000000110010",
6261 => "0000000000110010",
6262 => "0000000000110010",
6263 => "0000000000110010",
6264 => "0000000000110010",
6265 => "0000000000110010",
6266 => "0000000000110010",
6267 => "0000000000110010",
6268 => "0000000000110010",
6269 => "0000000000110010",
6270 => "0000000000110010",
6271 => "0000000000110010",
6272 => "0000000000110010",
6273 => "0000000000110010",
6274 => "0000000000110010",
6275 => "0000000000110010",
6276 => "0000000000110010",
6277 => "0000000000110010",
6278 => "0000000000110010",
6279 => "0000000000110010",
6280 => "0000000000110010",
6281 => "0000000000110010",
6282 => "0000000000110010",
6283 => "0000000000110010",
6284 => "0000000000110010",
6285 => "0000000000110010",
6286 => "0000000000110010",
6287 => "0000000000110010",
6288 => "0000000000110010",
6289 => "0000000000110010",
6290 => "0000000000110010",
6291 => "0000000000110011",
6292 => "0000000000110011",
6293 => "0000000000110011",
6294 => "0000000000110011",
6295 => "0000000000110011",
6296 => "0000000000110011",
6297 => "0000000000110011",
6298 => "0000000000110011",
6299 => "0000000000110011",
6300 => "0000000000110011",
6301 => "0000000000110011",
6302 => "0000000000110011",
6303 => "0000000000110011",
6304 => "0000000000110011",
6305 => "0000000000110011",
6306 => "0000000000110011",
6307 => "0000000000110011",
6308 => "0000000000110011",
6309 => "0000000000110011",
6310 => "0000000000110011",
6311 => "0000000000110011",
6312 => "0000000000110011",
6313 => "0000000000110011",
6314 => "0000000000110011",
6315 => "0000000000110011",
6316 => "0000000000110011",
6317 => "0000000000110011",
6318 => "0000000000110011",
6319 => "0000000000110011",
6320 => "0000000000110011",
6321 => "0000000000110011",
6322 => "0000000000110011",
6323 => "0000000000110011",
6324 => "0000000000110011",
6325 => "0000000000110011",
6326 => "0000000000110011",
6327 => "0000000000110011",
6328 => "0000000000110011",
6329 => "0000000000110011",
6330 => "0000000000110011",
6331 => "0000000000110011",
6332 => "0000000000110011",
6333 => "0000000000110011",
6334 => "0000000000110011",
6335 => "0000000000110011",
6336 => "0000000000110011",
6337 => "0000000000110011",
6338 => "0000000000110011",
6339 => "0000000000110011",
6340 => "0000000000110011",
6341 => "0000000000110011",
6342 => "0000000000110011",
6343 => "0000000000110011",
6344 => "0000000000110011",
6345 => "0000000000110011",
6346 => "0000000000110011",
6347 => "0000000000110011",
6348 => "0000000000110011",
6349 => "0000000000110011",
6350 => "0000000000110011",
6351 => "0000000000110011",
6352 => "0000000000110011",
6353 => "0000000000110011",
6354 => "0000000000110011",
6355 => "0000000000110011",
6356 => "0000000000110011",
6357 => "0000000000110011",
6358 => "0000000000110011",
6359 => "0000000000110011",
6360 => "0000000000110011",
6361 => "0000000000110011",
6362 => "0000000000110011",
6363 => "0000000000110011",
6364 => "0000000000110011",
6365 => "0000000000110011",
6366 => "0000000000110011",
6367 => "0000000000110011",
6368 => "0000000000110011",
6369 => "0000000000110011",
6370 => "0000000000110011",
6371 => "0000000000110100",
6372 => "0000000000110100",
6373 => "0000000000110100",
6374 => "0000000000110100",
6375 => "0000000000110100",
6376 => "0000000000110100",
6377 => "0000000000110100",
6378 => "0000000000110100",
6379 => "0000000000110100",
6380 => "0000000000110100",
6381 => "0000000000110100",
6382 => "0000000000110100",
6383 => "0000000000110100",
6384 => "0000000000110100",
6385 => "0000000000110100",
6386 => "0000000000110100",
6387 => "0000000000110100",
6388 => "0000000000110100",
6389 => "0000000000110100",
6390 => "0000000000110100",
6391 => "0000000000110100",
6392 => "0000000000110100",
6393 => "0000000000110100",
6394 => "0000000000110100",
6395 => "0000000000110100",
6396 => "0000000000110100",
6397 => "0000000000110100",
6398 => "0000000000110100",
6399 => "0000000000110100",
6400 => "0000000000110100",
6401 => "0000000000110100",
6402 => "0000000000110100",
6403 => "0000000000110100",
6404 => "0000000000110100",
6405 => "0000000000110100",
6406 => "0000000000110100",
6407 => "0000000000110100",
6408 => "0000000000110100",
6409 => "0000000000110100",
6410 => "0000000000110100",
6411 => "0000000000110100",
6412 => "0000000000110100",
6413 => "0000000000110100",
6414 => "0000000000110100",
6415 => "0000000000110100",
6416 => "0000000000110100",
6417 => "0000000000110100",
6418 => "0000000000110100",
6419 => "0000000000110100",
6420 => "0000000000110100",
6421 => "0000000000110100",
6422 => "0000000000110100",
6423 => "0000000000110100",
6424 => "0000000000110100",
6425 => "0000000000110100",
6426 => "0000000000110100",
6427 => "0000000000110100",
6428 => "0000000000110100",
6429 => "0000000000110100",
6430 => "0000000000110100",
6431 => "0000000000110100",
6432 => "0000000000110100",
6433 => "0000000000110100",
6434 => "0000000000110100",
6435 => "0000000000110100",
6436 => "0000000000110100",
6437 => "0000000000110100",
6438 => "0000000000110100",
6439 => "0000000000110100",
6440 => "0000000000110100",
6441 => "0000000000110100",
6442 => "0000000000110100",
6443 => "0000000000110100",
6444 => "0000000000110100",
6445 => "0000000000110100",
6446 => "0000000000110100",
6447 => "0000000000110100",
6448 => "0000000000110100",
6449 => "0000000000110101",
6450 => "0000000000110101",
6451 => "0000000000110101",
6452 => "0000000000110101",
6453 => "0000000000110101",
6454 => "0000000000110101",
6455 => "0000000000110101",
6456 => "0000000000110101",
6457 => "0000000000110101",
6458 => "0000000000110101",
6459 => "0000000000110101",
6460 => "0000000000110101",
6461 => "0000000000110101",
6462 => "0000000000110101",
6463 => "0000000000110101",
6464 => "0000000000110101",
6465 => "0000000000110101",
6466 => "0000000000110101",
6467 => "0000000000110101",
6468 => "0000000000110101",
6469 => "0000000000110101",
6470 => "0000000000110101",
6471 => "0000000000110101",
6472 => "0000000000110101",
6473 => "0000000000110101",
6474 => "0000000000110101",
6475 => "0000000000110101",
6476 => "0000000000110101",
6477 => "0000000000110101",
6478 => "0000000000110101",
6479 => "0000000000110101",
6480 => "0000000000110101",
6481 => "0000000000110101",
6482 => "0000000000110101",
6483 => "0000000000110101",
6484 => "0000000000110101",
6485 => "0000000000110101",
6486 => "0000000000110101",
6487 => "0000000000110101",
6488 => "0000000000110101",
6489 => "0000000000110101",
6490 => "0000000000110101",
6491 => "0000000000110101",
6492 => "0000000000110101",
6493 => "0000000000110101",
6494 => "0000000000110101",
6495 => "0000000000110101",
6496 => "0000000000110101",
6497 => "0000000000110101",
6498 => "0000000000110101",
6499 => "0000000000110101",
6500 => "0000000000110101",
6501 => "0000000000110101",
6502 => "0000000000110101",
6503 => "0000000000110101",
6504 => "0000000000110101",
6505 => "0000000000110101",
6506 => "0000000000110101",
6507 => "0000000000110101",
6508 => "0000000000110101",
6509 => "0000000000110101",
6510 => "0000000000110101",
6511 => "0000000000110101",
6512 => "0000000000110101",
6513 => "0000000000110101",
6514 => "0000000000110101",
6515 => "0000000000110101",
6516 => "0000000000110101",
6517 => "0000000000110101",
6518 => "0000000000110101",
6519 => "0000000000110101",
6520 => "0000000000110101",
6521 => "0000000000110101",
6522 => "0000000000110101",
6523 => "0000000000110101",
6524 => "0000000000110101",
6525 => "0000000000110101",
6526 => "0000000000110110",
6527 => "0000000000110110",
6528 => "0000000000110110",
6529 => "0000000000110110",
6530 => "0000000000110110",
6531 => "0000000000110110",
6532 => "0000000000110110",
6533 => "0000000000110110",
6534 => "0000000000110110",
6535 => "0000000000110110",
6536 => "0000000000110110",
6537 => "0000000000110110",
6538 => "0000000000110110",
6539 => "0000000000110110",
6540 => "0000000000110110",
6541 => "0000000000110110",
6542 => "0000000000110110",
6543 => "0000000000110110",
6544 => "0000000000110110",
6545 => "0000000000110110",
6546 => "0000000000110110",
6547 => "0000000000110110",
6548 => "0000000000110110",
6549 => "0000000000110110",
6550 => "0000000000110110",
6551 => "0000000000110110",
6552 => "0000000000110110",
6553 => "0000000000110110",
6554 => "0000000000110110",
6555 => "0000000000110110",
6556 => "0000000000110110",
6557 => "0000000000110110",
6558 => "0000000000110110",
6559 => "0000000000110110",
6560 => "0000000000110110",
6561 => "0000000000110110",
6562 => "0000000000110110",
6563 => "0000000000110110",
6564 => "0000000000110110",
6565 => "0000000000110110",
6566 => "0000000000110110",
6567 => "0000000000110110",
6568 => "0000000000110110",
6569 => "0000000000110110",
6570 => "0000000000110110",
6571 => "0000000000110110",
6572 => "0000000000110110",
6573 => "0000000000110110",
6574 => "0000000000110110",
6575 => "0000000000110110",
6576 => "0000000000110110",
6577 => "0000000000110110",
6578 => "0000000000110110",
6579 => "0000000000110110",
6580 => "0000000000110110",
6581 => "0000000000110110",
6582 => "0000000000110110",
6583 => "0000000000110110",
6584 => "0000000000110110",
6585 => "0000000000110110",
6586 => "0000000000110110",
6587 => "0000000000110110",
6588 => "0000000000110110",
6589 => "0000000000110110",
6590 => "0000000000110110",
6591 => "0000000000110110",
6592 => "0000000000110110",
6593 => "0000000000110110",
6594 => "0000000000110110",
6595 => "0000000000110110",
6596 => "0000000000110110",
6597 => "0000000000110110",
6598 => "0000000000110110",
6599 => "0000000000110110",
6600 => "0000000000110110",
6601 => "0000000000110111",
6602 => "0000000000110111",
6603 => "0000000000110111",
6604 => "0000000000110111",
6605 => "0000000000110111",
6606 => "0000000000110111",
6607 => "0000000000110111",
6608 => "0000000000110111",
6609 => "0000000000110111",
6610 => "0000000000110111",
6611 => "0000000000110111",
6612 => "0000000000110111",
6613 => "0000000000110111",
6614 => "0000000000110111",
6615 => "0000000000110111",
6616 => "0000000000110111",
6617 => "0000000000110111",
6618 => "0000000000110111",
6619 => "0000000000110111",
6620 => "0000000000110111",
6621 => "0000000000110111",
6622 => "0000000000110111",
6623 => "0000000000110111",
6624 => "0000000000110111",
6625 => "0000000000110111",
6626 => "0000000000110111",
6627 => "0000000000110111",
6628 => "0000000000110111",
6629 => "0000000000110111",
6630 => "0000000000110111",
6631 => "0000000000110111",
6632 => "0000000000110111",
6633 => "0000000000110111",
6634 => "0000000000110111",
6635 => "0000000000110111",
6636 => "0000000000110111",
6637 => "0000000000110111",
6638 => "0000000000110111",
6639 => "0000000000110111",
6640 => "0000000000110111",
6641 => "0000000000110111",
6642 => "0000000000110111",
6643 => "0000000000110111",
6644 => "0000000000110111",
6645 => "0000000000110111",
6646 => "0000000000110111",
6647 => "0000000000110111",
6648 => "0000000000110111",
6649 => "0000000000110111",
6650 => "0000000000110111",
6651 => "0000000000110111",
6652 => "0000000000110111",
6653 => "0000000000110111",
6654 => "0000000000110111",
6655 => "0000000000110111",
6656 => "0000000000110111",
6657 => "0000000000110111",
6658 => "0000000000110111",
6659 => "0000000000110111",
6660 => "0000000000110111",
6661 => "0000000000110111",
6662 => "0000000000110111",
6663 => "0000000000110111",
6664 => "0000000000110111",
6665 => "0000000000110111",
6666 => "0000000000110111",
6667 => "0000000000110111",
6668 => "0000000000110111",
6669 => "0000000000110111",
6670 => "0000000000110111",
6671 => "0000000000110111",
6672 => "0000000000110111",
6673 => "0000000000110111",
6674 => "0000000000110111",
6675 => "0000000000111000",
6676 => "0000000000111000",
6677 => "0000000000111000",
6678 => "0000000000111000",
6679 => "0000000000111000",
6680 => "0000000000111000",
6681 => "0000000000111000",
6682 => "0000000000111000",
6683 => "0000000000111000",
6684 => "0000000000111000",
6685 => "0000000000111000",
6686 => "0000000000111000",
6687 => "0000000000111000",
6688 => "0000000000111000",
6689 => "0000000000111000",
6690 => "0000000000111000",
6691 => "0000000000111000",
6692 => "0000000000111000",
6693 => "0000000000111000",
6694 => "0000000000111000",
6695 => "0000000000111000",
6696 => "0000000000111000",
6697 => "0000000000111000",
6698 => "0000000000111000",
6699 => "0000000000111000",
6700 => "0000000000111000",
6701 => "0000000000111000",
6702 => "0000000000111000",
6703 => "0000000000111000",
6704 => "0000000000111000",
6705 => "0000000000111000",
6706 => "0000000000111000",
6707 => "0000000000111000",
6708 => "0000000000111000",
6709 => "0000000000111000",
6710 => "0000000000111000",
6711 => "0000000000111000",
6712 => "0000000000111000",
6713 => "0000000000111000",
6714 => "0000000000111000",
6715 => "0000000000111000",
6716 => "0000000000111000",
6717 => "0000000000111000",
6718 => "0000000000111000",
6719 => "0000000000111000",
6720 => "0000000000111000",
6721 => "0000000000111000",
6722 => "0000000000111000",
6723 => "0000000000111000",
6724 => "0000000000111000",
6725 => "0000000000111000",
6726 => "0000000000111000",
6727 => "0000000000111000",
6728 => "0000000000111000",
6729 => "0000000000111000",
6730 => "0000000000111000",
6731 => "0000000000111000",
6732 => "0000000000111000",
6733 => "0000000000111000",
6734 => "0000000000111000",
6735 => "0000000000111000",
6736 => "0000000000111000",
6737 => "0000000000111000",
6738 => "0000000000111000",
6739 => "0000000000111000",
6740 => "0000000000111000",
6741 => "0000000000111000",
6742 => "0000000000111000",
6743 => "0000000000111000",
6744 => "0000000000111000",
6745 => "0000000000111000",
6746 => "0000000000111000",
6747 => "0000000000111000",
6748 => "0000000000111001",
6749 => "0000000000111001",
6750 => "0000000000111001",
6751 => "0000000000111001",
6752 => "0000000000111001",
6753 => "0000000000111001",
6754 => "0000000000111001",
6755 => "0000000000111001",
6756 => "0000000000111001",
6757 => "0000000000111001",
6758 => "0000000000111001",
6759 => "0000000000111001",
6760 => "0000000000111001",
6761 => "0000000000111001",
6762 => "0000000000111001",
6763 => "0000000000111001",
6764 => "0000000000111001",
6765 => "0000000000111001",
6766 => "0000000000111001",
6767 => "0000000000111001",
6768 => "0000000000111001",
6769 => "0000000000111001",
6770 => "0000000000111001",
6771 => "0000000000111001",
6772 => "0000000000111001",
6773 => "0000000000111001",
6774 => "0000000000111001",
6775 => "0000000000111001",
6776 => "0000000000111001",
6777 => "0000000000111001",
6778 => "0000000000111001",
6779 => "0000000000111001",
6780 => "0000000000111001",
6781 => "0000000000111001",
6782 => "0000000000111001",
6783 => "0000000000111001",
6784 => "0000000000111001",
6785 => "0000000000111001",
6786 => "0000000000111001",
6787 => "0000000000111001",
6788 => "0000000000111001",
6789 => "0000000000111001",
6790 => "0000000000111001",
6791 => "0000000000111001",
6792 => "0000000000111001",
6793 => "0000000000111001",
6794 => "0000000000111001",
6795 => "0000000000111001",
6796 => "0000000000111001",
6797 => "0000000000111001",
6798 => "0000000000111001",
6799 => "0000000000111001",
6800 => "0000000000111001",
6801 => "0000000000111001",
6802 => "0000000000111001",
6803 => "0000000000111001",
6804 => "0000000000111001",
6805 => "0000000000111001",
6806 => "0000000000111001",
6807 => "0000000000111001",
6808 => "0000000000111001",
6809 => "0000000000111001",
6810 => "0000000000111001",
6811 => "0000000000111001",
6812 => "0000000000111001",
6813 => "0000000000111001",
6814 => "0000000000111001",
6815 => "0000000000111001",
6816 => "0000000000111001",
6817 => "0000000000111001",
6818 => "0000000000111001",
6819 => "0000000000111010",
6820 => "0000000000111010",
6821 => "0000000000111010",
6822 => "0000000000111010",
6823 => "0000000000111010",
6824 => "0000000000111010",
6825 => "0000000000111010",
6826 => "0000000000111010",
6827 => "0000000000111010",
6828 => "0000000000111010",
6829 => "0000000000111010",
6830 => "0000000000111010",
6831 => "0000000000111010",
6832 => "0000000000111010",
6833 => "0000000000111010",
6834 => "0000000000111010",
6835 => "0000000000111010",
6836 => "0000000000111010",
6837 => "0000000000111010",
6838 => "0000000000111010",
6839 => "0000000000111010",
6840 => "0000000000111010",
6841 => "0000000000111010",
6842 => "0000000000111010",
6843 => "0000000000111010",
6844 => "0000000000111010",
6845 => "0000000000111010",
6846 => "0000000000111010",
6847 => "0000000000111010",
6848 => "0000000000111010",
6849 => "0000000000111010",
6850 => "0000000000111010",
6851 => "0000000000111010",
6852 => "0000000000111010",
6853 => "0000000000111010",
6854 => "0000000000111010",
6855 => "0000000000111010",
6856 => "0000000000111010",
6857 => "0000000000111010",
6858 => "0000000000111010",
6859 => "0000000000111010",
6860 => "0000000000111010",
6861 => "0000000000111010",
6862 => "0000000000111010",
6863 => "0000000000111010",
6864 => "0000000000111010",
6865 => "0000000000111010",
6866 => "0000000000111010",
6867 => "0000000000111010",
6868 => "0000000000111010",
6869 => "0000000000111010",
6870 => "0000000000111010",
6871 => "0000000000111010",
6872 => "0000000000111010",
6873 => "0000000000111010",
6874 => "0000000000111010",
6875 => "0000000000111010",
6876 => "0000000000111010",
6877 => "0000000000111010",
6878 => "0000000000111010",
6879 => "0000000000111010",
6880 => "0000000000111010",
6881 => "0000000000111010",
6882 => "0000000000111010",
6883 => "0000000000111010",
6884 => "0000000000111010",
6885 => "0000000000111010",
6886 => "0000000000111010",
6887 => "0000000000111010",
6888 => "0000000000111010",
6889 => "0000000000111011",
6890 => "0000000000111011",
6891 => "0000000000111011",
6892 => "0000000000111011",
6893 => "0000000000111011",
6894 => "0000000000111011",
6895 => "0000000000111011",
6896 => "0000000000111011",
6897 => "0000000000111011",
6898 => "0000000000111011",
6899 => "0000000000111011",
6900 => "0000000000111011",
6901 => "0000000000111011",
6902 => "0000000000111011",
6903 => "0000000000111011",
6904 => "0000000000111011",
6905 => "0000000000111011",
6906 => "0000000000111011",
6907 => "0000000000111011",
6908 => "0000000000111011",
6909 => "0000000000111011",
6910 => "0000000000111011",
6911 => "0000000000111011",
6912 => "0000000000111011",
6913 => "0000000000111011",
6914 => "0000000000111011",
6915 => "0000000000111011",
6916 => "0000000000111011",
6917 => "0000000000111011",
6918 => "0000000000111011",
6919 => "0000000000111011",
6920 => "0000000000111011",
6921 => "0000000000111011",
6922 => "0000000000111011",
6923 => "0000000000111011",
6924 => "0000000000111011",
6925 => "0000000000111011",
6926 => "0000000000111011",
6927 => "0000000000111011",
6928 => "0000000000111011",
6929 => "0000000000111011",
6930 => "0000000000111011",
6931 => "0000000000111011",
6932 => "0000000000111011",
6933 => "0000000000111011",
6934 => "0000000000111011",
6935 => "0000000000111011",
6936 => "0000000000111011",
6937 => "0000000000111011",
6938 => "0000000000111011",
6939 => "0000000000111011",
6940 => "0000000000111011",
6941 => "0000000000111011",
6942 => "0000000000111011",
6943 => "0000000000111011",
6944 => "0000000000111011",
6945 => "0000000000111011",
6946 => "0000000000111011",
6947 => "0000000000111011",
6948 => "0000000000111011",
6949 => "0000000000111011",
6950 => "0000000000111011",
6951 => "0000000000111011",
6952 => "0000000000111011",
6953 => "0000000000111011",
6954 => "0000000000111011",
6955 => "0000000000111011",
6956 => "0000000000111011",
6957 => "0000000000111011",
6958 => "0000000000111100",
6959 => "0000000000111100",
6960 => "0000000000111100",
6961 => "0000000000111100",
6962 => "0000000000111100",
6963 => "0000000000111100",
6964 => "0000000000111100",
6965 => "0000000000111100",
6966 => "0000000000111100",
6967 => "0000000000111100",
6968 => "0000000000111100",
6969 => "0000000000111100",
6970 => "0000000000111100",
6971 => "0000000000111100",
6972 => "0000000000111100",
6973 => "0000000000111100",
6974 => "0000000000111100",
6975 => "0000000000111100",
6976 => "0000000000111100",
6977 => "0000000000111100",
6978 => "0000000000111100",
6979 => "0000000000111100",
6980 => "0000000000111100",
6981 => "0000000000111100",
6982 => "0000000000111100",
6983 => "0000000000111100",
6984 => "0000000000111100",
6985 => "0000000000111100",
6986 => "0000000000111100",
6987 => "0000000000111100",
6988 => "0000000000111100",
6989 => "0000000000111100",
6990 => "0000000000111100",
6991 => "0000000000111100",
6992 => "0000000000111100",
6993 => "0000000000111100",
6994 => "0000000000111100",
6995 => "0000000000111100",
6996 => "0000000000111100",
6997 => "0000000000111100",
6998 => "0000000000111100",
6999 => "0000000000111100",
7000 => "0000000000111100",
7001 => "0000000000111100",
7002 => "0000000000111100",
7003 => "0000000000111100",
7004 => "0000000000111100",
7005 => "0000000000111100",
7006 => "0000000000111100",
7007 => "0000000000111100",
7008 => "0000000000111100",
7009 => "0000000000111100",
7010 => "0000000000111100",
7011 => "0000000000111100",
7012 => "0000000000111100",
7013 => "0000000000111100",
7014 => "0000000000111100",
7015 => "0000000000111100",
7016 => "0000000000111100",
7017 => "0000000000111100",
7018 => "0000000000111100",
7019 => "0000000000111100",
7020 => "0000000000111100",
7021 => "0000000000111100",
7022 => "0000000000111100",
7023 => "0000000000111100",
7024 => "0000000000111100",
7025 => "0000000000111100",
7026 => "0000000000111101",
7027 => "0000000000111101",
7028 => "0000000000111101",
7029 => "0000000000111101",
7030 => "0000000000111101",
7031 => "0000000000111101",
7032 => "0000000000111101",
7033 => "0000000000111101",
7034 => "0000000000111101",
7035 => "0000000000111101",
7036 => "0000000000111101",
7037 => "0000000000111101",
7038 => "0000000000111101",
7039 => "0000000000111101",
7040 => "0000000000111101",
7041 => "0000000000111101",
7042 => "0000000000111101",
7043 => "0000000000111101",
7044 => "0000000000111101",
7045 => "0000000000111101",
7046 => "0000000000111101",
7047 => "0000000000111101",
7048 => "0000000000111101",
7049 => "0000000000111101",
7050 => "0000000000111101",
7051 => "0000000000111101",
7052 => "0000000000111101",
7053 => "0000000000111101",
7054 => "0000000000111101",
7055 => "0000000000111101",
7056 => "0000000000111101",
7057 => "0000000000111101",
7058 => "0000000000111101",
7059 => "0000000000111101",
7060 => "0000000000111101",
7061 => "0000000000111101",
7062 => "0000000000111101",
7063 => "0000000000111101",
7064 => "0000000000111101",
7065 => "0000000000111101",
7066 => "0000000000111101",
7067 => "0000000000111101",
7068 => "0000000000111101",
7069 => "0000000000111101",
7070 => "0000000000111101",
7071 => "0000000000111101",
7072 => "0000000000111101",
7073 => "0000000000111101",
7074 => "0000000000111101",
7075 => "0000000000111101",
7076 => "0000000000111101",
7077 => "0000000000111101",
7078 => "0000000000111101",
7079 => "0000000000111101",
7080 => "0000000000111101",
7081 => "0000000000111101",
7082 => "0000000000111101",
7083 => "0000000000111101",
7084 => "0000000000111101",
7085 => "0000000000111101",
7086 => "0000000000111101",
7087 => "0000000000111101",
7088 => "0000000000111101",
7089 => "0000000000111101",
7090 => "0000000000111101",
7091 => "0000000000111101",
7092 => "0000000000111101",
7093 => "0000000000111110",
7094 => "0000000000111110",
7095 => "0000000000111110",
7096 => "0000000000111110",
7097 => "0000000000111110",
7098 => "0000000000111110",
7099 => "0000000000111110",
7100 => "0000000000111110",
7101 => "0000000000111110",
7102 => "0000000000111110",
7103 => "0000000000111110",
7104 => "0000000000111110",
7105 => "0000000000111110",
7106 => "0000000000111110",
7107 => "0000000000111110",
7108 => "0000000000111110",
7109 => "0000000000111110",
7110 => "0000000000111110",
7111 => "0000000000111110",
7112 => "0000000000111110",
7113 => "0000000000111110",
7114 => "0000000000111110",
7115 => "0000000000111110",
7116 => "0000000000111110",
7117 => "0000000000111110",
7118 => "0000000000111110",
7119 => "0000000000111110",
7120 => "0000000000111110",
7121 => "0000000000111110",
7122 => "0000000000111110",
7123 => "0000000000111110",
7124 => "0000000000111110",
7125 => "0000000000111110",
7126 => "0000000000111110",
7127 => "0000000000111110",
7128 => "0000000000111110",
7129 => "0000000000111110",
7130 => "0000000000111110",
7131 => "0000000000111110",
7132 => "0000000000111110",
7133 => "0000000000111110",
7134 => "0000000000111110",
7135 => "0000000000111110",
7136 => "0000000000111110",
7137 => "0000000000111110",
7138 => "0000000000111110",
7139 => "0000000000111110",
7140 => "0000000000111110",
7141 => "0000000000111110",
7142 => "0000000000111110",
7143 => "0000000000111110",
7144 => "0000000000111110",
7145 => "0000000000111110",
7146 => "0000000000111110",
7147 => "0000000000111110",
7148 => "0000000000111110",
7149 => "0000000000111110",
7150 => "0000000000111110",
7151 => "0000000000111110",
7152 => "0000000000111110",
7153 => "0000000000111110",
7154 => "0000000000111110",
7155 => "0000000000111110",
7156 => "0000000000111110",
7157 => "0000000000111110",
7158 => "0000000000111110",
7159 => "0000000000111111",
7160 => "0000000000111111",
7161 => "0000000000111111",
7162 => "0000000000111111",
7163 => "0000000000111111",
7164 => "0000000000111111",
7165 => "0000000000111111",
7166 => "0000000000111111",
7167 => "0000000000111111",
7168 => "0000000000111111",
7169 => "0000000000111111",
7170 => "0000000000111111",
7171 => "0000000000111111",
7172 => "0000000000111111",
7173 => "0000000000111111",
7174 => "0000000000111111",
7175 => "0000000000111111",
7176 => "0000000000111111",
7177 => "0000000000111111",
7178 => "0000000000111111",
7179 => "0000000000111111",
7180 => "0000000000111111",
7181 => "0000000000111111",
7182 => "0000000000111111",
7183 => "0000000000111111",
7184 => "0000000000111111",
7185 => "0000000000111111",
7186 => "0000000000111111",
7187 => "0000000000111111",
7188 => "0000000000111111",
7189 => "0000000000111111",
7190 => "0000000000111111",
7191 => "0000000000111111",
7192 => "0000000000111111",
7193 => "0000000000111111",
7194 => "0000000000111111",
7195 => "0000000000111111",
7196 => "0000000000111111",
7197 => "0000000000111111",
7198 => "0000000000111111",
7199 => "0000000000111111",
7200 => "0000000000111111",
7201 => "0000000000111111",
7202 => "0000000000111111",
7203 => "0000000000111111",
7204 => "0000000000111111",
7205 => "0000000000111111",
7206 => "0000000000111111",
7207 => "0000000000111111",
7208 => "0000000000111111",
7209 => "0000000000111111",
7210 => "0000000000111111",
7211 => "0000000000111111",
7212 => "0000000000111111",
7213 => "0000000000111111",
7214 => "0000000000111111",
7215 => "0000000000111111",
7216 => "0000000000111111",
7217 => "0000000000111111",
7218 => "0000000000111111",
7219 => "0000000000111111",
7220 => "0000000000111111",
7221 => "0000000000111111",
7222 => "0000000000111111",
7223 => "0000000001000000",
7224 => "0000000001000000",
7225 => "0000000001000000",
7226 => "0000000001000000",
7227 => "0000000001000000",
7228 => "0000000001000000",
7229 => "0000000001000000",
7230 => "0000000001000000",
7231 => "0000000001000000",
7232 => "0000000001000000",
7233 => "0000000001000000",
7234 => "0000000001000000",
7235 => "0000000001000000",
7236 => "0000000001000000",
7237 => "0000000001000000",
7238 => "0000000001000000",
7239 => "0000000001000000",
7240 => "0000000001000000",
7241 => "0000000001000000",
7242 => "0000000001000000",
7243 => "0000000001000000",
7244 => "0000000001000000",
7245 => "0000000001000000",
7246 => "0000000001000000",
7247 => "0000000001000000",
7248 => "0000000001000000",
7249 => "0000000001000000",
7250 => "0000000001000000",
7251 => "0000000001000000",
7252 => "0000000001000000",
7253 => "0000000001000000",
7254 => "0000000001000000",
7255 => "0000000001000000",
7256 => "0000000001000000",
7257 => "0000000001000000",
7258 => "0000000001000000",
7259 => "0000000001000000",
7260 => "0000000001000000",
7261 => "0000000001000000",
7262 => "0000000001000000",
7263 => "0000000001000000",
7264 => "0000000001000000",
7265 => "0000000001000000",
7266 => "0000000001000000",
7267 => "0000000001000000",
7268 => "0000000001000000",
7269 => "0000000001000000",
7270 => "0000000001000000",
7271 => "0000000001000000",
7272 => "0000000001000000",
7273 => "0000000001000000",
7274 => "0000000001000000",
7275 => "0000000001000000",
7276 => "0000000001000000",
7277 => "0000000001000000",
7278 => "0000000001000000",
7279 => "0000000001000000",
7280 => "0000000001000000",
7281 => "0000000001000000",
7282 => "0000000001000000",
7283 => "0000000001000000",
7284 => "0000000001000000",
7285 => "0000000001000000",
7286 => "0000000001000001",
7287 => "0000000001000001",
7288 => "0000000001000001",
7289 => "0000000001000001",
7290 => "0000000001000001",
7291 => "0000000001000001",
7292 => "0000000001000001",
7293 => "0000000001000001",
7294 => "0000000001000001",
7295 => "0000000001000001",
7296 => "0000000001000001",
7297 => "0000000001000001",
7298 => "0000000001000001",
7299 => "0000000001000001",
7300 => "0000000001000001",
7301 => "0000000001000001",
7302 => "0000000001000001",
7303 => "0000000001000001",
7304 => "0000000001000001",
7305 => "0000000001000001",
7306 => "0000000001000001",
7307 => "0000000001000001",
7308 => "0000000001000001",
7309 => "0000000001000001",
7310 => "0000000001000001",
7311 => "0000000001000001",
7312 => "0000000001000001",
7313 => "0000000001000001",
7314 => "0000000001000001",
7315 => "0000000001000001",
7316 => "0000000001000001",
7317 => "0000000001000001",
7318 => "0000000001000001",
7319 => "0000000001000001",
7320 => "0000000001000001",
7321 => "0000000001000001",
7322 => "0000000001000001",
7323 => "0000000001000001",
7324 => "0000000001000001",
7325 => "0000000001000001",
7326 => "0000000001000001",
7327 => "0000000001000001",
7328 => "0000000001000001",
7329 => "0000000001000001",
7330 => "0000000001000001",
7331 => "0000000001000001",
7332 => "0000000001000001",
7333 => "0000000001000001",
7334 => "0000000001000001",
7335 => "0000000001000001",
7336 => "0000000001000001",
7337 => "0000000001000001",
7338 => "0000000001000001",
7339 => "0000000001000001",
7340 => "0000000001000001",
7341 => "0000000001000001",
7342 => "0000000001000001",
7343 => "0000000001000001",
7344 => "0000000001000001",
7345 => "0000000001000001",
7346 => "0000000001000001",
7347 => "0000000001000001",
7348 => "0000000001000001",
7349 => "0000000001000010",
7350 => "0000000001000010",
7351 => "0000000001000010",
7352 => "0000000001000010",
7353 => "0000000001000010",
7354 => "0000000001000010",
7355 => "0000000001000010",
7356 => "0000000001000010",
7357 => "0000000001000010",
7358 => "0000000001000010",
7359 => "0000000001000010",
7360 => "0000000001000010",
7361 => "0000000001000010",
7362 => "0000000001000010",
7363 => "0000000001000010",
7364 => "0000000001000010",
7365 => "0000000001000010",
7366 => "0000000001000010",
7367 => "0000000001000010",
7368 => "0000000001000010",
7369 => "0000000001000010",
7370 => "0000000001000010",
7371 => "0000000001000010",
7372 => "0000000001000010",
7373 => "0000000001000010",
7374 => "0000000001000010",
7375 => "0000000001000010",
7376 => "0000000001000010",
7377 => "0000000001000010",
7378 => "0000000001000010",
7379 => "0000000001000010",
7380 => "0000000001000010",
7381 => "0000000001000010",
7382 => "0000000001000010",
7383 => "0000000001000010",
7384 => "0000000001000010",
7385 => "0000000001000010",
7386 => "0000000001000010",
7387 => "0000000001000010",
7388 => "0000000001000010",
7389 => "0000000001000010",
7390 => "0000000001000010",
7391 => "0000000001000010",
7392 => "0000000001000010",
7393 => "0000000001000010",
7394 => "0000000001000010",
7395 => "0000000001000010",
7396 => "0000000001000010",
7397 => "0000000001000010",
7398 => "0000000001000010",
7399 => "0000000001000010",
7400 => "0000000001000010",
7401 => "0000000001000010",
7402 => "0000000001000010",
7403 => "0000000001000010",
7404 => "0000000001000010",
7405 => "0000000001000010",
7406 => "0000000001000010",
7407 => "0000000001000010",
7408 => "0000000001000010",
7409 => "0000000001000010",
7410 => "0000000001000011",
7411 => "0000000001000011",
7412 => "0000000001000011",
7413 => "0000000001000011",
7414 => "0000000001000011",
7415 => "0000000001000011",
7416 => "0000000001000011",
7417 => "0000000001000011",
7418 => "0000000001000011",
7419 => "0000000001000011",
7420 => "0000000001000011",
7421 => "0000000001000011",
7422 => "0000000001000011",
7423 => "0000000001000011",
7424 => "0000000001000011",
7425 => "0000000001000011",
7426 => "0000000001000011",
7427 => "0000000001000011",
7428 => "0000000001000011",
7429 => "0000000001000011",
7430 => "0000000001000011",
7431 => "0000000001000011",
7432 => "0000000001000011",
7433 => "0000000001000011",
7434 => "0000000001000011",
7435 => "0000000001000011",
7436 => "0000000001000011",
7437 => "0000000001000011",
7438 => "0000000001000011",
7439 => "0000000001000011",
7440 => "0000000001000011",
7441 => "0000000001000011",
7442 => "0000000001000011",
7443 => "0000000001000011",
7444 => "0000000001000011",
7445 => "0000000001000011",
7446 => "0000000001000011",
7447 => "0000000001000011",
7448 => "0000000001000011",
7449 => "0000000001000011",
7450 => "0000000001000011",
7451 => "0000000001000011",
7452 => "0000000001000011",
7453 => "0000000001000011",
7454 => "0000000001000011",
7455 => "0000000001000011",
7456 => "0000000001000011",
7457 => "0000000001000011",
7458 => "0000000001000011",
7459 => "0000000001000011",
7460 => "0000000001000011",
7461 => "0000000001000011",
7462 => "0000000001000011",
7463 => "0000000001000011",
7464 => "0000000001000011",
7465 => "0000000001000011",
7466 => "0000000001000011",
7467 => "0000000001000011",
7468 => "0000000001000011",
7469 => "0000000001000011",
7470 => "0000000001000011",
7471 => "0000000001000100",
7472 => "0000000001000100",
7473 => "0000000001000100",
7474 => "0000000001000100",
7475 => "0000000001000100",
7476 => "0000000001000100",
7477 => "0000000001000100",
7478 => "0000000001000100",
7479 => "0000000001000100",
7480 => "0000000001000100",
7481 => "0000000001000100",
7482 => "0000000001000100",
7483 => "0000000001000100",
7484 => "0000000001000100",
7485 => "0000000001000100",
7486 => "0000000001000100",
7487 => "0000000001000100",
7488 => "0000000001000100",
7489 => "0000000001000100",
7490 => "0000000001000100",
7491 => "0000000001000100",
7492 => "0000000001000100",
7493 => "0000000001000100",
7494 => "0000000001000100",
7495 => "0000000001000100",
7496 => "0000000001000100",
7497 => "0000000001000100",
7498 => "0000000001000100",
7499 => "0000000001000100",
7500 => "0000000001000100",
7501 => "0000000001000100",
7502 => "0000000001000100",
7503 => "0000000001000100",
7504 => "0000000001000100",
7505 => "0000000001000100",
7506 => "0000000001000100",
7507 => "0000000001000100",
7508 => "0000000001000100",
7509 => "0000000001000100",
7510 => "0000000001000100",
7511 => "0000000001000100",
7512 => "0000000001000100",
7513 => "0000000001000100",
7514 => "0000000001000100",
7515 => "0000000001000100",
7516 => "0000000001000100",
7517 => "0000000001000100",
7518 => "0000000001000100",
7519 => "0000000001000100",
7520 => "0000000001000100",
7521 => "0000000001000100",
7522 => "0000000001000100",
7523 => "0000000001000100",
7524 => "0000000001000100",
7525 => "0000000001000100",
7526 => "0000000001000100",
7527 => "0000000001000100",
7528 => "0000000001000100",
7529 => "0000000001000100",
7530 => "0000000001000100",
7531 => "0000000001000101",
7532 => "0000000001000101",
7533 => "0000000001000101",
7534 => "0000000001000101",
7535 => "0000000001000101",
7536 => "0000000001000101",
7537 => "0000000001000101",
7538 => "0000000001000101",
7539 => "0000000001000101",
7540 => "0000000001000101",
7541 => "0000000001000101",
7542 => "0000000001000101",
7543 => "0000000001000101",
7544 => "0000000001000101",
7545 => "0000000001000101",
7546 => "0000000001000101",
7547 => "0000000001000101",
7548 => "0000000001000101",
7549 => "0000000001000101",
7550 => "0000000001000101",
7551 => "0000000001000101",
7552 => "0000000001000101",
7553 => "0000000001000101",
7554 => "0000000001000101",
7555 => "0000000001000101",
7556 => "0000000001000101",
7557 => "0000000001000101",
7558 => "0000000001000101",
7559 => "0000000001000101",
7560 => "0000000001000101",
7561 => "0000000001000101",
7562 => "0000000001000101",
7563 => "0000000001000101",
7564 => "0000000001000101",
7565 => "0000000001000101",
7566 => "0000000001000101",
7567 => "0000000001000101",
7568 => "0000000001000101",
7569 => "0000000001000101",
7570 => "0000000001000101",
7571 => "0000000001000101",
7572 => "0000000001000101",
7573 => "0000000001000101",
7574 => "0000000001000101",
7575 => "0000000001000101",
7576 => "0000000001000101",
7577 => "0000000001000101",
7578 => "0000000001000101",
7579 => "0000000001000101",
7580 => "0000000001000101",
7581 => "0000000001000101",
7582 => "0000000001000101",
7583 => "0000000001000101",
7584 => "0000000001000101",
7585 => "0000000001000101",
7586 => "0000000001000101",
7587 => "0000000001000101",
7588 => "0000000001000101",
7589 => "0000000001000101",
7590 => "0000000001000110",
7591 => "0000000001000110",
7592 => "0000000001000110",
7593 => "0000000001000110",
7594 => "0000000001000110",
7595 => "0000000001000110",
7596 => "0000000001000110",
7597 => "0000000001000110",
7598 => "0000000001000110",
7599 => "0000000001000110",
7600 => "0000000001000110",
7601 => "0000000001000110",
7602 => "0000000001000110",
7603 => "0000000001000110",
7604 => "0000000001000110",
7605 => "0000000001000110",
7606 => "0000000001000110",
7607 => "0000000001000110",
7608 => "0000000001000110",
7609 => "0000000001000110",
7610 => "0000000001000110",
7611 => "0000000001000110",
7612 => "0000000001000110",
7613 => "0000000001000110",
7614 => "0000000001000110",
7615 => "0000000001000110",
7616 => "0000000001000110",
7617 => "0000000001000110",
7618 => "0000000001000110",
7619 => "0000000001000110",
7620 => "0000000001000110",
7621 => "0000000001000110",
7622 => "0000000001000110",
7623 => "0000000001000110",
7624 => "0000000001000110",
7625 => "0000000001000110",
7626 => "0000000001000110",
7627 => "0000000001000110",
7628 => "0000000001000110",
7629 => "0000000001000110",
7630 => "0000000001000110",
7631 => "0000000001000110",
7632 => "0000000001000110",
7633 => "0000000001000110",
7634 => "0000000001000110",
7635 => "0000000001000110",
7636 => "0000000001000110",
7637 => "0000000001000110",
7638 => "0000000001000110",
7639 => "0000000001000110",
7640 => "0000000001000110",
7641 => "0000000001000110",
7642 => "0000000001000110",
7643 => "0000000001000110",
7644 => "0000000001000110",
7645 => "0000000001000110",
7646 => "0000000001000110",
7647 => "0000000001000110",
7648 => "0000000001000111",
7649 => "0000000001000111",
7650 => "0000000001000111",
7651 => "0000000001000111",
7652 => "0000000001000111",
7653 => "0000000001000111",
7654 => "0000000001000111",
7655 => "0000000001000111",
7656 => "0000000001000111",
7657 => "0000000001000111",
7658 => "0000000001000111",
7659 => "0000000001000111",
7660 => "0000000001000111",
7661 => "0000000001000111",
7662 => "0000000001000111",
7663 => "0000000001000111",
7664 => "0000000001000111",
7665 => "0000000001000111",
7666 => "0000000001000111",
7667 => "0000000001000111",
7668 => "0000000001000111",
7669 => "0000000001000111",
7670 => "0000000001000111",
7671 => "0000000001000111",
7672 => "0000000001000111",
7673 => "0000000001000111",
7674 => "0000000001000111",
7675 => "0000000001000111",
7676 => "0000000001000111",
7677 => "0000000001000111",
7678 => "0000000001000111",
7679 => "0000000001000111",
7680 => "0000000001000111",
7681 => "0000000001000111",
7682 => "0000000001000111",
7683 => "0000000001000111",
7684 => "0000000001000111",
7685 => "0000000001000111",
7686 => "0000000001000111",
7687 => "0000000001000111",
7688 => "0000000001000111",
7689 => "0000000001000111",
7690 => "0000000001000111",
7691 => "0000000001000111",
7692 => "0000000001000111",
7693 => "0000000001000111",
7694 => "0000000001000111",
7695 => "0000000001000111",
7696 => "0000000001000111",
7697 => "0000000001000111",
7698 => "0000000001000111",
7699 => "0000000001000111",
7700 => "0000000001000111",
7701 => "0000000001000111",
7702 => "0000000001000111",
7703 => "0000000001000111",
7704 => "0000000001000111",
7705 => "0000000001000111",
7706 => "0000000001001000",
7707 => "0000000001001000",
7708 => "0000000001001000",
7709 => "0000000001001000",
7710 => "0000000001001000",
7711 => "0000000001001000",
7712 => "0000000001001000",
7713 => "0000000001001000",
7714 => "0000000001001000",
7715 => "0000000001001000",
7716 => "0000000001001000",
7717 => "0000000001001000",
7718 => "0000000001001000",
7719 => "0000000001001000",
7720 => "0000000001001000",
7721 => "0000000001001000",
7722 => "0000000001001000",
7723 => "0000000001001000",
7724 => "0000000001001000",
7725 => "0000000001001000",
7726 => "0000000001001000",
7727 => "0000000001001000",
7728 => "0000000001001000",
7729 => "0000000001001000",
7730 => "0000000001001000",
7731 => "0000000001001000",
7732 => "0000000001001000",
7733 => "0000000001001000",
7734 => "0000000001001000",
7735 => "0000000001001000",
7736 => "0000000001001000",
7737 => "0000000001001000",
7738 => "0000000001001000",
7739 => "0000000001001000",
7740 => "0000000001001000",
7741 => "0000000001001000",
7742 => "0000000001001000",
7743 => "0000000001001000",
7744 => "0000000001001000",
7745 => "0000000001001000",
7746 => "0000000001001000",
7747 => "0000000001001000",
7748 => "0000000001001000",
7749 => "0000000001001000",
7750 => "0000000001001000",
7751 => "0000000001001000",
7752 => "0000000001001000",
7753 => "0000000001001000",
7754 => "0000000001001000",
7755 => "0000000001001000",
7756 => "0000000001001000",
7757 => "0000000001001000",
7758 => "0000000001001000",
7759 => "0000000001001000",
7760 => "0000000001001000",
7761 => "0000000001001000",
7762 => "0000000001001000",
7763 => "0000000001001001",
7764 => "0000000001001001",
7765 => "0000000001001001",
7766 => "0000000001001001",
7767 => "0000000001001001",
7768 => "0000000001001001",
7769 => "0000000001001001",
7770 => "0000000001001001",
7771 => "0000000001001001",
7772 => "0000000001001001",
7773 => "0000000001001001",
7774 => "0000000001001001",
7775 => "0000000001001001",
7776 => "0000000001001001",
7777 => "0000000001001001",
7778 => "0000000001001001",
7779 => "0000000001001001",
7780 => "0000000001001001",
7781 => "0000000001001001",
7782 => "0000000001001001",
7783 => "0000000001001001",
7784 => "0000000001001001",
7785 => "0000000001001001",
7786 => "0000000001001001",
7787 => "0000000001001001",
7788 => "0000000001001001",
7789 => "0000000001001001",
7790 => "0000000001001001",
7791 => "0000000001001001",
7792 => "0000000001001001",
7793 => "0000000001001001",
7794 => "0000000001001001",
7795 => "0000000001001001",
7796 => "0000000001001001",
7797 => "0000000001001001",
7798 => "0000000001001001",
7799 => "0000000001001001",
7800 => "0000000001001001",
7801 => "0000000001001001",
7802 => "0000000001001001",
7803 => "0000000001001001",
7804 => "0000000001001001",
7805 => "0000000001001001",
7806 => "0000000001001001",
7807 => "0000000001001001",
7808 => "0000000001001001",
7809 => "0000000001001001",
7810 => "0000000001001001",
7811 => "0000000001001001",
7812 => "0000000001001001",
7813 => "0000000001001001",
7814 => "0000000001001001",
7815 => "0000000001001001",
7816 => "0000000001001001",
7817 => "0000000001001001",
7818 => "0000000001001010",
7819 => "0000000001001010",
7820 => "0000000001001010",
7821 => "0000000001001010",
7822 => "0000000001001010",
7823 => "0000000001001010",
7824 => "0000000001001010",
7825 => "0000000001001010",
7826 => "0000000001001010",
7827 => "0000000001001010",
7828 => "0000000001001010",
7829 => "0000000001001010",
7830 => "0000000001001010",
7831 => "0000000001001010",
7832 => "0000000001001010",
7833 => "0000000001001010",
7834 => "0000000001001010",
7835 => "0000000001001010",
7836 => "0000000001001010",
7837 => "0000000001001010",
7838 => "0000000001001010",
7839 => "0000000001001010",
7840 => "0000000001001010",
7841 => "0000000001001010",
7842 => "0000000001001010",
7843 => "0000000001001010",
7844 => "0000000001001010",
7845 => "0000000001001010",
7846 => "0000000001001010",
7847 => "0000000001001010",
7848 => "0000000001001010",
7849 => "0000000001001010",
7850 => "0000000001001010",
7851 => "0000000001001010",
7852 => "0000000001001010",
7853 => "0000000001001010",
7854 => "0000000001001010",
7855 => "0000000001001010",
7856 => "0000000001001010",
7857 => "0000000001001010",
7858 => "0000000001001010",
7859 => "0000000001001010",
7860 => "0000000001001010",
7861 => "0000000001001010",
7862 => "0000000001001010",
7863 => "0000000001001010",
7864 => "0000000001001010",
7865 => "0000000001001010",
7866 => "0000000001001010",
7867 => "0000000001001010",
7868 => "0000000001001010",
7869 => "0000000001001010",
7870 => "0000000001001010",
7871 => "0000000001001010",
7872 => "0000000001001010",
7873 => "0000000001001010",
7874 => "0000000001001011",
7875 => "0000000001001011",
7876 => "0000000001001011",
7877 => "0000000001001011",
7878 => "0000000001001011",
7879 => "0000000001001011",
7880 => "0000000001001011",
7881 => "0000000001001011",
7882 => "0000000001001011",
7883 => "0000000001001011",
7884 => "0000000001001011",
7885 => "0000000001001011",
7886 => "0000000001001011",
7887 => "0000000001001011",
7888 => "0000000001001011",
7889 => "0000000001001011",
7890 => "0000000001001011",
7891 => "0000000001001011",
7892 => "0000000001001011",
7893 => "0000000001001011",
7894 => "0000000001001011",
7895 => "0000000001001011",
7896 => "0000000001001011",
7897 => "0000000001001011",
7898 => "0000000001001011",
7899 => "0000000001001011",
7900 => "0000000001001011",
7901 => "0000000001001011",
7902 => "0000000001001011",
7903 => "0000000001001011",
7904 => "0000000001001011",
7905 => "0000000001001011",
7906 => "0000000001001011",
7907 => "0000000001001011",
7908 => "0000000001001011",
7909 => "0000000001001011",
7910 => "0000000001001011",
7911 => "0000000001001011",
7912 => "0000000001001011",
7913 => "0000000001001011",
7914 => "0000000001001011",
7915 => "0000000001001011",
7916 => "0000000001001011",
7917 => "0000000001001011",
7918 => "0000000001001011",
7919 => "0000000001001011",
7920 => "0000000001001011",
7921 => "0000000001001011",
7922 => "0000000001001011",
7923 => "0000000001001011",
7924 => "0000000001001011",
7925 => "0000000001001011",
7926 => "0000000001001011",
7927 => "0000000001001011",
7928 => "0000000001001100",
7929 => "0000000001001100",
7930 => "0000000001001100",
7931 => "0000000001001100",
7932 => "0000000001001100",
7933 => "0000000001001100",
7934 => "0000000001001100",
7935 => "0000000001001100",
7936 => "0000000001001100",
7937 => "0000000001001100",
7938 => "0000000001001100",
7939 => "0000000001001100",
7940 => "0000000001001100",
7941 => "0000000001001100",
7942 => "0000000001001100",
7943 => "0000000001001100",
7944 => "0000000001001100",
7945 => "0000000001001100",
7946 => "0000000001001100",
7947 => "0000000001001100",
7948 => "0000000001001100",
7949 => "0000000001001100",
7950 => "0000000001001100",
7951 => "0000000001001100",
7952 => "0000000001001100",
7953 => "0000000001001100",
7954 => "0000000001001100",
7955 => "0000000001001100",
7956 => "0000000001001100",
7957 => "0000000001001100",
7958 => "0000000001001100",
7959 => "0000000001001100",
7960 => "0000000001001100",
7961 => "0000000001001100",
7962 => "0000000001001100",
7963 => "0000000001001100",
7964 => "0000000001001100",
7965 => "0000000001001100",
7966 => "0000000001001100",
7967 => "0000000001001100",
7968 => "0000000001001100",
7969 => "0000000001001100",
7970 => "0000000001001100",
7971 => "0000000001001100",
7972 => "0000000001001100",
7973 => "0000000001001100",
7974 => "0000000001001100",
7975 => "0000000001001100",
7976 => "0000000001001100",
7977 => "0000000001001100",
7978 => "0000000001001100",
7979 => "0000000001001100",
7980 => "0000000001001100",
7981 => "0000000001001100",
7982 => "0000000001001101",
7983 => "0000000001001101",
7984 => "0000000001001101",
7985 => "0000000001001101",
7986 => "0000000001001101",
7987 => "0000000001001101",
7988 => "0000000001001101",
7989 => "0000000001001101",
7990 => "0000000001001101",
7991 => "0000000001001101",
7992 => "0000000001001101",
7993 => "0000000001001101",
7994 => "0000000001001101",
7995 => "0000000001001101",
7996 => "0000000001001101",
7997 => "0000000001001101",
7998 => "0000000001001101",
7999 => "0000000001001101",
8000 => "0000000001001101",
8001 => "0000000001001101",
8002 => "0000000001001101",
8003 => "0000000001001101",
8004 => "0000000001001101",
8005 => "0000000001001101",
8006 => "0000000001001101",
8007 => "0000000001001101",
8008 => "0000000001001101",
8009 => "0000000001001101",
8010 => "0000000001001101",
8011 => "0000000001001101",
8012 => "0000000001001101",
8013 => "0000000001001101",
8014 => "0000000001001101",
8015 => "0000000001001101",
8016 => "0000000001001101",
8017 => "0000000001001101",
8018 => "0000000001001101",
8019 => "0000000001001101",
8020 => "0000000001001101",
8021 => "0000000001001101",
8022 => "0000000001001101",
8023 => "0000000001001101",
8024 => "0000000001001101",
8025 => "0000000001001101",
8026 => "0000000001001101",
8027 => "0000000001001101",
8028 => "0000000001001101",
8029 => "0000000001001101",
8030 => "0000000001001101",
8031 => "0000000001001101",
8032 => "0000000001001101",
8033 => "0000000001001101",
8034 => "0000000001001101",
8035 => "0000000001001110",
8036 => "0000000001001110",
8037 => "0000000001001110",
8038 => "0000000001001110",
8039 => "0000000001001110",
8040 => "0000000001001110",
8041 => "0000000001001110",
8042 => "0000000001001110",
8043 => "0000000001001110",
8044 => "0000000001001110",
8045 => "0000000001001110",
8046 => "0000000001001110",
8047 => "0000000001001110",
8048 => "0000000001001110",
8049 => "0000000001001110",
8050 => "0000000001001110",
8051 => "0000000001001110",
8052 => "0000000001001110",
8053 => "0000000001001110",
8054 => "0000000001001110",
8055 => "0000000001001110",
8056 => "0000000001001110",
8057 => "0000000001001110",
8058 => "0000000001001110",
8059 => "0000000001001110",
8060 => "0000000001001110",
8061 => "0000000001001110",
8062 => "0000000001001110",
8063 => "0000000001001110",
8064 => "0000000001001110",
8065 => "0000000001001110",
8066 => "0000000001001110",
8067 => "0000000001001110",
8068 => "0000000001001110",
8069 => "0000000001001110",
8070 => "0000000001001110",
8071 => "0000000001001110",
8072 => "0000000001001110",
8073 => "0000000001001110",
8074 => "0000000001001110",
8075 => "0000000001001110",
8076 => "0000000001001110",
8077 => "0000000001001110",
8078 => "0000000001001110",
8079 => "0000000001001110",
8080 => "0000000001001110",
8081 => "0000000001001110",
8082 => "0000000001001110",
8083 => "0000000001001110",
8084 => "0000000001001110",
8085 => "0000000001001110",
8086 => "0000000001001110",
8087 => "0000000001001111",
8088 => "0000000001001111",
8089 => "0000000001001111",
8090 => "0000000001001111",
8091 => "0000000001001111",
8092 => "0000000001001111",
8093 => "0000000001001111",
8094 => "0000000001001111",
8095 => "0000000001001111",
8096 => "0000000001001111",
8097 => "0000000001001111",
8098 => "0000000001001111",
8099 => "0000000001001111",
8100 => "0000000001001111",
8101 => "0000000001001111",
8102 => "0000000001001111",
8103 => "0000000001001111",
8104 => "0000000001001111",
8105 => "0000000001001111",
8106 => "0000000001001111",
8107 => "0000000001001111",
8108 => "0000000001001111",
8109 => "0000000001001111",
8110 => "0000000001001111",
8111 => "0000000001001111",
8112 => "0000000001001111",
8113 => "0000000001001111",
8114 => "0000000001001111",
8115 => "0000000001001111",
8116 => "0000000001001111",
8117 => "0000000001001111",
8118 => "0000000001001111",
8119 => "0000000001001111",
8120 => "0000000001001111",
8121 => "0000000001001111",
8122 => "0000000001001111",
8123 => "0000000001001111",
8124 => "0000000001001111",
8125 => "0000000001001111",
8126 => "0000000001001111",
8127 => "0000000001001111",
8128 => "0000000001001111",
8129 => "0000000001001111",
8130 => "0000000001001111",
8131 => "0000000001001111",
8132 => "0000000001001111",
8133 => "0000000001001111",
8134 => "0000000001001111",
8135 => "0000000001001111",
8136 => "0000000001001111",
8137 => "0000000001001111",
8138 => "0000000001001111",
8139 => "0000000001010000",
8140 => "0000000001010000",
8141 => "0000000001010000",
8142 => "0000000001010000",
8143 => "0000000001010000",
8144 => "0000000001010000",
8145 => "0000000001010000",
8146 => "0000000001010000",
8147 => "0000000001010000",
8148 => "0000000001010000",
8149 => "0000000001010000",
8150 => "0000000001010000",
8151 => "0000000001010000",
8152 => "0000000001010000",
8153 => "0000000001010000",
8154 => "0000000001010000",
8155 => "0000000001010000",
8156 => "0000000001010000",
8157 => "0000000001010000",
8158 => "0000000001010000",
8159 => "0000000001010000",
8160 => "0000000001010000",
8161 => "0000000001010000",
8162 => "0000000001010000",
8163 => "0000000001010000",
8164 => "0000000001010000",
8165 => "0000000001010000",
8166 => "0000000001010000",
8167 => "0000000001010000",
8168 => "0000000001010000",
8169 => "0000000001010000",
8170 => "0000000001010000",
8171 => "0000000001010000",
8172 => "0000000001010000",
8173 => "0000000001010000",
8174 => "0000000001010000",
8175 => "0000000001010000",
8176 => "0000000001010000",
8177 => "0000000001010000",
8178 => "0000000001010000",
8179 => "0000000001010000",
8180 => "0000000001010000",
8181 => "0000000001010000",
8182 => "0000000001010000",
8183 => "0000000001010000",
8184 => "0000000001010000",
8185 => "0000000001010000",
8186 => "0000000001010000",
8187 => "0000000001010000",
8188 => "0000000001010000",
8189 => "0000000001010000",
8190 => "0000000001010001",
8191 => "0000000001010001",
8192 => "0000000001010001",
8193 => "0000000001010001",
8194 => "0000000001010001",
8195 => "0000000001010001",
8196 => "0000000001010001",
8197 => "0000000001010001",
8198 => "0000000001010001",
8199 => "0000000001010001",
8200 => "0000000001010001",
8201 => "0000000001010001",
8202 => "0000000001010001",
8203 => "0000000001010001",
8204 => "0000000001010001",
8205 => "0000000001010001",
8206 => "0000000001010001",
8207 => "0000000001010001",
8208 => "0000000001010001",
8209 => "0000000001010001",
8210 => "0000000001010001",
8211 => "0000000001010001",
8212 => "0000000001010001",
8213 => "0000000001010001",
8214 => "0000000001010001",
8215 => "0000000001010001",
8216 => "0000000001010001",
8217 => "0000000001010001",
8218 => "0000000001010001",
8219 => "0000000001010001",
8220 => "0000000001010001",
8221 => "0000000001010001",
8222 => "0000000001010001",
8223 => "0000000001010001",
8224 => "0000000001010001",
8225 => "0000000001010001",
8226 => "0000000001010001",
8227 => "0000000001010001",
8228 => "0000000001010001",
8229 => "0000000001010001",
8230 => "0000000001010001",
8231 => "0000000001010001",
8232 => "0000000001010001",
8233 => "0000000001010001",
8234 => "0000000001010001",
8235 => "0000000001010001",
8236 => "0000000001010001",
8237 => "0000000001010001",
8238 => "0000000001010001",
8239 => "0000000001010001",
8240 => "0000000001010010",
8241 => "0000000001010010",
8242 => "0000000001010010",
8243 => "0000000001010010",
8244 => "0000000001010010",
8245 => "0000000001010010",
8246 => "0000000001010010",
8247 => "0000000001010010",
8248 => "0000000001010010",
8249 => "0000000001010010",
8250 => "0000000001010010",
8251 => "0000000001010010",
8252 => "0000000001010010",
8253 => "0000000001010010",
8254 => "0000000001010010",
8255 => "0000000001010010",
8256 => "0000000001010010",
8257 => "0000000001010010",
8258 => "0000000001010010",
8259 => "0000000001010010",
8260 => "0000000001010010",
8261 => "0000000001010010",
8262 => "0000000001010010",
8263 => "0000000001010010",
8264 => "0000000001010010",
8265 => "0000000001010010",
8266 => "0000000001010010",
8267 => "0000000001010010",
8268 => "0000000001010010",
8269 => "0000000001010010",
8270 => "0000000001010010",
8271 => "0000000001010010",
8272 => "0000000001010010",
8273 => "0000000001010010",
8274 => "0000000001010010",
8275 => "0000000001010010",
8276 => "0000000001010010",
8277 => "0000000001010010",
8278 => "0000000001010010",
8279 => "0000000001010010",
8280 => "0000000001010010",
8281 => "0000000001010010",
8282 => "0000000001010010",
8283 => "0000000001010010",
8284 => "0000000001010010",
8285 => "0000000001010010",
8286 => "0000000001010010",
8287 => "0000000001010010",
8288 => "0000000001010010",
8289 => "0000000001010010",
8290 => "0000000001010011",
8291 => "0000000001010011",
8292 => "0000000001010011",
8293 => "0000000001010011",
8294 => "0000000001010011",
8295 => "0000000001010011",
8296 => "0000000001010011",
8297 => "0000000001010011",
8298 => "0000000001010011",
8299 => "0000000001010011",
8300 => "0000000001010011",
8301 => "0000000001010011",
8302 => "0000000001010011",
8303 => "0000000001010011",
8304 => "0000000001010011",
8305 => "0000000001010011",
8306 => "0000000001010011",
8307 => "0000000001010011",
8308 => "0000000001010011",
8309 => "0000000001010011",
8310 => "0000000001010011",
8311 => "0000000001010011",
8312 => "0000000001010011",
8313 => "0000000001010011",
8314 => "0000000001010011",
8315 => "0000000001010011",
8316 => "0000000001010011",
8317 => "0000000001010011",
8318 => "0000000001010011",
8319 => "0000000001010011",
8320 => "0000000001010011",
8321 => "0000000001010011",
8322 => "0000000001010011",
8323 => "0000000001010011",
8324 => "0000000001010011",
8325 => "0000000001010011",
8326 => "0000000001010011",
8327 => "0000000001010011",
8328 => "0000000001010011",
8329 => "0000000001010011",
8330 => "0000000001010011",
8331 => "0000000001010011",
8332 => "0000000001010011",
8333 => "0000000001010011",
8334 => "0000000001010011",
8335 => "0000000001010011",
8336 => "0000000001010011",
8337 => "0000000001010011",
8338 => "0000000001010011",
8339 => "0000000001010100",
8340 => "0000000001010100",
8341 => "0000000001010100",
8342 => "0000000001010100",
8343 => "0000000001010100",
8344 => "0000000001010100",
8345 => "0000000001010100",
8346 => "0000000001010100",
8347 => "0000000001010100",
8348 => "0000000001010100",
8349 => "0000000001010100",
8350 => "0000000001010100",
8351 => "0000000001010100",
8352 => "0000000001010100",
8353 => "0000000001010100",
8354 => "0000000001010100",
8355 => "0000000001010100",
8356 => "0000000001010100",
8357 => "0000000001010100",
8358 => "0000000001010100",
8359 => "0000000001010100",
8360 => "0000000001010100",
8361 => "0000000001010100",
8362 => "0000000001010100",
8363 => "0000000001010100",
8364 => "0000000001010100",
8365 => "0000000001010100",
8366 => "0000000001010100",
8367 => "0000000001010100",
8368 => "0000000001010100",
8369 => "0000000001010100",
8370 => "0000000001010100",
8371 => "0000000001010100",
8372 => "0000000001010100",
8373 => "0000000001010100",
8374 => "0000000001010100",
8375 => "0000000001010100",
8376 => "0000000001010100",
8377 => "0000000001010100",
8378 => "0000000001010100",
8379 => "0000000001010100",
8380 => "0000000001010100",
8381 => "0000000001010100",
8382 => "0000000001010100",
8383 => "0000000001010100",
8384 => "0000000001010100",
8385 => "0000000001010100",
8386 => "0000000001010100",
8387 => "0000000001010100",
8388 => "0000000001010101",
8389 => "0000000001010101",
8390 => "0000000001010101",
8391 => "0000000001010101",
8392 => "0000000001010101",
8393 => "0000000001010101",
8394 => "0000000001010101",
8395 => "0000000001010101",
8396 => "0000000001010101",
8397 => "0000000001010101",
8398 => "0000000001010101",
8399 => "0000000001010101",
8400 => "0000000001010101",
8401 => "0000000001010101",
8402 => "0000000001010101",
8403 => "0000000001010101",
8404 => "0000000001010101",
8405 => "0000000001010101",
8406 => "0000000001010101",
8407 => "0000000001010101",
8408 => "0000000001010101",
8409 => "0000000001010101",
8410 => "0000000001010101",
8411 => "0000000001010101",
8412 => "0000000001010101",
8413 => "0000000001010101",
8414 => "0000000001010101",
8415 => "0000000001010101",
8416 => "0000000001010101",
8417 => "0000000001010101",
8418 => "0000000001010101",
8419 => "0000000001010101",
8420 => "0000000001010101",
8421 => "0000000001010101",
8422 => "0000000001010101",
8423 => "0000000001010101",
8424 => "0000000001010101",
8425 => "0000000001010101",
8426 => "0000000001010101",
8427 => "0000000001010101",
8428 => "0000000001010101",
8429 => "0000000001010101",
8430 => "0000000001010101",
8431 => "0000000001010101",
8432 => "0000000001010101",
8433 => "0000000001010101",
8434 => "0000000001010101",
8435 => "0000000001010101",
8436 => "0000000001010110",
8437 => "0000000001010110",
8438 => "0000000001010110",
8439 => "0000000001010110",
8440 => "0000000001010110",
8441 => "0000000001010110",
8442 => "0000000001010110",
8443 => "0000000001010110",
8444 => "0000000001010110",
8445 => "0000000001010110",
8446 => "0000000001010110",
8447 => "0000000001010110",
8448 => "0000000001010110",
8449 => "0000000001010110",
8450 => "0000000001010110",
8451 => "0000000001010110",
8452 => "0000000001010110",
8453 => "0000000001010110",
8454 => "0000000001010110",
8455 => "0000000001010110",
8456 => "0000000001010110",
8457 => "0000000001010110",
8458 => "0000000001010110",
8459 => "0000000001010110",
8460 => "0000000001010110",
8461 => "0000000001010110",
8462 => "0000000001010110",
8463 => "0000000001010110",
8464 => "0000000001010110",
8465 => "0000000001010110",
8466 => "0000000001010110",
8467 => "0000000001010110",
8468 => "0000000001010110",
8469 => "0000000001010110",
8470 => "0000000001010110",
8471 => "0000000001010110",
8472 => "0000000001010110",
8473 => "0000000001010110",
8474 => "0000000001010110",
8475 => "0000000001010110",
8476 => "0000000001010110",
8477 => "0000000001010110",
8478 => "0000000001010110",
8479 => "0000000001010110",
8480 => "0000000001010110",
8481 => "0000000001010110",
8482 => "0000000001010110",
8483 => "0000000001010111",
8484 => "0000000001010111",
8485 => "0000000001010111",
8486 => "0000000001010111",
8487 => "0000000001010111",
8488 => "0000000001010111",
8489 => "0000000001010111",
8490 => "0000000001010111",
8491 => "0000000001010111",
8492 => "0000000001010111",
8493 => "0000000001010111",
8494 => "0000000001010111",
8495 => "0000000001010111",
8496 => "0000000001010111",
8497 => "0000000001010111",
8498 => "0000000001010111",
8499 => "0000000001010111",
8500 => "0000000001010111",
8501 => "0000000001010111",
8502 => "0000000001010111",
8503 => "0000000001010111",
8504 => "0000000001010111",
8505 => "0000000001010111",
8506 => "0000000001010111",
8507 => "0000000001010111",
8508 => "0000000001010111",
8509 => "0000000001010111",
8510 => "0000000001010111",
8511 => "0000000001010111",
8512 => "0000000001010111",
8513 => "0000000001010111",
8514 => "0000000001010111",
8515 => "0000000001010111",
8516 => "0000000001010111",
8517 => "0000000001010111",
8518 => "0000000001010111",
8519 => "0000000001010111",
8520 => "0000000001010111",
8521 => "0000000001010111",
8522 => "0000000001010111",
8523 => "0000000001010111",
8524 => "0000000001010111",
8525 => "0000000001010111",
8526 => "0000000001010111",
8527 => "0000000001010111",
8528 => "0000000001010111",
8529 => "0000000001010111",
8530 => "0000000001011000",
8531 => "0000000001011000",
8532 => "0000000001011000",
8533 => "0000000001011000",
8534 => "0000000001011000",
8535 => "0000000001011000",
8536 => "0000000001011000",
8537 => "0000000001011000",
8538 => "0000000001011000",
8539 => "0000000001011000",
8540 => "0000000001011000",
8541 => "0000000001011000",
8542 => "0000000001011000",
8543 => "0000000001011000",
8544 => "0000000001011000",
8545 => "0000000001011000",
8546 => "0000000001011000",
8547 => "0000000001011000",
8548 => "0000000001011000",
8549 => "0000000001011000",
8550 => "0000000001011000",
8551 => "0000000001011000",
8552 => "0000000001011000",
8553 => "0000000001011000",
8554 => "0000000001011000",
8555 => "0000000001011000",
8556 => "0000000001011000",
8557 => "0000000001011000",
8558 => "0000000001011000",
8559 => "0000000001011000",
8560 => "0000000001011000",
8561 => "0000000001011000",
8562 => "0000000001011000",
8563 => "0000000001011000",
8564 => "0000000001011000",
8565 => "0000000001011000",
8566 => "0000000001011000",
8567 => "0000000001011000",
8568 => "0000000001011000",
8569 => "0000000001011000",
8570 => "0000000001011000",
8571 => "0000000001011000",
8572 => "0000000001011000",
8573 => "0000000001011000",
8574 => "0000000001011000",
8575 => "0000000001011000",
8576 => "0000000001011000",
8577 => "0000000001011001",
8578 => "0000000001011001",
8579 => "0000000001011001",
8580 => "0000000001011001",
8581 => "0000000001011001",
8582 => "0000000001011001",
8583 => "0000000001011001",
8584 => "0000000001011001",
8585 => "0000000001011001",
8586 => "0000000001011001",
8587 => "0000000001011001",
8588 => "0000000001011001",
8589 => "0000000001011001",
8590 => "0000000001011001",
8591 => "0000000001011001",
8592 => "0000000001011001",
8593 => "0000000001011001",
8594 => "0000000001011001",
8595 => "0000000001011001",
8596 => "0000000001011001",
8597 => "0000000001011001",
8598 => "0000000001011001",
8599 => "0000000001011001",
8600 => "0000000001011001",
8601 => "0000000001011001",
8602 => "0000000001011001",
8603 => "0000000001011001",
8604 => "0000000001011001",
8605 => "0000000001011001",
8606 => "0000000001011001",
8607 => "0000000001011001",
8608 => "0000000001011001",
8609 => "0000000001011001",
8610 => "0000000001011001",
8611 => "0000000001011001",
8612 => "0000000001011001",
8613 => "0000000001011001",
8614 => "0000000001011001",
8615 => "0000000001011001",
8616 => "0000000001011001",
8617 => "0000000001011001",
8618 => "0000000001011001",
8619 => "0000000001011001",
8620 => "0000000001011001",
8621 => "0000000001011001",
8622 => "0000000001011010",
8623 => "0000000001011010",
8624 => "0000000001011010",
8625 => "0000000001011010",
8626 => "0000000001011010",
8627 => "0000000001011010",
8628 => "0000000001011010",
8629 => "0000000001011010",
8630 => "0000000001011010",
8631 => "0000000001011010",
8632 => "0000000001011010",
8633 => "0000000001011010",
8634 => "0000000001011010",
8635 => "0000000001011010",
8636 => "0000000001011010",
8637 => "0000000001011010",
8638 => "0000000001011010",
8639 => "0000000001011010",
8640 => "0000000001011010",
8641 => "0000000001011010",
8642 => "0000000001011010",
8643 => "0000000001011010",
8644 => "0000000001011010",
8645 => "0000000001011010",
8646 => "0000000001011010",
8647 => "0000000001011010",
8648 => "0000000001011010",
8649 => "0000000001011010",
8650 => "0000000001011010",
8651 => "0000000001011010",
8652 => "0000000001011010",
8653 => "0000000001011010",
8654 => "0000000001011010",
8655 => "0000000001011010",
8656 => "0000000001011010",
8657 => "0000000001011010",
8658 => "0000000001011010",
8659 => "0000000001011010",
8660 => "0000000001011010",
8661 => "0000000001011010",
8662 => "0000000001011010",
8663 => "0000000001011010",
8664 => "0000000001011010",
8665 => "0000000001011010",
8666 => "0000000001011010",
8667 => "0000000001011010",
8668 => "0000000001011011",
8669 => "0000000001011011",
8670 => "0000000001011011",
8671 => "0000000001011011",
8672 => "0000000001011011",
8673 => "0000000001011011",
8674 => "0000000001011011",
8675 => "0000000001011011",
8676 => "0000000001011011",
8677 => "0000000001011011",
8678 => "0000000001011011",
8679 => "0000000001011011",
8680 => "0000000001011011",
8681 => "0000000001011011",
8682 => "0000000001011011",
8683 => "0000000001011011",
8684 => "0000000001011011",
8685 => "0000000001011011",
8686 => "0000000001011011",
8687 => "0000000001011011",
8688 => "0000000001011011",
8689 => "0000000001011011",
8690 => "0000000001011011",
8691 => "0000000001011011",
8692 => "0000000001011011",
8693 => "0000000001011011",
8694 => "0000000001011011",
8695 => "0000000001011011",
8696 => "0000000001011011",
8697 => "0000000001011011",
8698 => "0000000001011011",
8699 => "0000000001011011",
8700 => "0000000001011011",
8701 => "0000000001011011",
8702 => "0000000001011011",
8703 => "0000000001011011",
8704 => "0000000001011011",
8705 => "0000000001011011",
8706 => "0000000001011011",
8707 => "0000000001011011",
8708 => "0000000001011011",
8709 => "0000000001011011",
8710 => "0000000001011011",
8711 => "0000000001011011",
8712 => "0000000001011011",
8713 => "0000000001011100",
8714 => "0000000001011100",
8715 => "0000000001011100",
8716 => "0000000001011100",
8717 => "0000000001011100",
8718 => "0000000001011100",
8719 => "0000000001011100",
8720 => "0000000001011100",
8721 => "0000000001011100",
8722 => "0000000001011100",
8723 => "0000000001011100",
8724 => "0000000001011100",
8725 => "0000000001011100",
8726 => "0000000001011100",
8727 => "0000000001011100",
8728 => "0000000001011100",
8729 => "0000000001011100",
8730 => "0000000001011100",
8731 => "0000000001011100",
8732 => "0000000001011100",
8733 => "0000000001011100",
8734 => "0000000001011100",
8735 => "0000000001011100",
8736 => "0000000001011100",
8737 => "0000000001011100",
8738 => "0000000001011100",
8739 => "0000000001011100",
8740 => "0000000001011100",
8741 => "0000000001011100",
8742 => "0000000001011100",
8743 => "0000000001011100",
8744 => "0000000001011100",
8745 => "0000000001011100",
8746 => "0000000001011100",
8747 => "0000000001011100",
8748 => "0000000001011100",
8749 => "0000000001011100",
8750 => "0000000001011100",
8751 => "0000000001011100",
8752 => "0000000001011100",
8753 => "0000000001011100",
8754 => "0000000001011100",
8755 => "0000000001011100",
8756 => "0000000001011100",
8757 => "0000000001011101",
8758 => "0000000001011101",
8759 => "0000000001011101",
8760 => "0000000001011101",
8761 => "0000000001011101",
8762 => "0000000001011101",
8763 => "0000000001011101",
8764 => "0000000001011101",
8765 => "0000000001011101",
8766 => "0000000001011101",
8767 => "0000000001011101",
8768 => "0000000001011101",
8769 => "0000000001011101",
8770 => "0000000001011101",
8771 => "0000000001011101",
8772 => "0000000001011101",
8773 => "0000000001011101",
8774 => "0000000001011101",
8775 => "0000000001011101",
8776 => "0000000001011101",
8777 => "0000000001011101",
8778 => "0000000001011101",
8779 => "0000000001011101",
8780 => "0000000001011101",
8781 => "0000000001011101",
8782 => "0000000001011101",
8783 => "0000000001011101",
8784 => "0000000001011101",
8785 => "0000000001011101",
8786 => "0000000001011101",
8787 => "0000000001011101",
8788 => "0000000001011101",
8789 => "0000000001011101",
8790 => "0000000001011101",
8791 => "0000000001011101",
8792 => "0000000001011101",
8793 => "0000000001011101",
8794 => "0000000001011101",
8795 => "0000000001011101",
8796 => "0000000001011101",
8797 => "0000000001011101",
8798 => "0000000001011101",
8799 => "0000000001011101",
8800 => "0000000001011101",
8801 => "0000000001011110",
8802 => "0000000001011110",
8803 => "0000000001011110",
8804 => "0000000001011110",
8805 => "0000000001011110",
8806 => "0000000001011110",
8807 => "0000000001011110",
8808 => "0000000001011110",
8809 => "0000000001011110",
8810 => "0000000001011110",
8811 => "0000000001011110",
8812 => "0000000001011110",
8813 => "0000000001011110",
8814 => "0000000001011110",
8815 => "0000000001011110",
8816 => "0000000001011110",
8817 => "0000000001011110",
8818 => "0000000001011110",
8819 => "0000000001011110",
8820 => "0000000001011110",
8821 => "0000000001011110",
8822 => "0000000001011110",
8823 => "0000000001011110",
8824 => "0000000001011110",
8825 => "0000000001011110",
8826 => "0000000001011110",
8827 => "0000000001011110",
8828 => "0000000001011110",
8829 => "0000000001011110",
8830 => "0000000001011110",
8831 => "0000000001011110",
8832 => "0000000001011110",
8833 => "0000000001011110",
8834 => "0000000001011110",
8835 => "0000000001011110",
8836 => "0000000001011110",
8837 => "0000000001011110",
8838 => "0000000001011110",
8839 => "0000000001011110",
8840 => "0000000001011110",
8841 => "0000000001011110",
8842 => "0000000001011110",
8843 => "0000000001011110",
8844 => "0000000001011110",
8845 => "0000000001011111",
8846 => "0000000001011111",
8847 => "0000000001011111",
8848 => "0000000001011111",
8849 => "0000000001011111",
8850 => "0000000001011111",
8851 => "0000000001011111",
8852 => "0000000001011111",
8853 => "0000000001011111",
8854 => "0000000001011111",
8855 => "0000000001011111",
8856 => "0000000001011111",
8857 => "0000000001011111",
8858 => "0000000001011111",
8859 => "0000000001011111",
8860 => "0000000001011111",
8861 => "0000000001011111",
8862 => "0000000001011111",
8863 => "0000000001011111",
8864 => "0000000001011111",
8865 => "0000000001011111",
8866 => "0000000001011111",
8867 => "0000000001011111",
8868 => "0000000001011111",
8869 => "0000000001011111",
8870 => "0000000001011111",
8871 => "0000000001011111",
8872 => "0000000001011111",
8873 => "0000000001011111",
8874 => "0000000001011111",
8875 => "0000000001011111",
8876 => "0000000001011111",
8877 => "0000000001011111",
8878 => "0000000001011111",
8879 => "0000000001011111",
8880 => "0000000001011111",
8881 => "0000000001011111",
8882 => "0000000001011111",
8883 => "0000000001011111",
8884 => "0000000001011111",
8885 => "0000000001011111",
8886 => "0000000001011111",
8887 => "0000000001011111",
8888 => "0000000001100000",
8889 => "0000000001100000",
8890 => "0000000001100000",
8891 => "0000000001100000",
8892 => "0000000001100000",
8893 => "0000000001100000",
8894 => "0000000001100000",
8895 => "0000000001100000",
8896 => "0000000001100000",
8897 => "0000000001100000",
8898 => "0000000001100000",
8899 => "0000000001100000",
8900 => "0000000001100000",
8901 => "0000000001100000",
8902 => "0000000001100000",
8903 => "0000000001100000",
8904 => "0000000001100000",
8905 => "0000000001100000",
8906 => "0000000001100000",
8907 => "0000000001100000",
8908 => "0000000001100000",
8909 => "0000000001100000",
8910 => "0000000001100000",
8911 => "0000000001100000",
8912 => "0000000001100000",
8913 => "0000000001100000",
8914 => "0000000001100000",
8915 => "0000000001100000",
8916 => "0000000001100000",
8917 => "0000000001100000",
8918 => "0000000001100000",
8919 => "0000000001100000",
8920 => "0000000001100000",
8921 => "0000000001100000",
8922 => "0000000001100000",
8923 => "0000000001100000",
8924 => "0000000001100000",
8925 => "0000000001100000",
8926 => "0000000001100000",
8927 => "0000000001100000",
8928 => "0000000001100000",
8929 => "0000000001100000",
8930 => "0000000001100001",
8931 => "0000000001100001",
8932 => "0000000001100001",
8933 => "0000000001100001",
8934 => "0000000001100001",
8935 => "0000000001100001",
8936 => "0000000001100001",
8937 => "0000000001100001",
8938 => "0000000001100001",
8939 => "0000000001100001",
8940 => "0000000001100001",
8941 => "0000000001100001",
8942 => "0000000001100001",
8943 => "0000000001100001",
8944 => "0000000001100001",
8945 => "0000000001100001",
8946 => "0000000001100001",
8947 => "0000000001100001",
8948 => "0000000001100001",
8949 => "0000000001100001",
8950 => "0000000001100001",
8951 => "0000000001100001",
8952 => "0000000001100001",
8953 => "0000000001100001",
8954 => "0000000001100001",
8955 => "0000000001100001",
8956 => "0000000001100001",
8957 => "0000000001100001",
8958 => "0000000001100001",
8959 => "0000000001100001",
8960 => "0000000001100001",
8961 => "0000000001100001",
8962 => "0000000001100001",
8963 => "0000000001100001",
8964 => "0000000001100001",
8965 => "0000000001100001",
8966 => "0000000001100001",
8967 => "0000000001100001",
8968 => "0000000001100001",
8969 => "0000000001100001",
8970 => "0000000001100001",
8971 => "0000000001100001",
8972 => "0000000001100010",
8973 => "0000000001100010",
8974 => "0000000001100010",
8975 => "0000000001100010",
8976 => "0000000001100010",
8977 => "0000000001100010",
8978 => "0000000001100010",
8979 => "0000000001100010",
8980 => "0000000001100010",
8981 => "0000000001100010",
8982 => "0000000001100010",
8983 => "0000000001100010",
8984 => "0000000001100010",
8985 => "0000000001100010",
8986 => "0000000001100010",
8987 => "0000000001100010",
8988 => "0000000001100010",
8989 => "0000000001100010",
8990 => "0000000001100010",
8991 => "0000000001100010",
8992 => "0000000001100010",
8993 => "0000000001100010",
8994 => "0000000001100010",
8995 => "0000000001100010",
8996 => "0000000001100010",
8997 => "0000000001100010",
8998 => "0000000001100010",
8999 => "0000000001100010",
9000 => "0000000001100010",
9001 => "0000000001100010",
9002 => "0000000001100010",
9003 => "0000000001100010",
9004 => "0000000001100010",
9005 => "0000000001100010",
9006 => "0000000001100010",
9007 => "0000000001100010",
9008 => "0000000001100010",
9009 => "0000000001100010",
9010 => "0000000001100010",
9011 => "0000000001100010",
9012 => "0000000001100010",
9013 => "0000000001100010",
9014 => "0000000001100011",
9015 => "0000000001100011",
9016 => "0000000001100011",
9017 => "0000000001100011",
9018 => "0000000001100011",
9019 => "0000000001100011",
9020 => "0000000001100011",
9021 => "0000000001100011",
9022 => "0000000001100011",
9023 => "0000000001100011",
9024 => "0000000001100011",
9025 => "0000000001100011",
9026 => "0000000001100011",
9027 => "0000000001100011",
9028 => "0000000001100011",
9029 => "0000000001100011",
9030 => "0000000001100011",
9031 => "0000000001100011",
9032 => "0000000001100011",
9033 => "0000000001100011",
9034 => "0000000001100011",
9035 => "0000000001100011",
9036 => "0000000001100011",
9037 => "0000000001100011",
9038 => "0000000001100011",
9039 => "0000000001100011",
9040 => "0000000001100011",
9041 => "0000000001100011",
9042 => "0000000001100011",
9043 => "0000000001100011",
9044 => "0000000001100011",
9045 => "0000000001100011",
9046 => "0000000001100011",
9047 => "0000000001100011",
9048 => "0000000001100011",
9049 => "0000000001100011",
9050 => "0000000001100011",
9051 => "0000000001100011",
9052 => "0000000001100011",
9053 => "0000000001100011",
9054 => "0000000001100011",
9055 => "0000000001100100",
9056 => "0000000001100100",
9057 => "0000000001100100",
9058 => "0000000001100100",
9059 => "0000000001100100",
9060 => "0000000001100100",
9061 => "0000000001100100",
9062 => "0000000001100100",
9063 => "0000000001100100",
9064 => "0000000001100100",
9065 => "0000000001100100",
9066 => "0000000001100100",
9067 => "0000000001100100",
9068 => "0000000001100100",
9069 => "0000000001100100",
9070 => "0000000001100100",
9071 => "0000000001100100",
9072 => "0000000001100100",
9073 => "0000000001100100",
9074 => "0000000001100100",
9075 => "0000000001100100",
9076 => "0000000001100100",
9077 => "0000000001100100",
9078 => "0000000001100100",
9079 => "0000000001100100",
9080 => "0000000001100100",
9081 => "0000000001100100",
9082 => "0000000001100100",
9083 => "0000000001100100",
9084 => "0000000001100100",
9085 => "0000000001100100",
9086 => "0000000001100100",
9087 => "0000000001100100",
9088 => "0000000001100100",
9089 => "0000000001100100",
9090 => "0000000001100100",
9091 => "0000000001100100",
9092 => "0000000001100100",
9093 => "0000000001100100",
9094 => "0000000001100100",
9095 => "0000000001100100",
9096 => "0000000001100101",
9097 => "0000000001100101",
9098 => "0000000001100101",
9099 => "0000000001100101",
9100 => "0000000001100101",
9101 => "0000000001100101",
9102 => "0000000001100101",
9103 => "0000000001100101",
9104 => "0000000001100101",
9105 => "0000000001100101",
9106 => "0000000001100101",
9107 => "0000000001100101",
9108 => "0000000001100101",
9109 => "0000000001100101",
9110 => "0000000001100101",
9111 => "0000000001100101",
9112 => "0000000001100101",
9113 => "0000000001100101",
9114 => "0000000001100101",
9115 => "0000000001100101",
9116 => "0000000001100101",
9117 => "0000000001100101",
9118 => "0000000001100101",
9119 => "0000000001100101",
9120 => "0000000001100101",
9121 => "0000000001100101",
9122 => "0000000001100101",
9123 => "0000000001100101",
9124 => "0000000001100101",
9125 => "0000000001100101",
9126 => "0000000001100101",
9127 => "0000000001100101",
9128 => "0000000001100101",
9129 => "0000000001100101",
9130 => "0000000001100101",
9131 => "0000000001100101",
9132 => "0000000001100101",
9133 => "0000000001100101",
9134 => "0000000001100101",
9135 => "0000000001100101",
9136 => "0000000001100101",
9137 => "0000000001100110",
9138 => "0000000001100110",
9139 => "0000000001100110",
9140 => "0000000001100110",
9141 => "0000000001100110",
9142 => "0000000001100110",
9143 => "0000000001100110",
9144 => "0000000001100110",
9145 => "0000000001100110",
9146 => "0000000001100110",
9147 => "0000000001100110",
9148 => "0000000001100110",
9149 => "0000000001100110",
9150 => "0000000001100110",
9151 => "0000000001100110",
9152 => "0000000001100110",
9153 => "0000000001100110",
9154 => "0000000001100110",
9155 => "0000000001100110",
9156 => "0000000001100110",
9157 => "0000000001100110",
9158 => "0000000001100110",
9159 => "0000000001100110",
9160 => "0000000001100110",
9161 => "0000000001100110",
9162 => "0000000001100110",
9163 => "0000000001100110",
9164 => "0000000001100110",
9165 => "0000000001100110",
9166 => "0000000001100110",
9167 => "0000000001100110",
9168 => "0000000001100110",
9169 => "0000000001100110",
9170 => "0000000001100110",
9171 => "0000000001100110",
9172 => "0000000001100110",
9173 => "0000000001100110",
9174 => "0000000001100110",
9175 => "0000000001100110",
9176 => "0000000001100110",
9177 => "0000000001100111",
9178 => "0000000001100111",
9179 => "0000000001100111",
9180 => "0000000001100111",
9181 => "0000000001100111",
9182 => "0000000001100111",
9183 => "0000000001100111",
9184 => "0000000001100111",
9185 => "0000000001100111",
9186 => "0000000001100111",
9187 => "0000000001100111",
9188 => "0000000001100111",
9189 => "0000000001100111",
9190 => "0000000001100111",
9191 => "0000000001100111",
9192 => "0000000001100111",
9193 => "0000000001100111",
9194 => "0000000001100111",
9195 => "0000000001100111",
9196 => "0000000001100111",
9197 => "0000000001100111",
9198 => "0000000001100111",
9199 => "0000000001100111",
9200 => "0000000001100111",
9201 => "0000000001100111",
9202 => "0000000001100111",
9203 => "0000000001100111",
9204 => "0000000001100111",
9205 => "0000000001100111",
9206 => "0000000001100111",
9207 => "0000000001100111",
9208 => "0000000001100111",
9209 => "0000000001100111",
9210 => "0000000001100111",
9211 => "0000000001100111",
9212 => "0000000001100111",
9213 => "0000000001100111",
9214 => "0000000001100111",
9215 => "0000000001100111",
9216 => "0000000001100111",
9217 => "0000000001101000",
9218 => "0000000001101000",
9219 => "0000000001101000",
9220 => "0000000001101000",
9221 => "0000000001101000",
9222 => "0000000001101000",
9223 => "0000000001101000",
9224 => "0000000001101000",
9225 => "0000000001101000",
9226 => "0000000001101000",
9227 => "0000000001101000",
9228 => "0000000001101000",
9229 => "0000000001101000",
9230 => "0000000001101000",
9231 => "0000000001101000",
9232 => "0000000001101000",
9233 => "0000000001101000",
9234 => "0000000001101000",
9235 => "0000000001101000",
9236 => "0000000001101000",
9237 => "0000000001101000",
9238 => "0000000001101000",
9239 => "0000000001101000",
9240 => "0000000001101000",
9241 => "0000000001101000",
9242 => "0000000001101000",
9243 => "0000000001101000",
9244 => "0000000001101000",
9245 => "0000000001101000",
9246 => "0000000001101000",
9247 => "0000000001101000",
9248 => "0000000001101000",
9249 => "0000000001101000",
9250 => "0000000001101000",
9251 => "0000000001101000",
9252 => "0000000001101000",
9253 => "0000000001101000",
9254 => "0000000001101000",
9255 => "0000000001101000",
9256 => "0000000001101001",
9257 => "0000000001101001",
9258 => "0000000001101001",
9259 => "0000000001101001",
9260 => "0000000001101001",
9261 => "0000000001101001",
9262 => "0000000001101001",
9263 => "0000000001101001",
9264 => "0000000001101001",
9265 => "0000000001101001",
9266 => "0000000001101001",
9267 => "0000000001101001",
9268 => "0000000001101001",
9269 => "0000000001101001",
9270 => "0000000001101001",
9271 => "0000000001101001",
9272 => "0000000001101001",
9273 => "0000000001101001",
9274 => "0000000001101001",
9275 => "0000000001101001",
9276 => "0000000001101001",
9277 => "0000000001101001",
9278 => "0000000001101001",
9279 => "0000000001101001",
9280 => "0000000001101001",
9281 => "0000000001101001",
9282 => "0000000001101001",
9283 => "0000000001101001",
9284 => "0000000001101001",
9285 => "0000000001101001",
9286 => "0000000001101001",
9287 => "0000000001101001",
9288 => "0000000001101001",
9289 => "0000000001101001",
9290 => "0000000001101001",
9291 => "0000000001101001",
9292 => "0000000001101001",
9293 => "0000000001101001",
9294 => "0000000001101001",
9295 => "0000000001101010",
9296 => "0000000001101010",
9297 => "0000000001101010",
9298 => "0000000001101010",
9299 => "0000000001101010",
9300 => "0000000001101010",
9301 => "0000000001101010",
9302 => "0000000001101010",
9303 => "0000000001101010",
9304 => "0000000001101010",
9305 => "0000000001101010",
9306 => "0000000001101010",
9307 => "0000000001101010",
9308 => "0000000001101010",
9309 => "0000000001101010",
9310 => "0000000001101010",
9311 => "0000000001101010",
9312 => "0000000001101010",
9313 => "0000000001101010",
9314 => "0000000001101010",
9315 => "0000000001101010",
9316 => "0000000001101010",
9317 => "0000000001101010",
9318 => "0000000001101010",
9319 => "0000000001101010",
9320 => "0000000001101010",
9321 => "0000000001101010",
9322 => "0000000001101010",
9323 => "0000000001101010",
9324 => "0000000001101010",
9325 => "0000000001101010",
9326 => "0000000001101010",
9327 => "0000000001101010",
9328 => "0000000001101010",
9329 => "0000000001101010",
9330 => "0000000001101010",
9331 => "0000000001101010",
9332 => "0000000001101010",
9333 => "0000000001101011",
9334 => "0000000001101011",
9335 => "0000000001101011",
9336 => "0000000001101011",
9337 => "0000000001101011",
9338 => "0000000001101011",
9339 => "0000000001101011",
9340 => "0000000001101011",
9341 => "0000000001101011",
9342 => "0000000001101011",
9343 => "0000000001101011",
9344 => "0000000001101011",
9345 => "0000000001101011",
9346 => "0000000001101011",
9347 => "0000000001101011",
9348 => "0000000001101011",
9349 => "0000000001101011",
9350 => "0000000001101011",
9351 => "0000000001101011",
9352 => "0000000001101011",
9353 => "0000000001101011",
9354 => "0000000001101011",
9355 => "0000000001101011",
9356 => "0000000001101011",
9357 => "0000000001101011",
9358 => "0000000001101011",
9359 => "0000000001101011",
9360 => "0000000001101011",
9361 => "0000000001101011",
9362 => "0000000001101011",
9363 => "0000000001101011",
9364 => "0000000001101011",
9365 => "0000000001101011",
9366 => "0000000001101011",
9367 => "0000000001101011",
9368 => "0000000001101011",
9369 => "0000000001101011",
9370 => "0000000001101011",
9371 => "0000000001101011",
9372 => "0000000001101100",
9373 => "0000000001101100",
9374 => "0000000001101100",
9375 => "0000000001101100",
9376 => "0000000001101100",
9377 => "0000000001101100",
9378 => "0000000001101100",
9379 => "0000000001101100",
9380 => "0000000001101100",
9381 => "0000000001101100",
9382 => "0000000001101100",
9383 => "0000000001101100",
9384 => "0000000001101100",
9385 => "0000000001101100",
9386 => "0000000001101100",
9387 => "0000000001101100",
9388 => "0000000001101100",
9389 => "0000000001101100",
9390 => "0000000001101100",
9391 => "0000000001101100",
9392 => "0000000001101100",
9393 => "0000000001101100",
9394 => "0000000001101100",
9395 => "0000000001101100",
9396 => "0000000001101100",
9397 => "0000000001101100",
9398 => "0000000001101100",
9399 => "0000000001101100",
9400 => "0000000001101100",
9401 => "0000000001101100",
9402 => "0000000001101100",
9403 => "0000000001101100",
9404 => "0000000001101100",
9405 => "0000000001101100",
9406 => "0000000001101100",
9407 => "0000000001101100",
9408 => "0000000001101100",
9409 => "0000000001101100",
9410 => "0000000001101101",
9411 => "0000000001101101",
9412 => "0000000001101101",
9413 => "0000000001101101",
9414 => "0000000001101101",
9415 => "0000000001101101",
9416 => "0000000001101101",
9417 => "0000000001101101",
9418 => "0000000001101101",
9419 => "0000000001101101",
9420 => "0000000001101101",
9421 => "0000000001101101",
9422 => "0000000001101101",
9423 => "0000000001101101",
9424 => "0000000001101101",
9425 => "0000000001101101",
9426 => "0000000001101101",
9427 => "0000000001101101",
9428 => "0000000001101101",
9429 => "0000000001101101",
9430 => "0000000001101101",
9431 => "0000000001101101",
9432 => "0000000001101101",
9433 => "0000000001101101",
9434 => "0000000001101101",
9435 => "0000000001101101",
9436 => "0000000001101101",
9437 => "0000000001101101",
9438 => "0000000001101101",
9439 => "0000000001101101",
9440 => "0000000001101101",
9441 => "0000000001101101",
9442 => "0000000001101101",
9443 => "0000000001101101",
9444 => "0000000001101101",
9445 => "0000000001101101",
9446 => "0000000001101101",
9447 => "0000000001101110",
9448 => "0000000001101110",
9449 => "0000000001101110",
9450 => "0000000001101110",
9451 => "0000000001101110",
9452 => "0000000001101110",
9453 => "0000000001101110",
9454 => "0000000001101110",
9455 => "0000000001101110",
9456 => "0000000001101110",
9457 => "0000000001101110",
9458 => "0000000001101110",
9459 => "0000000001101110",
9460 => "0000000001101110",
9461 => "0000000001101110",
9462 => "0000000001101110",
9463 => "0000000001101110",
9464 => "0000000001101110",
9465 => "0000000001101110",
9466 => "0000000001101110",
9467 => "0000000001101110",
9468 => "0000000001101110",
9469 => "0000000001101110",
9470 => "0000000001101110",
9471 => "0000000001101110",
9472 => "0000000001101110",
9473 => "0000000001101110",
9474 => "0000000001101110",
9475 => "0000000001101110",
9476 => "0000000001101110",
9477 => "0000000001101110",
9478 => "0000000001101110",
9479 => "0000000001101110",
9480 => "0000000001101110",
9481 => "0000000001101110",
9482 => "0000000001101110",
9483 => "0000000001101110",
9484 => "0000000001101111",
9485 => "0000000001101111",
9486 => "0000000001101111",
9487 => "0000000001101111",
9488 => "0000000001101111",
9489 => "0000000001101111",
9490 => "0000000001101111",
9491 => "0000000001101111",
9492 => "0000000001101111",
9493 => "0000000001101111",
9494 => "0000000001101111",
9495 => "0000000001101111",
9496 => "0000000001101111",
9497 => "0000000001101111",
9498 => "0000000001101111",
9499 => "0000000001101111",
9500 => "0000000001101111",
9501 => "0000000001101111",
9502 => "0000000001101111",
9503 => "0000000001101111",
9504 => "0000000001101111",
9505 => "0000000001101111",
9506 => "0000000001101111",
9507 => "0000000001101111",
9508 => "0000000001101111",
9509 => "0000000001101111",
9510 => "0000000001101111",
9511 => "0000000001101111",
9512 => "0000000001101111",
9513 => "0000000001101111",
9514 => "0000000001101111",
9515 => "0000000001101111",
9516 => "0000000001101111",
9517 => "0000000001101111",
9518 => "0000000001101111",
9519 => "0000000001101111",
9520 => "0000000001101111",
9521 => "0000000001110000",
9522 => "0000000001110000",
9523 => "0000000001110000",
9524 => "0000000001110000",
9525 => "0000000001110000",
9526 => "0000000001110000",
9527 => "0000000001110000",
9528 => "0000000001110000",
9529 => "0000000001110000",
9530 => "0000000001110000",
9531 => "0000000001110000",
9532 => "0000000001110000",
9533 => "0000000001110000",
9534 => "0000000001110000",
9535 => "0000000001110000",
9536 => "0000000001110000",
9537 => "0000000001110000",
9538 => "0000000001110000",
9539 => "0000000001110000",
9540 => "0000000001110000",
9541 => "0000000001110000",
9542 => "0000000001110000",
9543 => "0000000001110000",
9544 => "0000000001110000",
9545 => "0000000001110000",
9546 => "0000000001110000",
9547 => "0000000001110000",
9548 => "0000000001110000",
9549 => "0000000001110000",
9550 => "0000000001110000",
9551 => "0000000001110000",
9552 => "0000000001110000",
9553 => "0000000001110000",
9554 => "0000000001110000",
9555 => "0000000001110000",
9556 => "0000000001110000",
9557 => "0000000001110000",
9558 => "0000000001110001",
9559 => "0000000001110001",
9560 => "0000000001110001",
9561 => "0000000001110001",
9562 => "0000000001110001",
9563 => "0000000001110001",
9564 => "0000000001110001",
9565 => "0000000001110001",
9566 => "0000000001110001",
9567 => "0000000001110001",
9568 => "0000000001110001",
9569 => "0000000001110001",
9570 => "0000000001110001",
9571 => "0000000001110001",
9572 => "0000000001110001",
9573 => "0000000001110001",
9574 => "0000000001110001",
9575 => "0000000001110001",
9576 => "0000000001110001",
9577 => "0000000001110001",
9578 => "0000000001110001",
9579 => "0000000001110001",
9580 => "0000000001110001",
9581 => "0000000001110001",
9582 => "0000000001110001",
9583 => "0000000001110001",
9584 => "0000000001110001",
9585 => "0000000001110001",
9586 => "0000000001110001",
9587 => "0000000001110001",
9588 => "0000000001110001",
9589 => "0000000001110001",
9590 => "0000000001110001",
9591 => "0000000001110001",
9592 => "0000000001110001",
9593 => "0000000001110001",
9594 => "0000000001110010",
9595 => "0000000001110010",
9596 => "0000000001110010",
9597 => "0000000001110010",
9598 => "0000000001110010",
9599 => "0000000001110010",
9600 => "0000000001110010",
9601 => "0000000001110010",
9602 => "0000000001110010",
9603 => "0000000001110010",
9604 => "0000000001110010",
9605 => "0000000001110010",
9606 => "0000000001110010",
9607 => "0000000001110010",
9608 => "0000000001110010",
9609 => "0000000001110010",
9610 => "0000000001110010",
9611 => "0000000001110010",
9612 => "0000000001110010",
9613 => "0000000001110010",
9614 => "0000000001110010",
9615 => "0000000001110010",
9616 => "0000000001110010",
9617 => "0000000001110010",
9618 => "0000000001110010",
9619 => "0000000001110010",
9620 => "0000000001110010",
9621 => "0000000001110010",
9622 => "0000000001110010",
9623 => "0000000001110010",
9624 => "0000000001110010",
9625 => "0000000001110010",
9626 => "0000000001110010",
9627 => "0000000001110010",
9628 => "0000000001110010",
9629 => "0000000001110010",
9630 => "0000000001110011",
9631 => "0000000001110011",
9632 => "0000000001110011",
9633 => "0000000001110011",
9634 => "0000000001110011",
9635 => "0000000001110011",
9636 => "0000000001110011",
9637 => "0000000001110011",
9638 => "0000000001110011",
9639 => "0000000001110011",
9640 => "0000000001110011",
9641 => "0000000001110011",
9642 => "0000000001110011",
9643 => "0000000001110011",
9644 => "0000000001110011",
9645 => "0000000001110011",
9646 => "0000000001110011",
9647 => "0000000001110011",
9648 => "0000000001110011",
9649 => "0000000001110011",
9650 => "0000000001110011",
9651 => "0000000001110011",
9652 => "0000000001110011",
9653 => "0000000001110011",
9654 => "0000000001110011",
9655 => "0000000001110011",
9656 => "0000000001110011",
9657 => "0000000001110011",
9658 => "0000000001110011",
9659 => "0000000001110011",
9660 => "0000000001110011",
9661 => "0000000001110011",
9662 => "0000000001110011",
9663 => "0000000001110011",
9664 => "0000000001110011",
9665 => "0000000001110011",
9666 => "0000000001110100",
9667 => "0000000001110100",
9668 => "0000000001110100",
9669 => "0000000001110100",
9670 => "0000000001110100",
9671 => "0000000001110100",
9672 => "0000000001110100",
9673 => "0000000001110100",
9674 => "0000000001110100",
9675 => "0000000001110100",
9676 => "0000000001110100",
9677 => "0000000001110100",
9678 => "0000000001110100",
9679 => "0000000001110100",
9680 => "0000000001110100",
9681 => "0000000001110100",
9682 => "0000000001110100",
9683 => "0000000001110100",
9684 => "0000000001110100",
9685 => "0000000001110100",
9686 => "0000000001110100",
9687 => "0000000001110100",
9688 => "0000000001110100",
9689 => "0000000001110100",
9690 => "0000000001110100",
9691 => "0000000001110100",
9692 => "0000000001110100",
9693 => "0000000001110100",
9694 => "0000000001110100",
9695 => "0000000001110100",
9696 => "0000000001110100",
9697 => "0000000001110100",
9698 => "0000000001110100",
9699 => "0000000001110100",
9700 => "0000000001110100",
9701 => "0000000001110101",
9702 => "0000000001110101",
9703 => "0000000001110101",
9704 => "0000000001110101",
9705 => "0000000001110101",
9706 => "0000000001110101",
9707 => "0000000001110101",
9708 => "0000000001110101",
9709 => "0000000001110101",
9710 => "0000000001110101",
9711 => "0000000001110101",
9712 => "0000000001110101",
9713 => "0000000001110101",
9714 => "0000000001110101",
9715 => "0000000001110101",
9716 => "0000000001110101",
9717 => "0000000001110101",
9718 => "0000000001110101",
9719 => "0000000001110101",
9720 => "0000000001110101",
9721 => "0000000001110101",
9722 => "0000000001110101",
9723 => "0000000001110101",
9724 => "0000000001110101",
9725 => "0000000001110101",
9726 => "0000000001110101",
9727 => "0000000001110101",
9728 => "0000000001110101",
9729 => "0000000001110101",
9730 => "0000000001110101",
9731 => "0000000001110101",
9732 => "0000000001110101",
9733 => "0000000001110101",
9734 => "0000000001110101",
9735 => "0000000001110101",
9736 => "0000000001110110",
9737 => "0000000001110110",
9738 => "0000000001110110",
9739 => "0000000001110110",
9740 => "0000000001110110",
9741 => "0000000001110110",
9742 => "0000000001110110",
9743 => "0000000001110110",
9744 => "0000000001110110",
9745 => "0000000001110110",
9746 => "0000000001110110",
9747 => "0000000001110110",
9748 => "0000000001110110",
9749 => "0000000001110110",
9750 => "0000000001110110",
9751 => "0000000001110110",
9752 => "0000000001110110",
9753 => "0000000001110110",
9754 => "0000000001110110",
9755 => "0000000001110110",
9756 => "0000000001110110",
9757 => "0000000001110110",
9758 => "0000000001110110",
9759 => "0000000001110110",
9760 => "0000000001110110",
9761 => "0000000001110110",
9762 => "0000000001110110",
9763 => "0000000001110110",
9764 => "0000000001110110",
9765 => "0000000001110110",
9766 => "0000000001110110",
9767 => "0000000001110110",
9768 => "0000000001110110",
9769 => "0000000001110110",
9770 => "0000000001110110",
9771 => "0000000001110111",
9772 => "0000000001110111",
9773 => "0000000001110111",
9774 => "0000000001110111",
9775 => "0000000001110111",
9776 => "0000000001110111",
9777 => "0000000001110111",
9778 => "0000000001110111",
9779 => "0000000001110111",
9780 => "0000000001110111",
9781 => "0000000001110111",
9782 => "0000000001110111",
9783 => "0000000001110111",
9784 => "0000000001110111",
9785 => "0000000001110111",
9786 => "0000000001110111",
9787 => "0000000001110111",
9788 => "0000000001110111",
9789 => "0000000001110111",
9790 => "0000000001110111",
9791 => "0000000001110111",
9792 => "0000000001110111",
9793 => "0000000001110111",
9794 => "0000000001110111",
9795 => "0000000001110111",
9796 => "0000000001110111",
9797 => "0000000001110111",
9798 => "0000000001110111",
9799 => "0000000001110111",
9800 => "0000000001110111",
9801 => "0000000001110111",
9802 => "0000000001110111",
9803 => "0000000001110111",
9804 => "0000000001110111",
9805 => "0000000001111000",
9806 => "0000000001111000",
9807 => "0000000001111000",
9808 => "0000000001111000",
9809 => "0000000001111000",
9810 => "0000000001111000",
9811 => "0000000001111000",
9812 => "0000000001111000",
9813 => "0000000001111000",
9814 => "0000000001111000",
9815 => "0000000001111000",
9816 => "0000000001111000",
9817 => "0000000001111000",
9818 => "0000000001111000",
9819 => "0000000001111000",
9820 => "0000000001111000",
9821 => "0000000001111000",
9822 => "0000000001111000",
9823 => "0000000001111000",
9824 => "0000000001111000",
9825 => "0000000001111000",
9826 => "0000000001111000",
9827 => "0000000001111000",
9828 => "0000000001111000",
9829 => "0000000001111000",
9830 => "0000000001111000",
9831 => "0000000001111000",
9832 => "0000000001111000",
9833 => "0000000001111000",
9834 => "0000000001111000",
9835 => "0000000001111000",
9836 => "0000000001111000",
9837 => "0000000001111000",
9838 => "0000000001111000",
9839 => "0000000001111001",
9840 => "0000000001111001",
9841 => "0000000001111001",
9842 => "0000000001111001",
9843 => "0000000001111001",
9844 => "0000000001111001",
9845 => "0000000001111001",
9846 => "0000000001111001",
9847 => "0000000001111001",
9848 => "0000000001111001",
9849 => "0000000001111001",
9850 => "0000000001111001",
9851 => "0000000001111001",
9852 => "0000000001111001",
9853 => "0000000001111001",
9854 => "0000000001111001",
9855 => "0000000001111001",
9856 => "0000000001111001",
9857 => "0000000001111001",
9858 => "0000000001111001",
9859 => "0000000001111001",
9860 => "0000000001111001",
9861 => "0000000001111001",
9862 => "0000000001111001",
9863 => "0000000001111001",
9864 => "0000000001111001",
9865 => "0000000001111001",
9866 => "0000000001111001",
9867 => "0000000001111001",
9868 => "0000000001111001",
9869 => "0000000001111001",
9870 => "0000000001111001",
9871 => "0000000001111001",
9872 => "0000000001111001",
9873 => "0000000001111010",
9874 => "0000000001111010",
9875 => "0000000001111010",
9876 => "0000000001111010",
9877 => "0000000001111010",
9878 => "0000000001111010",
9879 => "0000000001111010",
9880 => "0000000001111010",
9881 => "0000000001111010",
9882 => "0000000001111010",
9883 => "0000000001111010",
9884 => "0000000001111010",
9885 => "0000000001111010",
9886 => "0000000001111010",
9887 => "0000000001111010",
9888 => "0000000001111010",
9889 => "0000000001111010",
9890 => "0000000001111010",
9891 => "0000000001111010",
9892 => "0000000001111010",
9893 => "0000000001111010",
9894 => "0000000001111010",
9895 => "0000000001111010",
9896 => "0000000001111010",
9897 => "0000000001111010",
9898 => "0000000001111010",
9899 => "0000000001111010",
9900 => "0000000001111010",
9901 => "0000000001111010",
9902 => "0000000001111010",
9903 => "0000000001111010",
9904 => "0000000001111010",
9905 => "0000000001111010",
9906 => "0000000001111011",
9907 => "0000000001111011",
9908 => "0000000001111011",
9909 => "0000000001111011",
9910 => "0000000001111011",
9911 => "0000000001111011",
9912 => "0000000001111011",
9913 => "0000000001111011",
9914 => "0000000001111011",
9915 => "0000000001111011",
9916 => "0000000001111011",
9917 => "0000000001111011",
9918 => "0000000001111011",
9919 => "0000000001111011",
9920 => "0000000001111011",
9921 => "0000000001111011",
9922 => "0000000001111011",
9923 => "0000000001111011",
9924 => "0000000001111011",
9925 => "0000000001111011",
9926 => "0000000001111011",
9927 => "0000000001111011",
9928 => "0000000001111011",
9929 => "0000000001111011",
9930 => "0000000001111011",
9931 => "0000000001111011",
9932 => "0000000001111011",
9933 => "0000000001111011",
9934 => "0000000001111011",
9935 => "0000000001111011",
9936 => "0000000001111011",
9937 => "0000000001111011",
9938 => "0000000001111011",
9939 => "0000000001111011",
9940 => "0000000001111100",
9941 => "0000000001111100",
9942 => "0000000001111100",
9943 => "0000000001111100",
9944 => "0000000001111100",
9945 => "0000000001111100",
9946 => "0000000001111100",
9947 => "0000000001111100",
9948 => "0000000001111100",
9949 => "0000000001111100",
9950 => "0000000001111100",
9951 => "0000000001111100",
9952 => "0000000001111100",
9953 => "0000000001111100",
9954 => "0000000001111100",
9955 => "0000000001111100",
9956 => "0000000001111100",
9957 => "0000000001111100",
9958 => "0000000001111100",
9959 => "0000000001111100",
9960 => "0000000001111100",
9961 => "0000000001111100",
9962 => "0000000001111100",
9963 => "0000000001111100",
9964 => "0000000001111100",
9965 => "0000000001111100",
9966 => "0000000001111100",
9967 => "0000000001111100",
9968 => "0000000001111100",
9969 => "0000000001111100",
9970 => "0000000001111100",
9971 => "0000000001111100",
9972 => "0000000001111100",
9973 => "0000000001111101",
9974 => "0000000001111101",
9975 => "0000000001111101",
9976 => "0000000001111101",
9977 => "0000000001111101",
9978 => "0000000001111101",
9979 => "0000000001111101",
9980 => "0000000001111101",
9981 => "0000000001111101",
9982 => "0000000001111101",
9983 => "0000000001111101",
9984 => "0000000001111101",
9985 => "0000000001111101",
9986 => "0000000001111101",
9987 => "0000000001111101",
9988 => "0000000001111101",
9989 => "0000000001111101",
9990 => "0000000001111101",
9991 => "0000000001111101",
9992 => "0000000001111101",
9993 => "0000000001111101",
9994 => "0000000001111101",
9995 => "0000000001111101",
9996 => "0000000001111101",
9997 => "0000000001111101",
9998 => "0000000001111101",
9999 => "0000000001111101",
10000 => "0000000001111101",
10001 => "0000000001111101",
10002 => "0000000001111101",
10003 => "0000000001111101",
10004 => "0000000001111101",
10005 => "0000000001111101",
10006 => "0000000001111110",
10007 => "0000000001111110",
10008 => "0000000001111110",
10009 => "0000000001111110",
10010 => "0000000001111110",
10011 => "0000000001111110",
10012 => "0000000001111110",
10013 => "0000000001111110",
10014 => "0000000001111110",
10015 => "0000000001111110",
10016 => "0000000001111110",
10017 => "0000000001111110",
10018 => "0000000001111110",
10019 => "0000000001111110",
10020 => "0000000001111110",
10021 => "0000000001111110",
10022 => "0000000001111110",
10023 => "0000000001111110",
10024 => "0000000001111110",
10025 => "0000000001111110",
10026 => "0000000001111110",
10027 => "0000000001111110",
10028 => "0000000001111110",
10029 => "0000000001111110",
10030 => "0000000001111110",
10031 => "0000000001111110",
10032 => "0000000001111110",
10033 => "0000000001111110",
10034 => "0000000001111110",
10035 => "0000000001111110",
10036 => "0000000001111110",
10037 => "0000000001111110",
10038 => "0000000001111111",
10039 => "0000000001111111",
10040 => "0000000001111111",
10041 => "0000000001111111",
10042 => "0000000001111111",
10043 => "0000000001111111",
10044 => "0000000001111111",
10045 => "0000000001111111",
10046 => "0000000001111111",
10047 => "0000000001111111",
10048 => "0000000001111111",
10049 => "0000000001111111",
10050 => "0000000001111111",
10051 => "0000000001111111",
10052 => "0000000001111111",
10053 => "0000000001111111",
10054 => "0000000001111111",
10055 => "0000000001111111",
10056 => "0000000001111111",
10057 => "0000000001111111",
10058 => "0000000001111111",
10059 => "0000000001111111",
10060 => "0000000001111111",
10061 => "0000000001111111",
10062 => "0000000001111111",
10063 => "0000000001111111",
10064 => "0000000001111111",
10065 => "0000000001111111",
10066 => "0000000001111111",
10067 => "0000000001111111",
10068 => "0000000001111111",
10069 => "0000000001111111",
10070 => "0000000010000000",
10071 => "0000000010000000",
10072 => "0000000010000000",
10073 => "0000000010000000",
10074 => "0000000010000000",
10075 => "0000000010000000",
10076 => "0000000010000000",
10077 => "0000000010000000",
10078 => "0000000010000000",
10079 => "0000000010000000",
10080 => "0000000010000000",
10081 => "0000000010000000",
10082 => "0000000010000000",
10083 => "0000000010000000",
10084 => "0000000010000000",
10085 => "0000000010000000",
10086 => "0000000010000000",
10087 => "0000000010000000",
10088 => "0000000010000000",
10089 => "0000000010000000",
10090 => "0000000010000000",
10091 => "0000000010000000",
10092 => "0000000010000000",
10093 => "0000000010000000",
10094 => "0000000010000000",
10095 => "0000000010000000",
10096 => "0000000010000000",
10097 => "0000000010000000",
10098 => "0000000010000000",
10099 => "0000000010000000",
10100 => "0000000010000000",
10101 => "0000000010000001",
10102 => "0000000010000001",
10103 => "0000000010000001",
10104 => "0000000010000001",
10105 => "0000000010000001",
10106 => "0000000010000001",
10107 => "0000000010000001",
10108 => "0000000010000001",
10109 => "0000000010000001",
10110 => "0000000010000001",
10111 => "0000000010000001",
10112 => "0000000010000001",
10113 => "0000000010000001",
10114 => "0000000010000001",
10115 => "0000000010000001",
10116 => "0000000010000001",
10117 => "0000000010000001",
10118 => "0000000010000001",
10119 => "0000000010000001",
10120 => "0000000010000001",
10121 => "0000000010000001",
10122 => "0000000010000001",
10123 => "0000000010000001",
10124 => "0000000010000001",
10125 => "0000000010000001",
10126 => "0000000010000001",
10127 => "0000000010000001",
10128 => "0000000010000001",
10129 => "0000000010000001",
10130 => "0000000010000001",
10131 => "0000000010000001",
10132 => "0000000010000001",
10133 => "0000000010000010",
10134 => "0000000010000010",
10135 => "0000000010000010",
10136 => "0000000010000010",
10137 => "0000000010000010",
10138 => "0000000010000010",
10139 => "0000000010000010",
10140 => "0000000010000010",
10141 => "0000000010000010",
10142 => "0000000010000010",
10143 => "0000000010000010",
10144 => "0000000010000010",
10145 => "0000000010000010",
10146 => "0000000010000010",
10147 => "0000000010000010",
10148 => "0000000010000010",
10149 => "0000000010000010",
10150 => "0000000010000010",
10151 => "0000000010000010",
10152 => "0000000010000010",
10153 => "0000000010000010",
10154 => "0000000010000010",
10155 => "0000000010000010",
10156 => "0000000010000010",
10157 => "0000000010000010",
10158 => "0000000010000010",
10159 => "0000000010000010",
10160 => "0000000010000010",
10161 => "0000000010000010",
10162 => "0000000010000010",
10163 => "0000000010000010",
10164 => "0000000010000010",
10165 => "0000000010000011",
10166 => "0000000010000011",
10167 => "0000000010000011",
10168 => "0000000010000011",
10169 => "0000000010000011",
10170 => "0000000010000011",
10171 => "0000000010000011",
10172 => "0000000010000011",
10173 => "0000000010000011",
10174 => "0000000010000011",
10175 => "0000000010000011",
10176 => "0000000010000011",
10177 => "0000000010000011",
10178 => "0000000010000011",
10179 => "0000000010000011",
10180 => "0000000010000011",
10181 => "0000000010000011",
10182 => "0000000010000011",
10183 => "0000000010000011",
10184 => "0000000010000011",
10185 => "0000000010000011",
10186 => "0000000010000011",
10187 => "0000000010000011",
10188 => "0000000010000011",
10189 => "0000000010000011",
10190 => "0000000010000011",
10191 => "0000000010000011",
10192 => "0000000010000011",
10193 => "0000000010000011",
10194 => "0000000010000011",
10195 => "0000000010000011",
10196 => "0000000010000100",
10197 => "0000000010000100",
10198 => "0000000010000100",
10199 => "0000000010000100",
10200 => "0000000010000100",
10201 => "0000000010000100",
10202 => "0000000010000100",
10203 => "0000000010000100",
10204 => "0000000010000100",
10205 => "0000000010000100",
10206 => "0000000010000100",
10207 => "0000000010000100",
10208 => "0000000010000100",
10209 => "0000000010000100",
10210 => "0000000010000100",
10211 => "0000000010000100",
10212 => "0000000010000100",
10213 => "0000000010000100",
10214 => "0000000010000100",
10215 => "0000000010000100",
10216 => "0000000010000100",
10217 => "0000000010000100",
10218 => "0000000010000100",
10219 => "0000000010000100",
10220 => "0000000010000100",
10221 => "0000000010000100",
10222 => "0000000010000100",
10223 => "0000000010000100",
10224 => "0000000010000100",
10225 => "0000000010000100",
10226 => "0000000010000100",
10227 => "0000000010000101",
10228 => "0000000010000101",
10229 => "0000000010000101",
10230 => "0000000010000101",
10231 => "0000000010000101",
10232 => "0000000010000101",
10233 => "0000000010000101",
10234 => "0000000010000101",
10235 => "0000000010000101",
10236 => "0000000010000101",
10237 => "0000000010000101",
10238 => "0000000010000101",
10239 => "0000000010000101",
10240 => "0000000010000101",
10241 => "0000000010000101",
10242 => "0000000010000101",
10243 => "0000000010000101",
10244 => "0000000010000101",
10245 => "0000000010000101",
10246 => "0000000010000101",
10247 => "0000000010000101",
10248 => "0000000010000101",
10249 => "0000000010000101",
10250 => "0000000010000101",
10251 => "0000000010000101",
10252 => "0000000010000101",
10253 => "0000000010000101",
10254 => "0000000010000101",
10255 => "0000000010000101",
10256 => "0000000010000101",
10257 => "0000000010000101",
10258 => "0000000010000110",
10259 => "0000000010000110",
10260 => "0000000010000110",
10261 => "0000000010000110",
10262 => "0000000010000110",
10263 => "0000000010000110",
10264 => "0000000010000110",
10265 => "0000000010000110",
10266 => "0000000010000110",
10267 => "0000000010000110",
10268 => "0000000010000110",
10269 => "0000000010000110",
10270 => "0000000010000110",
10271 => "0000000010000110",
10272 => "0000000010000110",
10273 => "0000000010000110",
10274 => "0000000010000110",
10275 => "0000000010000110",
10276 => "0000000010000110",
10277 => "0000000010000110",
10278 => "0000000010000110",
10279 => "0000000010000110",
10280 => "0000000010000110",
10281 => "0000000010000110",
10282 => "0000000010000110",
10283 => "0000000010000110",
10284 => "0000000010000110",
10285 => "0000000010000110",
10286 => "0000000010000110",
10287 => "0000000010000110",
10288 => "0000000010000111",
10289 => "0000000010000111",
10290 => "0000000010000111",
10291 => "0000000010000111",
10292 => "0000000010000111",
10293 => "0000000010000111",
10294 => "0000000010000111",
10295 => "0000000010000111",
10296 => "0000000010000111",
10297 => "0000000010000111",
10298 => "0000000010000111",
10299 => "0000000010000111",
10300 => "0000000010000111",
10301 => "0000000010000111",
10302 => "0000000010000111",
10303 => "0000000010000111",
10304 => "0000000010000111",
10305 => "0000000010000111",
10306 => "0000000010000111",
10307 => "0000000010000111",
10308 => "0000000010000111",
10309 => "0000000010000111",
10310 => "0000000010000111",
10311 => "0000000010000111",
10312 => "0000000010000111",
10313 => "0000000010000111",
10314 => "0000000010000111",
10315 => "0000000010000111",
10316 => "0000000010000111",
10317 => "0000000010000111",
10318 => "0000000010000111",
10319 => "0000000010001000",
10320 => "0000000010001000",
10321 => "0000000010001000",
10322 => "0000000010001000",
10323 => "0000000010001000",
10324 => "0000000010001000",
10325 => "0000000010001000",
10326 => "0000000010001000",
10327 => "0000000010001000",
10328 => "0000000010001000",
10329 => "0000000010001000",
10330 => "0000000010001000",
10331 => "0000000010001000",
10332 => "0000000010001000",
10333 => "0000000010001000",
10334 => "0000000010001000",
10335 => "0000000010001000",
10336 => "0000000010001000",
10337 => "0000000010001000",
10338 => "0000000010001000",
10339 => "0000000010001000",
10340 => "0000000010001000",
10341 => "0000000010001000",
10342 => "0000000010001000",
10343 => "0000000010001000",
10344 => "0000000010001000",
10345 => "0000000010001000",
10346 => "0000000010001000",
10347 => "0000000010001000",
10348 => "0000000010001000",
10349 => "0000000010001001",
10350 => "0000000010001001",
10351 => "0000000010001001",
10352 => "0000000010001001",
10353 => "0000000010001001",
10354 => "0000000010001001",
10355 => "0000000010001001",
10356 => "0000000010001001",
10357 => "0000000010001001",
10358 => "0000000010001001",
10359 => "0000000010001001",
10360 => "0000000010001001",
10361 => "0000000010001001",
10362 => "0000000010001001",
10363 => "0000000010001001",
10364 => "0000000010001001",
10365 => "0000000010001001",
10366 => "0000000010001001",
10367 => "0000000010001001",
10368 => "0000000010001001",
10369 => "0000000010001001",
10370 => "0000000010001001",
10371 => "0000000010001001",
10372 => "0000000010001001",
10373 => "0000000010001001",
10374 => "0000000010001001",
10375 => "0000000010001001",
10376 => "0000000010001001",
10377 => "0000000010001001",
10378 => "0000000010001001",
10379 => "0000000010001010",
10380 => "0000000010001010",
10381 => "0000000010001010",
10382 => "0000000010001010",
10383 => "0000000010001010",
10384 => "0000000010001010",
10385 => "0000000010001010",
10386 => "0000000010001010",
10387 => "0000000010001010",
10388 => "0000000010001010",
10389 => "0000000010001010",
10390 => "0000000010001010",
10391 => "0000000010001010",
10392 => "0000000010001010",
10393 => "0000000010001010",
10394 => "0000000010001010",
10395 => "0000000010001010",
10396 => "0000000010001010",
10397 => "0000000010001010",
10398 => "0000000010001010",
10399 => "0000000010001010",
10400 => "0000000010001010",
10401 => "0000000010001010",
10402 => "0000000010001010",
10403 => "0000000010001010",
10404 => "0000000010001010",
10405 => "0000000010001010",
10406 => "0000000010001010",
10407 => "0000000010001010",
10408 => "0000000010001010",
10409 => "0000000010001011",
10410 => "0000000010001011",
10411 => "0000000010001011",
10412 => "0000000010001011",
10413 => "0000000010001011",
10414 => "0000000010001011",
10415 => "0000000010001011",
10416 => "0000000010001011",
10417 => "0000000010001011",
10418 => "0000000010001011",
10419 => "0000000010001011",
10420 => "0000000010001011",
10421 => "0000000010001011",
10422 => "0000000010001011",
10423 => "0000000010001011",
10424 => "0000000010001011",
10425 => "0000000010001011",
10426 => "0000000010001011",
10427 => "0000000010001011",
10428 => "0000000010001011",
10429 => "0000000010001011",
10430 => "0000000010001011",
10431 => "0000000010001011",
10432 => "0000000010001011",
10433 => "0000000010001011",
10434 => "0000000010001011",
10435 => "0000000010001011",
10436 => "0000000010001011",
10437 => "0000000010001011",
10438 => "0000000010001100",
10439 => "0000000010001100",
10440 => "0000000010001100",
10441 => "0000000010001100",
10442 => "0000000010001100",
10443 => "0000000010001100",
10444 => "0000000010001100",
10445 => "0000000010001100",
10446 => "0000000010001100",
10447 => "0000000010001100",
10448 => "0000000010001100",
10449 => "0000000010001100",
10450 => "0000000010001100",
10451 => "0000000010001100",
10452 => "0000000010001100",
10453 => "0000000010001100",
10454 => "0000000010001100",
10455 => "0000000010001100",
10456 => "0000000010001100",
10457 => "0000000010001100",
10458 => "0000000010001100",
10459 => "0000000010001100",
10460 => "0000000010001100",
10461 => "0000000010001100",
10462 => "0000000010001100",
10463 => "0000000010001100",
10464 => "0000000010001100",
10465 => "0000000010001100",
10466 => "0000000010001100",
10467 => "0000000010001101",
10468 => "0000000010001101",
10469 => "0000000010001101",
10470 => "0000000010001101",
10471 => "0000000010001101",
10472 => "0000000010001101",
10473 => "0000000010001101",
10474 => "0000000010001101",
10475 => "0000000010001101",
10476 => "0000000010001101",
10477 => "0000000010001101",
10478 => "0000000010001101",
10479 => "0000000010001101",
10480 => "0000000010001101",
10481 => "0000000010001101",
10482 => "0000000010001101",
10483 => "0000000010001101",
10484 => "0000000010001101",
10485 => "0000000010001101",
10486 => "0000000010001101",
10487 => "0000000010001101",
10488 => "0000000010001101",
10489 => "0000000010001101",
10490 => "0000000010001101",
10491 => "0000000010001101",
10492 => "0000000010001101",
10493 => "0000000010001101",
10494 => "0000000010001101",
10495 => "0000000010001101",
10496 => "0000000010001110",
10497 => "0000000010001110",
10498 => "0000000010001110",
10499 => "0000000010001110",
10500 => "0000000010001110",
10501 => "0000000010001110",
10502 => "0000000010001110",
10503 => "0000000010001110",
10504 => "0000000010001110",
10505 => "0000000010001110",
10506 => "0000000010001110",
10507 => "0000000010001110",
10508 => "0000000010001110",
10509 => "0000000010001110",
10510 => "0000000010001110",
10511 => "0000000010001110",
10512 => "0000000010001110",
10513 => "0000000010001110",
10514 => "0000000010001110",
10515 => "0000000010001110",
10516 => "0000000010001110",
10517 => "0000000010001110",
10518 => "0000000010001110",
10519 => "0000000010001110",
10520 => "0000000010001110",
10521 => "0000000010001110",
10522 => "0000000010001110",
10523 => "0000000010001110",
10524 => "0000000010001110",
10525 => "0000000010001111",
10526 => "0000000010001111",
10527 => "0000000010001111",
10528 => "0000000010001111",
10529 => "0000000010001111",
10530 => "0000000010001111",
10531 => "0000000010001111",
10532 => "0000000010001111",
10533 => "0000000010001111",
10534 => "0000000010001111",
10535 => "0000000010001111",
10536 => "0000000010001111",
10537 => "0000000010001111",
10538 => "0000000010001111",
10539 => "0000000010001111",
10540 => "0000000010001111",
10541 => "0000000010001111",
10542 => "0000000010001111",
10543 => "0000000010001111",
10544 => "0000000010001111",
10545 => "0000000010001111",
10546 => "0000000010001111",
10547 => "0000000010001111",
10548 => "0000000010001111",
10549 => "0000000010001111",
10550 => "0000000010001111",
10551 => "0000000010001111",
10552 => "0000000010001111",
10553 => "0000000010001111",
10554 => "0000000010010000",
10555 => "0000000010010000",
10556 => "0000000010010000",
10557 => "0000000010010000",
10558 => "0000000010010000",
10559 => "0000000010010000",
10560 => "0000000010010000",
10561 => "0000000010010000",
10562 => "0000000010010000",
10563 => "0000000010010000",
10564 => "0000000010010000",
10565 => "0000000010010000",
10566 => "0000000010010000",
10567 => "0000000010010000",
10568 => "0000000010010000",
10569 => "0000000010010000",
10570 => "0000000010010000",
10571 => "0000000010010000",
10572 => "0000000010010000",
10573 => "0000000010010000",
10574 => "0000000010010000",
10575 => "0000000010010000",
10576 => "0000000010010000",
10577 => "0000000010010000",
10578 => "0000000010010000",
10579 => "0000000010010000",
10580 => "0000000010010000",
10581 => "0000000010010000",
10582 => "0000000010010001",
10583 => "0000000010010001",
10584 => "0000000010010001",
10585 => "0000000010010001",
10586 => "0000000010010001",
10587 => "0000000010010001",
10588 => "0000000010010001",
10589 => "0000000010010001",
10590 => "0000000010010001",
10591 => "0000000010010001",
10592 => "0000000010010001",
10593 => "0000000010010001",
10594 => "0000000010010001",
10595 => "0000000010010001",
10596 => "0000000010010001",
10597 => "0000000010010001",
10598 => "0000000010010001",
10599 => "0000000010010001",
10600 => "0000000010010001",
10601 => "0000000010010001",
10602 => "0000000010010001",
10603 => "0000000010010001",
10604 => "0000000010010001",
10605 => "0000000010010001",
10606 => "0000000010010001",
10607 => "0000000010010001",
10608 => "0000000010010001",
10609 => "0000000010010001",
10610 => "0000000010010001",
10611 => "0000000010010010",
10612 => "0000000010010010",
10613 => "0000000010010010",
10614 => "0000000010010010",
10615 => "0000000010010010",
10616 => "0000000010010010",
10617 => "0000000010010010",
10618 => "0000000010010010",
10619 => "0000000010010010",
10620 => "0000000010010010",
10621 => "0000000010010010",
10622 => "0000000010010010",
10623 => "0000000010010010",
10624 => "0000000010010010",
10625 => "0000000010010010",
10626 => "0000000010010010",
10627 => "0000000010010010",
10628 => "0000000010010010",
10629 => "0000000010010010",
10630 => "0000000010010010",
10631 => "0000000010010010",
10632 => "0000000010010010",
10633 => "0000000010010010",
10634 => "0000000010010010",
10635 => "0000000010010010",
10636 => "0000000010010010",
10637 => "0000000010010010",
10638 => "0000000010010010",
10639 => "0000000010010011",
10640 => "0000000010010011",
10641 => "0000000010010011",
10642 => "0000000010010011",
10643 => "0000000010010011",
10644 => "0000000010010011",
10645 => "0000000010010011",
10646 => "0000000010010011",
10647 => "0000000010010011",
10648 => "0000000010010011",
10649 => "0000000010010011",
10650 => "0000000010010011",
10651 => "0000000010010011",
10652 => "0000000010010011",
10653 => "0000000010010011",
10654 => "0000000010010011",
10655 => "0000000010010011",
10656 => "0000000010010011",
10657 => "0000000010010011",
10658 => "0000000010010011",
10659 => "0000000010010011",
10660 => "0000000010010011",
10661 => "0000000010010011",
10662 => "0000000010010011",
10663 => "0000000010010011",
10664 => "0000000010010011",
10665 => "0000000010010011",
10666 => "0000000010010011",
10667 => "0000000010010100",
10668 => "0000000010010100",
10669 => "0000000010010100",
10670 => "0000000010010100",
10671 => "0000000010010100",
10672 => "0000000010010100",
10673 => "0000000010010100",
10674 => "0000000010010100",
10675 => "0000000010010100",
10676 => "0000000010010100",
10677 => "0000000010010100",
10678 => "0000000010010100",
10679 => "0000000010010100",
10680 => "0000000010010100",
10681 => "0000000010010100",
10682 => "0000000010010100",
10683 => "0000000010010100",
10684 => "0000000010010100",
10685 => "0000000010010100",
10686 => "0000000010010100",
10687 => "0000000010010100",
10688 => "0000000010010100",
10689 => "0000000010010100",
10690 => "0000000010010100",
10691 => "0000000010010100",
10692 => "0000000010010100",
10693 => "0000000010010100",
10694 => "0000000010010101",
10695 => "0000000010010101",
10696 => "0000000010010101",
10697 => "0000000010010101",
10698 => "0000000010010101",
10699 => "0000000010010101",
10700 => "0000000010010101",
10701 => "0000000010010101",
10702 => "0000000010010101",
10703 => "0000000010010101",
10704 => "0000000010010101",
10705 => "0000000010010101",
10706 => "0000000010010101",
10707 => "0000000010010101",
10708 => "0000000010010101",
10709 => "0000000010010101",
10710 => "0000000010010101",
10711 => "0000000010010101",
10712 => "0000000010010101",
10713 => "0000000010010101",
10714 => "0000000010010101",
10715 => "0000000010010101",
10716 => "0000000010010101",
10717 => "0000000010010101",
10718 => "0000000010010101",
10719 => "0000000010010101",
10720 => "0000000010010101",
10721 => "0000000010010101",
10722 => "0000000010010110",
10723 => "0000000010010110",
10724 => "0000000010010110",
10725 => "0000000010010110",
10726 => "0000000010010110",
10727 => "0000000010010110",
10728 => "0000000010010110",
10729 => "0000000010010110",
10730 => "0000000010010110",
10731 => "0000000010010110",
10732 => "0000000010010110",
10733 => "0000000010010110",
10734 => "0000000010010110",
10735 => "0000000010010110",
10736 => "0000000010010110",
10737 => "0000000010010110",
10738 => "0000000010010110",
10739 => "0000000010010110",
10740 => "0000000010010110",
10741 => "0000000010010110",
10742 => "0000000010010110",
10743 => "0000000010010110",
10744 => "0000000010010110",
10745 => "0000000010010110",
10746 => "0000000010010110",
10747 => "0000000010010110",
10748 => "0000000010010110",
10749 => "0000000010010111",
10750 => "0000000010010111",
10751 => "0000000010010111",
10752 => "0000000010010111",
10753 => "0000000010010111",
10754 => "0000000010010111",
10755 => "0000000010010111",
10756 => "0000000010010111",
10757 => "0000000010010111",
10758 => "0000000010010111",
10759 => "0000000010010111",
10760 => "0000000010010111",
10761 => "0000000010010111",
10762 => "0000000010010111",
10763 => "0000000010010111",
10764 => "0000000010010111",
10765 => "0000000010010111",
10766 => "0000000010010111",
10767 => "0000000010010111",
10768 => "0000000010010111",
10769 => "0000000010010111",
10770 => "0000000010010111",
10771 => "0000000010010111",
10772 => "0000000010010111",
10773 => "0000000010010111",
10774 => "0000000010010111",
10775 => "0000000010010111",
10776 => "0000000010010111",
10777 => "0000000010011000",
10778 => "0000000010011000",
10779 => "0000000010011000",
10780 => "0000000010011000",
10781 => "0000000010011000",
10782 => "0000000010011000",
10783 => "0000000010011000",
10784 => "0000000010011000",
10785 => "0000000010011000",
10786 => "0000000010011000",
10787 => "0000000010011000",
10788 => "0000000010011000",
10789 => "0000000010011000",
10790 => "0000000010011000",
10791 => "0000000010011000",
10792 => "0000000010011000",
10793 => "0000000010011000",
10794 => "0000000010011000",
10795 => "0000000010011000",
10796 => "0000000010011000",
10797 => "0000000010011000",
10798 => "0000000010011000",
10799 => "0000000010011000",
10800 => "0000000010011000",
10801 => "0000000010011000",
10802 => "0000000010011000",
10803 => "0000000010011000",
10804 => "0000000010011001",
10805 => "0000000010011001",
10806 => "0000000010011001",
10807 => "0000000010011001",
10808 => "0000000010011001",
10809 => "0000000010011001",
10810 => "0000000010011001",
10811 => "0000000010011001",
10812 => "0000000010011001",
10813 => "0000000010011001",
10814 => "0000000010011001",
10815 => "0000000010011001",
10816 => "0000000010011001",
10817 => "0000000010011001",
10818 => "0000000010011001",
10819 => "0000000010011001",
10820 => "0000000010011001",
10821 => "0000000010011001",
10822 => "0000000010011001",
10823 => "0000000010011001",
10824 => "0000000010011001",
10825 => "0000000010011001",
10826 => "0000000010011001",
10827 => "0000000010011001",
10828 => "0000000010011001",
10829 => "0000000010011001",
10830 => "0000000010011010",
10831 => "0000000010011010",
10832 => "0000000010011010",
10833 => "0000000010011010",
10834 => "0000000010011010",
10835 => "0000000010011010",
10836 => "0000000010011010",
10837 => "0000000010011010",
10838 => "0000000010011010",
10839 => "0000000010011010",
10840 => "0000000010011010",
10841 => "0000000010011010",
10842 => "0000000010011010",
10843 => "0000000010011010",
10844 => "0000000010011010",
10845 => "0000000010011010",
10846 => "0000000010011010",
10847 => "0000000010011010",
10848 => "0000000010011010",
10849 => "0000000010011010",
10850 => "0000000010011010",
10851 => "0000000010011010",
10852 => "0000000010011010",
10853 => "0000000010011010",
10854 => "0000000010011010",
10855 => "0000000010011010",
10856 => "0000000010011010",
10857 => "0000000010011011",
10858 => "0000000010011011",
10859 => "0000000010011011",
10860 => "0000000010011011",
10861 => "0000000010011011",
10862 => "0000000010011011",
10863 => "0000000010011011",
10864 => "0000000010011011",
10865 => "0000000010011011",
10866 => "0000000010011011",
10867 => "0000000010011011",
10868 => "0000000010011011",
10869 => "0000000010011011",
10870 => "0000000010011011",
10871 => "0000000010011011",
10872 => "0000000010011011",
10873 => "0000000010011011",
10874 => "0000000010011011",
10875 => "0000000010011011",
10876 => "0000000010011011",
10877 => "0000000010011011",
10878 => "0000000010011011",
10879 => "0000000010011011",
10880 => "0000000010011011",
10881 => "0000000010011011",
10882 => "0000000010011011",
10883 => "0000000010011100",
10884 => "0000000010011100",
10885 => "0000000010011100",
10886 => "0000000010011100",
10887 => "0000000010011100",
10888 => "0000000010011100",
10889 => "0000000010011100",
10890 => "0000000010011100",
10891 => "0000000010011100",
10892 => "0000000010011100",
10893 => "0000000010011100",
10894 => "0000000010011100",
10895 => "0000000010011100",
10896 => "0000000010011100",
10897 => "0000000010011100",
10898 => "0000000010011100",
10899 => "0000000010011100",
10900 => "0000000010011100",
10901 => "0000000010011100",
10902 => "0000000010011100",
10903 => "0000000010011100",
10904 => "0000000010011100",
10905 => "0000000010011100",
10906 => "0000000010011100",
10907 => "0000000010011100",
10908 => "0000000010011100",
10909 => "0000000010011100",
10910 => "0000000010011101",
10911 => "0000000010011101",
10912 => "0000000010011101",
10913 => "0000000010011101",
10914 => "0000000010011101",
10915 => "0000000010011101",
10916 => "0000000010011101",
10917 => "0000000010011101",
10918 => "0000000010011101",
10919 => "0000000010011101",
10920 => "0000000010011101",
10921 => "0000000010011101",
10922 => "0000000010011101",
10923 => "0000000010011101",
10924 => "0000000010011101",
10925 => "0000000010011101",
10926 => "0000000010011101",
10927 => "0000000010011101",
10928 => "0000000010011101",
10929 => "0000000010011101",
10930 => "0000000010011101",
10931 => "0000000010011101",
10932 => "0000000010011101",
10933 => "0000000010011101",
10934 => "0000000010011101",
10935 => "0000000010011101",
10936 => "0000000010011110",
10937 => "0000000010011110",
10938 => "0000000010011110",
10939 => "0000000010011110",
10940 => "0000000010011110",
10941 => "0000000010011110",
10942 => "0000000010011110",
10943 => "0000000010011110",
10944 => "0000000010011110",
10945 => "0000000010011110",
10946 => "0000000010011110",
10947 => "0000000010011110",
10948 => "0000000010011110",
10949 => "0000000010011110",
10950 => "0000000010011110",
10951 => "0000000010011110",
10952 => "0000000010011110",
10953 => "0000000010011110",
10954 => "0000000010011110",
10955 => "0000000010011110",
10956 => "0000000010011110",
10957 => "0000000010011110",
10958 => "0000000010011110",
10959 => "0000000010011110",
10960 => "0000000010011110",
10961 => "0000000010011110",
10962 => "0000000010011111",
10963 => "0000000010011111",
10964 => "0000000010011111",
10965 => "0000000010011111",
10966 => "0000000010011111",
10967 => "0000000010011111",
10968 => "0000000010011111",
10969 => "0000000010011111",
10970 => "0000000010011111",
10971 => "0000000010011111",
10972 => "0000000010011111",
10973 => "0000000010011111",
10974 => "0000000010011111",
10975 => "0000000010011111",
10976 => "0000000010011111",
10977 => "0000000010011111",
10978 => "0000000010011111",
10979 => "0000000010011111",
10980 => "0000000010011111",
10981 => "0000000010011111",
10982 => "0000000010011111",
10983 => "0000000010011111",
10984 => "0000000010011111",
10985 => "0000000010011111",
10986 => "0000000010011111",
10987 => "0000000010011111",
10988 => "0000000010100000",
10989 => "0000000010100000",
10990 => "0000000010100000",
10991 => "0000000010100000",
10992 => "0000000010100000",
10993 => "0000000010100000",
10994 => "0000000010100000",
10995 => "0000000010100000",
10996 => "0000000010100000",
10997 => "0000000010100000",
10998 => "0000000010100000",
10999 => "0000000010100000",
11000 => "0000000010100000",
11001 => "0000000010100000",
11002 => "0000000010100000",
11003 => "0000000010100000",
11004 => "0000000010100000",
11005 => "0000000010100000",
11006 => "0000000010100000",
11007 => "0000000010100000",
11008 => "0000000010100000",
11009 => "0000000010100000",
11010 => "0000000010100000",
11011 => "0000000010100000",
11012 => "0000000010100000",
11013 => "0000000010100001",
11014 => "0000000010100001",
11015 => "0000000010100001",
11016 => "0000000010100001",
11017 => "0000000010100001",
11018 => "0000000010100001",
11019 => "0000000010100001",
11020 => "0000000010100001",
11021 => "0000000010100001",
11022 => "0000000010100001",
11023 => "0000000010100001",
11024 => "0000000010100001",
11025 => "0000000010100001",
11026 => "0000000010100001",
11027 => "0000000010100001",
11028 => "0000000010100001",
11029 => "0000000010100001",
11030 => "0000000010100001",
11031 => "0000000010100001",
11032 => "0000000010100001",
11033 => "0000000010100001",
11034 => "0000000010100001",
11035 => "0000000010100001",
11036 => "0000000010100001",
11037 => "0000000010100001",
11038 => "0000000010100001",
11039 => "0000000010100010",
11040 => "0000000010100010",
11041 => "0000000010100010",
11042 => "0000000010100010",
11043 => "0000000010100010",
11044 => "0000000010100010",
11045 => "0000000010100010",
11046 => "0000000010100010",
11047 => "0000000010100010",
11048 => "0000000010100010",
11049 => "0000000010100010",
11050 => "0000000010100010",
11051 => "0000000010100010",
11052 => "0000000010100010",
11053 => "0000000010100010",
11054 => "0000000010100010",
11055 => "0000000010100010",
11056 => "0000000010100010",
11057 => "0000000010100010",
11058 => "0000000010100010",
11059 => "0000000010100010",
11060 => "0000000010100010",
11061 => "0000000010100010",
11062 => "0000000010100010",
11063 => "0000000010100010",
11064 => "0000000010100011",
11065 => "0000000010100011",
11066 => "0000000010100011",
11067 => "0000000010100011",
11068 => "0000000010100011",
11069 => "0000000010100011",
11070 => "0000000010100011",
11071 => "0000000010100011",
11072 => "0000000010100011",
11073 => "0000000010100011",
11074 => "0000000010100011",
11075 => "0000000010100011",
11076 => "0000000010100011",
11077 => "0000000010100011",
11078 => "0000000010100011",
11079 => "0000000010100011",
11080 => "0000000010100011",
11081 => "0000000010100011",
11082 => "0000000010100011",
11083 => "0000000010100011",
11084 => "0000000010100011",
11085 => "0000000010100011",
11086 => "0000000010100011",
11087 => "0000000010100011",
11088 => "0000000010100011",
11089 => "0000000010100100",
11090 => "0000000010100100",
11091 => "0000000010100100",
11092 => "0000000010100100",
11093 => "0000000010100100",
11094 => "0000000010100100",
11095 => "0000000010100100",
11096 => "0000000010100100",
11097 => "0000000010100100",
11098 => "0000000010100100",
11099 => "0000000010100100",
11100 => "0000000010100100",
11101 => "0000000010100100",
11102 => "0000000010100100",
11103 => "0000000010100100",
11104 => "0000000010100100",
11105 => "0000000010100100",
11106 => "0000000010100100",
11107 => "0000000010100100",
11108 => "0000000010100100",
11109 => "0000000010100100",
11110 => "0000000010100100",
11111 => "0000000010100100",
11112 => "0000000010100100",
11113 => "0000000010100100",
11114 => "0000000010100101",
11115 => "0000000010100101",
11116 => "0000000010100101",
11117 => "0000000010100101",
11118 => "0000000010100101",
11119 => "0000000010100101",
11120 => "0000000010100101",
11121 => "0000000010100101",
11122 => "0000000010100101",
11123 => "0000000010100101",
11124 => "0000000010100101",
11125 => "0000000010100101",
11126 => "0000000010100101",
11127 => "0000000010100101",
11128 => "0000000010100101",
11129 => "0000000010100101",
11130 => "0000000010100101",
11131 => "0000000010100101",
11132 => "0000000010100101",
11133 => "0000000010100101",
11134 => "0000000010100101",
11135 => "0000000010100101",
11136 => "0000000010100101",
11137 => "0000000010100101",
11138 => "0000000010100101",
11139 => "0000000010100110",
11140 => "0000000010100110",
11141 => "0000000010100110",
11142 => "0000000010100110",
11143 => "0000000010100110",
11144 => "0000000010100110",
11145 => "0000000010100110",
11146 => "0000000010100110",
11147 => "0000000010100110",
11148 => "0000000010100110",
11149 => "0000000010100110",
11150 => "0000000010100110",
11151 => "0000000010100110",
11152 => "0000000010100110",
11153 => "0000000010100110",
11154 => "0000000010100110",
11155 => "0000000010100110",
11156 => "0000000010100110",
11157 => "0000000010100110",
11158 => "0000000010100110",
11159 => "0000000010100110",
11160 => "0000000010100110",
11161 => "0000000010100110",
11162 => "0000000010100110",
11163 => "0000000010100110",
11164 => "0000000010100111",
11165 => "0000000010100111",
11166 => "0000000010100111",
11167 => "0000000010100111",
11168 => "0000000010100111",
11169 => "0000000010100111",
11170 => "0000000010100111",
11171 => "0000000010100111",
11172 => "0000000010100111",
11173 => "0000000010100111",
11174 => "0000000010100111",
11175 => "0000000010100111",
11176 => "0000000010100111",
11177 => "0000000010100111",
11178 => "0000000010100111",
11179 => "0000000010100111",
11180 => "0000000010100111",
11181 => "0000000010100111",
11182 => "0000000010100111",
11183 => "0000000010100111",
11184 => "0000000010100111",
11185 => "0000000010100111",
11186 => "0000000010100111",
11187 => "0000000010100111",
11188 => "0000000010100111",
11189 => "0000000010101000",
11190 => "0000000010101000",
11191 => "0000000010101000",
11192 => "0000000010101000",
11193 => "0000000010101000",
11194 => "0000000010101000",
11195 => "0000000010101000",
11196 => "0000000010101000",
11197 => "0000000010101000",
11198 => "0000000010101000",
11199 => "0000000010101000",
11200 => "0000000010101000",
11201 => "0000000010101000",
11202 => "0000000010101000",
11203 => "0000000010101000",
11204 => "0000000010101000",
11205 => "0000000010101000",
11206 => "0000000010101000",
11207 => "0000000010101000",
11208 => "0000000010101000",
11209 => "0000000010101000",
11210 => "0000000010101000",
11211 => "0000000010101000",
11212 => "0000000010101000",
11213 => "0000000010101001",
11214 => "0000000010101001",
11215 => "0000000010101001",
11216 => "0000000010101001",
11217 => "0000000010101001",
11218 => "0000000010101001",
11219 => "0000000010101001",
11220 => "0000000010101001",
11221 => "0000000010101001",
11222 => "0000000010101001",
11223 => "0000000010101001",
11224 => "0000000010101001",
11225 => "0000000010101001",
11226 => "0000000010101001",
11227 => "0000000010101001",
11228 => "0000000010101001",
11229 => "0000000010101001",
11230 => "0000000010101001",
11231 => "0000000010101001",
11232 => "0000000010101001",
11233 => "0000000010101001",
11234 => "0000000010101001",
11235 => "0000000010101001",
11236 => "0000000010101001",
11237 => "0000000010101010",
11238 => "0000000010101010",
11239 => "0000000010101010",
11240 => "0000000010101010",
11241 => "0000000010101010",
11242 => "0000000010101010",
11243 => "0000000010101010",
11244 => "0000000010101010",
11245 => "0000000010101010",
11246 => "0000000010101010",
11247 => "0000000010101010",
11248 => "0000000010101010",
11249 => "0000000010101010",
11250 => "0000000010101010",
11251 => "0000000010101010",
11252 => "0000000010101010",
11253 => "0000000010101010",
11254 => "0000000010101010",
11255 => "0000000010101010",
11256 => "0000000010101010",
11257 => "0000000010101010",
11258 => "0000000010101010",
11259 => "0000000010101010",
11260 => "0000000010101010",
11261 => "0000000010101010",
11262 => "0000000010101011",
11263 => "0000000010101011",
11264 => "0000000010101011",
11265 => "0000000010101011",
11266 => "0000000010101011",
11267 => "0000000010101011",
11268 => "0000000010101011",
11269 => "0000000010101011",
11270 => "0000000010101011",
11271 => "0000000010101011",
11272 => "0000000010101011",
11273 => "0000000010101011",
11274 => "0000000010101011",
11275 => "0000000010101011",
11276 => "0000000010101011",
11277 => "0000000010101011",
11278 => "0000000010101011",
11279 => "0000000010101011",
11280 => "0000000010101011",
11281 => "0000000010101011",
11282 => "0000000010101011",
11283 => "0000000010101011",
11284 => "0000000010101011",
11285 => "0000000010101011",
11286 => "0000000010101100",
11287 => "0000000010101100",
11288 => "0000000010101100",
11289 => "0000000010101100",
11290 => "0000000010101100",
11291 => "0000000010101100",
11292 => "0000000010101100",
11293 => "0000000010101100",
11294 => "0000000010101100",
11295 => "0000000010101100",
11296 => "0000000010101100",
11297 => "0000000010101100",
11298 => "0000000010101100",
11299 => "0000000010101100",
11300 => "0000000010101100",
11301 => "0000000010101100",
11302 => "0000000010101100",
11303 => "0000000010101100",
11304 => "0000000010101100",
11305 => "0000000010101100",
11306 => "0000000010101100",
11307 => "0000000010101100",
11308 => "0000000010101100",
11309 => "0000000010101101",
11310 => "0000000010101101",
11311 => "0000000010101101",
11312 => "0000000010101101",
11313 => "0000000010101101",
11314 => "0000000010101101",
11315 => "0000000010101101",
11316 => "0000000010101101",
11317 => "0000000010101101",
11318 => "0000000010101101",
11319 => "0000000010101101",
11320 => "0000000010101101",
11321 => "0000000010101101",
11322 => "0000000010101101",
11323 => "0000000010101101",
11324 => "0000000010101101",
11325 => "0000000010101101",
11326 => "0000000010101101",
11327 => "0000000010101101",
11328 => "0000000010101101",
11329 => "0000000010101101",
11330 => "0000000010101101",
11331 => "0000000010101101",
11332 => "0000000010101101",
11333 => "0000000010101110",
11334 => "0000000010101110",
11335 => "0000000010101110",
11336 => "0000000010101110",
11337 => "0000000010101110",
11338 => "0000000010101110",
11339 => "0000000010101110",
11340 => "0000000010101110",
11341 => "0000000010101110",
11342 => "0000000010101110",
11343 => "0000000010101110",
11344 => "0000000010101110",
11345 => "0000000010101110",
11346 => "0000000010101110",
11347 => "0000000010101110",
11348 => "0000000010101110",
11349 => "0000000010101110",
11350 => "0000000010101110",
11351 => "0000000010101110",
11352 => "0000000010101110",
11353 => "0000000010101110",
11354 => "0000000010101110",
11355 => "0000000010101110",
11356 => "0000000010101110",
11357 => "0000000010101111",
11358 => "0000000010101111",
11359 => "0000000010101111",
11360 => "0000000010101111",
11361 => "0000000010101111",
11362 => "0000000010101111",
11363 => "0000000010101111",
11364 => "0000000010101111",
11365 => "0000000010101111",
11366 => "0000000010101111",
11367 => "0000000010101111",
11368 => "0000000010101111",
11369 => "0000000010101111",
11370 => "0000000010101111",
11371 => "0000000010101111",
11372 => "0000000010101111",
11373 => "0000000010101111",
11374 => "0000000010101111",
11375 => "0000000010101111",
11376 => "0000000010101111",
11377 => "0000000010101111",
11378 => "0000000010101111",
11379 => "0000000010101111",
11380 => "0000000010110000",
11381 => "0000000010110000",
11382 => "0000000010110000",
11383 => "0000000010110000",
11384 => "0000000010110000",
11385 => "0000000010110000",
11386 => "0000000010110000",
11387 => "0000000010110000",
11388 => "0000000010110000",
11389 => "0000000010110000",
11390 => "0000000010110000",
11391 => "0000000010110000",
11392 => "0000000010110000",
11393 => "0000000010110000",
11394 => "0000000010110000",
11395 => "0000000010110000",
11396 => "0000000010110000",
11397 => "0000000010110000",
11398 => "0000000010110000",
11399 => "0000000010110000",
11400 => "0000000010110000",
11401 => "0000000010110000",
11402 => "0000000010110000",
11403 => "0000000010110000",
11404 => "0000000010110001",
11405 => "0000000010110001",
11406 => "0000000010110001",
11407 => "0000000010110001",
11408 => "0000000010110001",
11409 => "0000000010110001",
11410 => "0000000010110001",
11411 => "0000000010110001",
11412 => "0000000010110001",
11413 => "0000000010110001",
11414 => "0000000010110001",
11415 => "0000000010110001",
11416 => "0000000010110001",
11417 => "0000000010110001",
11418 => "0000000010110001",
11419 => "0000000010110001",
11420 => "0000000010110001",
11421 => "0000000010110001",
11422 => "0000000010110001",
11423 => "0000000010110001",
11424 => "0000000010110001",
11425 => "0000000010110001",
11426 => "0000000010110001",
11427 => "0000000010110010",
11428 => "0000000010110010",
11429 => "0000000010110010",
11430 => "0000000010110010",
11431 => "0000000010110010",
11432 => "0000000010110010",
11433 => "0000000010110010",
11434 => "0000000010110010",
11435 => "0000000010110010",
11436 => "0000000010110010",
11437 => "0000000010110010",
11438 => "0000000010110010",
11439 => "0000000010110010",
11440 => "0000000010110010",
11441 => "0000000010110010",
11442 => "0000000010110010",
11443 => "0000000010110010",
11444 => "0000000010110010",
11445 => "0000000010110010",
11446 => "0000000010110010",
11447 => "0000000010110010",
11448 => "0000000010110010",
11449 => "0000000010110010",
11450 => "0000000010110011",
11451 => "0000000010110011",
11452 => "0000000010110011",
11453 => "0000000010110011",
11454 => "0000000010110011",
11455 => "0000000010110011",
11456 => "0000000010110011",
11457 => "0000000010110011",
11458 => "0000000010110011",
11459 => "0000000010110011",
11460 => "0000000010110011",
11461 => "0000000010110011",
11462 => "0000000010110011",
11463 => "0000000010110011",
11464 => "0000000010110011",
11465 => "0000000010110011",
11466 => "0000000010110011",
11467 => "0000000010110011",
11468 => "0000000010110011",
11469 => "0000000010110011",
11470 => "0000000010110011",
11471 => "0000000010110011",
11472 => "0000000010110011",
11473 => "0000000010110100",
11474 => "0000000010110100",
11475 => "0000000010110100",
11476 => "0000000010110100",
11477 => "0000000010110100",
11478 => "0000000010110100",
11479 => "0000000010110100",
11480 => "0000000010110100",
11481 => "0000000010110100",
11482 => "0000000010110100",
11483 => "0000000010110100",
11484 => "0000000010110100",
11485 => "0000000010110100",
11486 => "0000000010110100",
11487 => "0000000010110100",
11488 => "0000000010110100",
11489 => "0000000010110100",
11490 => "0000000010110100",
11491 => "0000000010110100",
11492 => "0000000010110100",
11493 => "0000000010110100",
11494 => "0000000010110100",
11495 => "0000000010110100",
11496 => "0000000010110101",
11497 => "0000000010110101",
11498 => "0000000010110101",
11499 => "0000000010110101",
11500 => "0000000010110101",
11501 => "0000000010110101",
11502 => "0000000010110101",
11503 => "0000000010110101",
11504 => "0000000010110101",
11505 => "0000000010110101",
11506 => "0000000010110101",
11507 => "0000000010110101",
11508 => "0000000010110101",
11509 => "0000000010110101",
11510 => "0000000010110101",
11511 => "0000000010110101",
11512 => "0000000010110101",
11513 => "0000000010110101",
11514 => "0000000010110101",
11515 => "0000000010110101",
11516 => "0000000010110101",
11517 => "0000000010110101",
11518 => "0000000010110110",
11519 => "0000000010110110",
11520 => "0000000010110110",
11521 => "0000000010110110",
11522 => "0000000010110110",
11523 => "0000000010110110",
11524 => "0000000010110110",
11525 => "0000000010110110",
11526 => "0000000010110110",
11527 => "0000000010110110",
11528 => "0000000010110110",
11529 => "0000000010110110",
11530 => "0000000010110110",
11531 => "0000000010110110",
11532 => "0000000010110110",
11533 => "0000000010110110",
11534 => "0000000010110110",
11535 => "0000000010110110",
11536 => "0000000010110110",
11537 => "0000000010110110",
11538 => "0000000010110110",
11539 => "0000000010110110",
11540 => "0000000010110110",
11541 => "0000000010110111",
11542 => "0000000010110111",
11543 => "0000000010110111",
11544 => "0000000010110111",
11545 => "0000000010110111",
11546 => "0000000010110111",
11547 => "0000000010110111",
11548 => "0000000010110111",
11549 => "0000000010110111",
11550 => "0000000010110111",
11551 => "0000000010110111",
11552 => "0000000010110111",
11553 => "0000000010110111",
11554 => "0000000010110111",
11555 => "0000000010110111",
11556 => "0000000010110111",
11557 => "0000000010110111",
11558 => "0000000010110111",
11559 => "0000000010110111",
11560 => "0000000010110111",
11561 => "0000000010110111",
11562 => "0000000010110111",
11563 => "0000000010111000",
11564 => "0000000010111000",
11565 => "0000000010111000",
11566 => "0000000010111000",
11567 => "0000000010111000",
11568 => "0000000010111000",
11569 => "0000000010111000",
11570 => "0000000010111000",
11571 => "0000000010111000",
11572 => "0000000010111000",
11573 => "0000000010111000",
11574 => "0000000010111000",
11575 => "0000000010111000",
11576 => "0000000010111000",
11577 => "0000000010111000",
11578 => "0000000010111000",
11579 => "0000000010111000",
11580 => "0000000010111000",
11581 => "0000000010111000",
11582 => "0000000010111000",
11583 => "0000000010111000",
11584 => "0000000010111000",
11585 => "0000000010111000",
11586 => "0000000010111001",
11587 => "0000000010111001",
11588 => "0000000010111001",
11589 => "0000000010111001",
11590 => "0000000010111001",
11591 => "0000000010111001",
11592 => "0000000010111001",
11593 => "0000000010111001",
11594 => "0000000010111001",
11595 => "0000000010111001",
11596 => "0000000010111001",
11597 => "0000000010111001",
11598 => "0000000010111001",
11599 => "0000000010111001",
11600 => "0000000010111001",
11601 => "0000000010111001",
11602 => "0000000010111001",
11603 => "0000000010111001",
11604 => "0000000010111001",
11605 => "0000000010111001",
11606 => "0000000010111001",
11607 => "0000000010111001",
11608 => "0000000010111010",
11609 => "0000000010111010",
11610 => "0000000010111010",
11611 => "0000000010111010",
11612 => "0000000010111010",
11613 => "0000000010111010",
11614 => "0000000010111010",
11615 => "0000000010111010",
11616 => "0000000010111010",
11617 => "0000000010111010",
11618 => "0000000010111010",
11619 => "0000000010111010",
11620 => "0000000010111010",
11621 => "0000000010111010",
11622 => "0000000010111010",
11623 => "0000000010111010",
11624 => "0000000010111010",
11625 => "0000000010111010",
11626 => "0000000010111010",
11627 => "0000000010111010",
11628 => "0000000010111010",
11629 => "0000000010111010",
11630 => "0000000010111011",
11631 => "0000000010111011",
11632 => "0000000010111011",
11633 => "0000000010111011",
11634 => "0000000010111011",
11635 => "0000000010111011",
11636 => "0000000010111011",
11637 => "0000000010111011",
11638 => "0000000010111011",
11639 => "0000000010111011",
11640 => "0000000010111011",
11641 => "0000000010111011",
11642 => "0000000010111011",
11643 => "0000000010111011",
11644 => "0000000010111011",
11645 => "0000000010111011",
11646 => "0000000010111011",
11647 => "0000000010111011",
11648 => "0000000010111011",
11649 => "0000000010111011",
11650 => "0000000010111011",
11651 => "0000000010111011",
11652 => "0000000010111100",
11653 => "0000000010111100",
11654 => "0000000010111100",
11655 => "0000000010111100",
11656 => "0000000010111100",
11657 => "0000000010111100",
11658 => "0000000010111100",
11659 => "0000000010111100",
11660 => "0000000010111100",
11661 => "0000000010111100",
11662 => "0000000010111100",
11663 => "0000000010111100",
11664 => "0000000010111100",
11665 => "0000000010111100",
11666 => "0000000010111100",
11667 => "0000000010111100",
11668 => "0000000010111100",
11669 => "0000000010111100",
11670 => "0000000010111100",
11671 => "0000000010111100",
11672 => "0000000010111100",
11673 => "0000000010111100",
11674 => "0000000010111101",
11675 => "0000000010111101",
11676 => "0000000010111101",
11677 => "0000000010111101",
11678 => "0000000010111101",
11679 => "0000000010111101",
11680 => "0000000010111101",
11681 => "0000000010111101",
11682 => "0000000010111101",
11683 => "0000000010111101",
11684 => "0000000010111101",
11685 => "0000000010111101",
11686 => "0000000010111101",
11687 => "0000000010111101",
11688 => "0000000010111101",
11689 => "0000000010111101",
11690 => "0000000010111101",
11691 => "0000000010111101",
11692 => "0000000010111101",
11693 => "0000000010111101",
11694 => "0000000010111101",
11695 => "0000000010111101",
11696 => "0000000010111110",
11697 => "0000000010111110",
11698 => "0000000010111110",
11699 => "0000000010111110",
11700 => "0000000010111110",
11701 => "0000000010111110",
11702 => "0000000010111110",
11703 => "0000000010111110",
11704 => "0000000010111110",
11705 => "0000000010111110",
11706 => "0000000010111110",
11707 => "0000000010111110",
11708 => "0000000010111110",
11709 => "0000000010111110",
11710 => "0000000010111110",
11711 => "0000000010111110",
11712 => "0000000010111110",
11713 => "0000000010111110",
11714 => "0000000010111110",
11715 => "0000000010111110",
11716 => "0000000010111110",
11717 => "0000000010111111",
11718 => "0000000010111111",
11719 => "0000000010111111",
11720 => "0000000010111111",
11721 => "0000000010111111",
11722 => "0000000010111111",
11723 => "0000000010111111",
11724 => "0000000010111111",
11725 => "0000000010111111",
11726 => "0000000010111111",
11727 => "0000000010111111",
11728 => "0000000010111111",
11729 => "0000000010111111",
11730 => "0000000010111111",
11731 => "0000000010111111",
11732 => "0000000010111111",
11733 => "0000000010111111",
11734 => "0000000010111111",
11735 => "0000000010111111",
11736 => "0000000010111111",
11737 => "0000000010111111",
11738 => "0000000010111111",
11739 => "0000000011000000",
11740 => "0000000011000000",
11741 => "0000000011000000",
11742 => "0000000011000000",
11743 => "0000000011000000",
11744 => "0000000011000000",
11745 => "0000000011000000",
11746 => "0000000011000000",
11747 => "0000000011000000",
11748 => "0000000011000000",
11749 => "0000000011000000",
11750 => "0000000011000000",
11751 => "0000000011000000",
11752 => "0000000011000000",
11753 => "0000000011000000",
11754 => "0000000011000000",
11755 => "0000000011000000",
11756 => "0000000011000000",
11757 => "0000000011000000",
11758 => "0000000011000000",
11759 => "0000000011000000",
11760 => "0000000011000001",
11761 => "0000000011000001",
11762 => "0000000011000001",
11763 => "0000000011000001",
11764 => "0000000011000001",
11765 => "0000000011000001",
11766 => "0000000011000001",
11767 => "0000000011000001",
11768 => "0000000011000001",
11769 => "0000000011000001",
11770 => "0000000011000001",
11771 => "0000000011000001",
11772 => "0000000011000001",
11773 => "0000000011000001",
11774 => "0000000011000001",
11775 => "0000000011000001",
11776 => "0000000011000001",
11777 => "0000000011000001",
11778 => "0000000011000001",
11779 => "0000000011000001",
11780 => "0000000011000001",
11781 => "0000000011000010",
11782 => "0000000011000010",
11783 => "0000000011000010",
11784 => "0000000011000010",
11785 => "0000000011000010",
11786 => "0000000011000010",
11787 => "0000000011000010",
11788 => "0000000011000010",
11789 => "0000000011000010",
11790 => "0000000011000010",
11791 => "0000000011000010",
11792 => "0000000011000010",
11793 => "0000000011000010",
11794 => "0000000011000010",
11795 => "0000000011000010",
11796 => "0000000011000010",
11797 => "0000000011000010",
11798 => "0000000011000010",
11799 => "0000000011000010",
11800 => "0000000011000010",
11801 => "0000000011000010",
11802 => "0000000011000010",
11803 => "0000000011000011",
11804 => "0000000011000011",
11805 => "0000000011000011",
11806 => "0000000011000011",
11807 => "0000000011000011",
11808 => "0000000011000011",
11809 => "0000000011000011",
11810 => "0000000011000011",
11811 => "0000000011000011",
11812 => "0000000011000011",
11813 => "0000000011000011",
11814 => "0000000011000011",
11815 => "0000000011000011",
11816 => "0000000011000011",
11817 => "0000000011000011",
11818 => "0000000011000011",
11819 => "0000000011000011",
11820 => "0000000011000011",
11821 => "0000000011000011",
11822 => "0000000011000011",
11823 => "0000000011000011",
11824 => "0000000011000100",
11825 => "0000000011000100",
11826 => "0000000011000100",
11827 => "0000000011000100",
11828 => "0000000011000100",
11829 => "0000000011000100",
11830 => "0000000011000100",
11831 => "0000000011000100",
11832 => "0000000011000100",
11833 => "0000000011000100",
11834 => "0000000011000100",
11835 => "0000000011000100",
11836 => "0000000011000100",
11837 => "0000000011000100",
11838 => "0000000011000100",
11839 => "0000000011000100",
11840 => "0000000011000100",
11841 => "0000000011000100",
11842 => "0000000011000100",
11843 => "0000000011000100",
11844 => "0000000011000100",
11845 => "0000000011000101",
11846 => "0000000011000101",
11847 => "0000000011000101",
11848 => "0000000011000101",
11849 => "0000000011000101",
11850 => "0000000011000101",
11851 => "0000000011000101",
11852 => "0000000011000101",
11853 => "0000000011000101",
11854 => "0000000011000101",
11855 => "0000000011000101",
11856 => "0000000011000101",
11857 => "0000000011000101",
11858 => "0000000011000101",
11859 => "0000000011000101",
11860 => "0000000011000101",
11861 => "0000000011000101",
11862 => "0000000011000101",
11863 => "0000000011000101",
11864 => "0000000011000101",
11865 => "0000000011000101",
11866 => "0000000011000110",
11867 => "0000000011000110",
11868 => "0000000011000110",
11869 => "0000000011000110",
11870 => "0000000011000110",
11871 => "0000000011000110",
11872 => "0000000011000110",
11873 => "0000000011000110",
11874 => "0000000011000110",
11875 => "0000000011000110",
11876 => "0000000011000110",
11877 => "0000000011000110",
11878 => "0000000011000110",
11879 => "0000000011000110",
11880 => "0000000011000110",
11881 => "0000000011000110",
11882 => "0000000011000110",
11883 => "0000000011000110",
11884 => "0000000011000110",
11885 => "0000000011000110",
11886 => "0000000011000111",
11887 => "0000000011000111",
11888 => "0000000011000111",
11889 => "0000000011000111",
11890 => "0000000011000111",
11891 => "0000000011000111",
11892 => "0000000011000111",
11893 => "0000000011000111",
11894 => "0000000011000111",
11895 => "0000000011000111",
11896 => "0000000011000111",
11897 => "0000000011000111",
11898 => "0000000011000111",
11899 => "0000000011000111",
11900 => "0000000011000111",
11901 => "0000000011000111",
11902 => "0000000011000111",
11903 => "0000000011000111",
11904 => "0000000011000111",
11905 => "0000000011000111",
11906 => "0000000011000111",
11907 => "0000000011001000",
11908 => "0000000011001000",
11909 => "0000000011001000",
11910 => "0000000011001000",
11911 => "0000000011001000",
11912 => "0000000011001000",
11913 => "0000000011001000",
11914 => "0000000011001000",
11915 => "0000000011001000",
11916 => "0000000011001000",
11917 => "0000000011001000",
11918 => "0000000011001000",
11919 => "0000000011001000",
11920 => "0000000011001000",
11921 => "0000000011001000",
11922 => "0000000011001000",
11923 => "0000000011001000",
11924 => "0000000011001000",
11925 => "0000000011001000",
11926 => "0000000011001000",
11927 => "0000000011001000",
11928 => "0000000011001001",
11929 => "0000000011001001",
11930 => "0000000011001001",
11931 => "0000000011001001",
11932 => "0000000011001001",
11933 => "0000000011001001",
11934 => "0000000011001001",
11935 => "0000000011001001",
11936 => "0000000011001001",
11937 => "0000000011001001",
11938 => "0000000011001001",
11939 => "0000000011001001",
11940 => "0000000011001001",
11941 => "0000000011001001",
11942 => "0000000011001001",
11943 => "0000000011001001",
11944 => "0000000011001001",
11945 => "0000000011001001",
11946 => "0000000011001001",
11947 => "0000000011001001",
11948 => "0000000011001010",
11949 => "0000000011001010",
11950 => "0000000011001010",
11951 => "0000000011001010",
11952 => "0000000011001010",
11953 => "0000000011001010",
11954 => "0000000011001010",
11955 => "0000000011001010",
11956 => "0000000011001010",
11957 => "0000000011001010",
11958 => "0000000011001010",
11959 => "0000000011001010",
11960 => "0000000011001010",
11961 => "0000000011001010",
11962 => "0000000011001010",
11963 => "0000000011001010",
11964 => "0000000011001010",
11965 => "0000000011001010",
11966 => "0000000011001010",
11967 => "0000000011001010",
11968 => "0000000011001011",
11969 => "0000000011001011",
11970 => "0000000011001011",
11971 => "0000000011001011",
11972 => "0000000011001011",
11973 => "0000000011001011",
11974 => "0000000011001011",
11975 => "0000000011001011",
11976 => "0000000011001011",
11977 => "0000000011001011",
11978 => "0000000011001011",
11979 => "0000000011001011",
11980 => "0000000011001011",
11981 => "0000000011001011",
11982 => "0000000011001011",
11983 => "0000000011001011",
11984 => "0000000011001011",
11985 => "0000000011001011",
11986 => "0000000011001011",
11987 => "0000000011001011",
11988 => "0000000011001011",
11989 => "0000000011001100",
11990 => "0000000011001100",
11991 => "0000000011001100",
11992 => "0000000011001100",
11993 => "0000000011001100",
11994 => "0000000011001100",
11995 => "0000000011001100",
11996 => "0000000011001100",
11997 => "0000000011001100",
11998 => "0000000011001100",
11999 => "0000000011001100",
12000 => "0000000011001100",
12001 => "0000000011001100",
12002 => "0000000011001100",
12003 => "0000000011001100",
12004 => "0000000011001100",
12005 => "0000000011001100",
12006 => "0000000011001100",
12007 => "0000000011001100",
12008 => "0000000011001100",
12009 => "0000000011001101",
12010 => "0000000011001101",
12011 => "0000000011001101",
12012 => "0000000011001101",
12013 => "0000000011001101",
12014 => "0000000011001101",
12015 => "0000000011001101",
12016 => "0000000011001101",
12017 => "0000000011001101",
12018 => "0000000011001101",
12019 => "0000000011001101",
12020 => "0000000011001101",
12021 => "0000000011001101",
12022 => "0000000011001101",
12023 => "0000000011001101",
12024 => "0000000011001101",
12025 => "0000000011001101",
12026 => "0000000011001101",
12027 => "0000000011001101",
12028 => "0000000011001101",
12029 => "0000000011001110",
12030 => "0000000011001110",
12031 => "0000000011001110",
12032 => "0000000011001110",
12033 => "0000000011001110",
12034 => "0000000011001110",
12035 => "0000000011001110",
12036 => "0000000011001110",
12037 => "0000000011001110",
12038 => "0000000011001110",
12039 => "0000000011001110",
12040 => "0000000011001110",
12041 => "0000000011001110",
12042 => "0000000011001110",
12043 => "0000000011001110",
12044 => "0000000011001110",
12045 => "0000000011001110",
12046 => "0000000011001110",
12047 => "0000000011001110",
12048 => "0000000011001110",
12049 => "0000000011001111",
12050 => "0000000011001111",
12051 => "0000000011001111",
12052 => "0000000011001111",
12053 => "0000000011001111",
12054 => "0000000011001111",
12055 => "0000000011001111",
12056 => "0000000011001111",
12057 => "0000000011001111",
12058 => "0000000011001111",
12059 => "0000000011001111",
12060 => "0000000011001111",
12061 => "0000000011001111",
12062 => "0000000011001111",
12063 => "0000000011001111",
12064 => "0000000011001111",
12065 => "0000000011001111",
12066 => "0000000011001111",
12067 => "0000000011001111",
12068 => "0000000011001111",
12069 => "0000000011010000",
12070 => "0000000011010000",
12071 => "0000000011010000",
12072 => "0000000011010000",
12073 => "0000000011010000",
12074 => "0000000011010000",
12075 => "0000000011010000",
12076 => "0000000011010000",
12077 => "0000000011010000",
12078 => "0000000011010000",
12079 => "0000000011010000",
12080 => "0000000011010000",
12081 => "0000000011010000",
12082 => "0000000011010000",
12083 => "0000000011010000",
12084 => "0000000011010000",
12085 => "0000000011010000",
12086 => "0000000011010000",
12087 => "0000000011010000",
12088 => "0000000011010000",
12089 => "0000000011010001",
12090 => "0000000011010001",
12091 => "0000000011010001",
12092 => "0000000011010001",
12093 => "0000000011010001",
12094 => "0000000011010001",
12095 => "0000000011010001",
12096 => "0000000011010001",
12097 => "0000000011010001",
12098 => "0000000011010001",
12099 => "0000000011010001",
12100 => "0000000011010001",
12101 => "0000000011010001",
12102 => "0000000011010001",
12103 => "0000000011010001",
12104 => "0000000011010001",
12105 => "0000000011010001",
12106 => "0000000011010001",
12107 => "0000000011010001",
12108 => "0000000011010010",
12109 => "0000000011010010",
12110 => "0000000011010010",
12111 => "0000000011010010",
12112 => "0000000011010010",
12113 => "0000000011010010",
12114 => "0000000011010010",
12115 => "0000000011010010",
12116 => "0000000011010010",
12117 => "0000000011010010",
12118 => "0000000011010010",
12119 => "0000000011010010",
12120 => "0000000011010010",
12121 => "0000000011010010",
12122 => "0000000011010010",
12123 => "0000000011010010",
12124 => "0000000011010010",
12125 => "0000000011010010",
12126 => "0000000011010010",
12127 => "0000000011010010",
12128 => "0000000011010011",
12129 => "0000000011010011",
12130 => "0000000011010011",
12131 => "0000000011010011",
12132 => "0000000011010011",
12133 => "0000000011010011",
12134 => "0000000011010011",
12135 => "0000000011010011",
12136 => "0000000011010011",
12137 => "0000000011010011",
12138 => "0000000011010011",
12139 => "0000000011010011",
12140 => "0000000011010011",
12141 => "0000000011010011",
12142 => "0000000011010011",
12143 => "0000000011010011",
12144 => "0000000011010011",
12145 => "0000000011010011",
12146 => "0000000011010011",
12147 => "0000000011010100",
12148 => "0000000011010100",
12149 => "0000000011010100",
12150 => "0000000011010100",
12151 => "0000000011010100",
12152 => "0000000011010100",
12153 => "0000000011010100",
12154 => "0000000011010100",
12155 => "0000000011010100",
12156 => "0000000011010100",
12157 => "0000000011010100",
12158 => "0000000011010100",
12159 => "0000000011010100",
12160 => "0000000011010100",
12161 => "0000000011010100",
12162 => "0000000011010100",
12163 => "0000000011010100",
12164 => "0000000011010100",
12165 => "0000000011010100",
12166 => "0000000011010100",
12167 => "0000000011010101",
12168 => "0000000011010101",
12169 => "0000000011010101",
12170 => "0000000011010101",
12171 => "0000000011010101",
12172 => "0000000011010101",
12173 => "0000000011010101",
12174 => "0000000011010101",
12175 => "0000000011010101",
12176 => "0000000011010101",
12177 => "0000000011010101",
12178 => "0000000011010101",
12179 => "0000000011010101",
12180 => "0000000011010101",
12181 => "0000000011010101",
12182 => "0000000011010101",
12183 => "0000000011010101",
12184 => "0000000011010101",
12185 => "0000000011010101",
12186 => "0000000011010110",
12187 => "0000000011010110",
12188 => "0000000011010110",
12189 => "0000000011010110",
12190 => "0000000011010110",
12191 => "0000000011010110",
12192 => "0000000011010110",
12193 => "0000000011010110",
12194 => "0000000011010110",
12195 => "0000000011010110",
12196 => "0000000011010110",
12197 => "0000000011010110",
12198 => "0000000011010110",
12199 => "0000000011010110",
12200 => "0000000011010110",
12201 => "0000000011010110",
12202 => "0000000011010110",
12203 => "0000000011010110",
12204 => "0000000011010110",
12205 => "0000000011010111",
12206 => "0000000011010111",
12207 => "0000000011010111",
12208 => "0000000011010111",
12209 => "0000000011010111",
12210 => "0000000011010111",
12211 => "0000000011010111",
12212 => "0000000011010111",
12213 => "0000000011010111",
12214 => "0000000011010111",
12215 => "0000000011010111",
12216 => "0000000011010111",
12217 => "0000000011010111",
12218 => "0000000011010111",
12219 => "0000000011010111",
12220 => "0000000011010111",
12221 => "0000000011010111",
12222 => "0000000011010111",
12223 => "0000000011010111",
12224 => "0000000011011000",
12225 => "0000000011011000",
12226 => "0000000011011000",
12227 => "0000000011011000",
12228 => "0000000011011000",
12229 => "0000000011011000",
12230 => "0000000011011000",
12231 => "0000000011011000",
12232 => "0000000011011000",
12233 => "0000000011011000",
12234 => "0000000011011000",
12235 => "0000000011011000",
12236 => "0000000011011000",
12237 => "0000000011011000",
12238 => "0000000011011000",
12239 => "0000000011011000",
12240 => "0000000011011000",
12241 => "0000000011011000",
12242 => "0000000011011000",
12243 => "0000000011011001",
12244 => "0000000011011001",
12245 => "0000000011011001",
12246 => "0000000011011001",
12247 => "0000000011011001",
12248 => "0000000011011001",
12249 => "0000000011011001",
12250 => "0000000011011001",
12251 => "0000000011011001",
12252 => "0000000011011001",
12253 => "0000000011011001",
12254 => "0000000011011001",
12255 => "0000000011011001",
12256 => "0000000011011001",
12257 => "0000000011011001",
12258 => "0000000011011001",
12259 => "0000000011011001",
12260 => "0000000011011001",
12261 => "0000000011011001",
12262 => "0000000011011010",
12263 => "0000000011011010",
12264 => "0000000011011010",
12265 => "0000000011011010",
12266 => "0000000011011010",
12267 => "0000000011011010",
12268 => "0000000011011010",
12269 => "0000000011011010",
12270 => "0000000011011010",
12271 => "0000000011011010",
12272 => "0000000011011010",
12273 => "0000000011011010",
12274 => "0000000011011010",
12275 => "0000000011011010",
12276 => "0000000011011010",
12277 => "0000000011011010",
12278 => "0000000011011010",
12279 => "0000000011011010",
12280 => "0000000011011010",
12281 => "0000000011011011",
12282 => "0000000011011011",
12283 => "0000000011011011",
12284 => "0000000011011011",
12285 => "0000000011011011",
12286 => "0000000011011011",
12287 => "0000000011011011",
12288 => "0000000011011011",
12289 => "0000000011011011",
12290 => "0000000011011011",
12291 => "0000000011011011",
12292 => "0000000011011011",
12293 => "0000000011011011",
12294 => "0000000011011011",
12295 => "0000000011011011",
12296 => "0000000011011011",
12297 => "0000000011011011",
12298 => "0000000011011011",
12299 => "0000000011011011",
12300 => "0000000011011100",
12301 => "0000000011011100",
12302 => "0000000011011100",
12303 => "0000000011011100",
12304 => "0000000011011100",
12305 => "0000000011011100",
12306 => "0000000011011100",
12307 => "0000000011011100",
12308 => "0000000011011100",
12309 => "0000000011011100",
12310 => "0000000011011100",
12311 => "0000000011011100",
12312 => "0000000011011100",
12313 => "0000000011011100",
12314 => "0000000011011100",
12315 => "0000000011011100",
12316 => "0000000011011100",
12317 => "0000000011011100",
12318 => "0000000011011100",
12319 => "0000000011011101",
12320 => "0000000011011101",
12321 => "0000000011011101",
12322 => "0000000011011101",
12323 => "0000000011011101",
12324 => "0000000011011101",
12325 => "0000000011011101",
12326 => "0000000011011101",
12327 => "0000000011011101",
12328 => "0000000011011101",
12329 => "0000000011011101",
12330 => "0000000011011101",
12331 => "0000000011011101",
12332 => "0000000011011101",
12333 => "0000000011011101",
12334 => "0000000011011101",
12335 => "0000000011011101",
12336 => "0000000011011101",
12337 => "0000000011011110",
12338 => "0000000011011110",
12339 => "0000000011011110",
12340 => "0000000011011110",
12341 => "0000000011011110",
12342 => "0000000011011110",
12343 => "0000000011011110",
12344 => "0000000011011110",
12345 => "0000000011011110",
12346 => "0000000011011110",
12347 => "0000000011011110",
12348 => "0000000011011110",
12349 => "0000000011011110",
12350 => "0000000011011110",
12351 => "0000000011011110",
12352 => "0000000011011110",
12353 => "0000000011011110",
12354 => "0000000011011110",
12355 => "0000000011011110",
12356 => "0000000011011111",
12357 => "0000000011011111",
12358 => "0000000011011111",
12359 => "0000000011011111",
12360 => "0000000011011111",
12361 => "0000000011011111",
12362 => "0000000011011111",
12363 => "0000000011011111",
12364 => "0000000011011111",
12365 => "0000000011011111",
12366 => "0000000011011111",
12367 => "0000000011011111",
12368 => "0000000011011111",
12369 => "0000000011011111",
12370 => "0000000011011111",
12371 => "0000000011011111",
12372 => "0000000011011111",
12373 => "0000000011011111",
12374 => "0000000011100000",
12375 => "0000000011100000",
12376 => "0000000011100000",
12377 => "0000000011100000",
12378 => "0000000011100000",
12379 => "0000000011100000",
12380 => "0000000011100000",
12381 => "0000000011100000",
12382 => "0000000011100000",
12383 => "0000000011100000",
12384 => "0000000011100000",
12385 => "0000000011100000",
12386 => "0000000011100000",
12387 => "0000000011100000",
12388 => "0000000011100000",
12389 => "0000000011100000",
12390 => "0000000011100000",
12391 => "0000000011100000",
12392 => "0000000011100000",
12393 => "0000000011100001",
12394 => "0000000011100001",
12395 => "0000000011100001",
12396 => "0000000011100001",
12397 => "0000000011100001",
12398 => "0000000011100001",
12399 => "0000000011100001",
12400 => "0000000011100001",
12401 => "0000000011100001",
12402 => "0000000011100001",
12403 => "0000000011100001",
12404 => "0000000011100001",
12405 => "0000000011100001",
12406 => "0000000011100001",
12407 => "0000000011100001",
12408 => "0000000011100001",
12409 => "0000000011100001",
12410 => "0000000011100001",
12411 => "0000000011100010",
12412 => "0000000011100010",
12413 => "0000000011100010",
12414 => "0000000011100010",
12415 => "0000000011100010",
12416 => "0000000011100010",
12417 => "0000000011100010",
12418 => "0000000011100010",
12419 => "0000000011100010",
12420 => "0000000011100010",
12421 => "0000000011100010",
12422 => "0000000011100010",
12423 => "0000000011100010",
12424 => "0000000011100010",
12425 => "0000000011100010",
12426 => "0000000011100010",
12427 => "0000000011100010",
12428 => "0000000011100010",
12429 => "0000000011100011",
12430 => "0000000011100011",
12431 => "0000000011100011",
12432 => "0000000011100011",
12433 => "0000000011100011",
12434 => "0000000011100011",
12435 => "0000000011100011",
12436 => "0000000011100011",
12437 => "0000000011100011",
12438 => "0000000011100011",
12439 => "0000000011100011",
12440 => "0000000011100011",
12441 => "0000000011100011",
12442 => "0000000011100011",
12443 => "0000000011100011",
12444 => "0000000011100011",
12445 => "0000000011100011",
12446 => "0000000011100011",
12447 => "0000000011100100",
12448 => "0000000011100100",
12449 => "0000000011100100",
12450 => "0000000011100100",
12451 => "0000000011100100",
12452 => "0000000011100100",
12453 => "0000000011100100",
12454 => "0000000011100100",
12455 => "0000000011100100",
12456 => "0000000011100100",
12457 => "0000000011100100",
12458 => "0000000011100100",
12459 => "0000000011100100",
12460 => "0000000011100100",
12461 => "0000000011100100",
12462 => "0000000011100100",
12463 => "0000000011100100",
12464 => "0000000011100100",
12465 => "0000000011100101",
12466 => "0000000011100101",
12467 => "0000000011100101",
12468 => "0000000011100101",
12469 => "0000000011100101",
12470 => "0000000011100101",
12471 => "0000000011100101",
12472 => "0000000011100101",
12473 => "0000000011100101",
12474 => "0000000011100101",
12475 => "0000000011100101",
12476 => "0000000011100101",
12477 => "0000000011100101",
12478 => "0000000011100101",
12479 => "0000000011100101",
12480 => "0000000011100101",
12481 => "0000000011100101",
12482 => "0000000011100101",
12483 => "0000000011100110",
12484 => "0000000011100110",
12485 => "0000000011100110",
12486 => "0000000011100110",
12487 => "0000000011100110",
12488 => "0000000011100110",
12489 => "0000000011100110",
12490 => "0000000011100110",
12491 => "0000000011100110",
12492 => "0000000011100110",
12493 => "0000000011100110",
12494 => "0000000011100110",
12495 => "0000000011100110",
12496 => "0000000011100110",
12497 => "0000000011100110",
12498 => "0000000011100110",
12499 => "0000000011100110",
12500 => "0000000011100110",
12501 => "0000000011100111",
12502 => "0000000011100111",
12503 => "0000000011100111",
12504 => "0000000011100111",
12505 => "0000000011100111",
12506 => "0000000011100111",
12507 => "0000000011100111",
12508 => "0000000011100111",
12509 => "0000000011100111",
12510 => "0000000011100111",
12511 => "0000000011100111",
12512 => "0000000011100111",
12513 => "0000000011100111",
12514 => "0000000011100111",
12515 => "0000000011100111",
12516 => "0000000011100111",
12517 => "0000000011100111",
12518 => "0000000011100111",
12519 => "0000000011101000",
12520 => "0000000011101000",
12521 => "0000000011101000",
12522 => "0000000011101000",
12523 => "0000000011101000",
12524 => "0000000011101000",
12525 => "0000000011101000",
12526 => "0000000011101000",
12527 => "0000000011101000",
12528 => "0000000011101000",
12529 => "0000000011101000",
12530 => "0000000011101000",
12531 => "0000000011101000",
12532 => "0000000011101000",
12533 => "0000000011101000",
12534 => "0000000011101000",
12535 => "0000000011101000",
12536 => "0000000011101000",
12537 => "0000000011101001",
12538 => "0000000011101001",
12539 => "0000000011101001",
12540 => "0000000011101001",
12541 => "0000000011101001",
12542 => "0000000011101001",
12543 => "0000000011101001",
12544 => "0000000011101001",
12545 => "0000000011101001",
12546 => "0000000011101001",
12547 => "0000000011101001",
12548 => "0000000011101001",
12549 => "0000000011101001",
12550 => "0000000011101001",
12551 => "0000000011101001",
12552 => "0000000011101001",
12553 => "0000000011101001",
12554 => "0000000011101001",
12555 => "0000000011101010",
12556 => "0000000011101010",
12557 => "0000000011101010",
12558 => "0000000011101010",
12559 => "0000000011101010",
12560 => "0000000011101010",
12561 => "0000000011101010",
12562 => "0000000011101010",
12563 => "0000000011101010",
12564 => "0000000011101010",
12565 => "0000000011101010",
12566 => "0000000011101010",
12567 => "0000000011101010",
12568 => "0000000011101010",
12569 => "0000000011101010",
12570 => "0000000011101010",
12571 => "0000000011101010",
12572 => "0000000011101011",
12573 => "0000000011101011",
12574 => "0000000011101011",
12575 => "0000000011101011",
12576 => "0000000011101011",
12577 => "0000000011101011",
12578 => "0000000011101011",
12579 => "0000000011101011",
12580 => "0000000011101011",
12581 => "0000000011101011",
12582 => "0000000011101011",
12583 => "0000000011101011",
12584 => "0000000011101011",
12585 => "0000000011101011",
12586 => "0000000011101011",
12587 => "0000000011101011",
12588 => "0000000011101011",
12589 => "0000000011101011",
12590 => "0000000011101100",
12591 => "0000000011101100",
12592 => "0000000011101100",
12593 => "0000000011101100",
12594 => "0000000011101100",
12595 => "0000000011101100",
12596 => "0000000011101100",
12597 => "0000000011101100",
12598 => "0000000011101100",
12599 => "0000000011101100",
12600 => "0000000011101100",
12601 => "0000000011101100",
12602 => "0000000011101100",
12603 => "0000000011101100",
12604 => "0000000011101100",
12605 => "0000000011101100",
12606 => "0000000011101100",
12607 => "0000000011101101",
12608 => "0000000011101101",
12609 => "0000000011101101",
12610 => "0000000011101101",
12611 => "0000000011101101",
12612 => "0000000011101101",
12613 => "0000000011101101",
12614 => "0000000011101101",
12615 => "0000000011101101",
12616 => "0000000011101101",
12617 => "0000000011101101",
12618 => "0000000011101101",
12619 => "0000000011101101",
12620 => "0000000011101101",
12621 => "0000000011101101",
12622 => "0000000011101101",
12623 => "0000000011101101",
12624 => "0000000011101101",
12625 => "0000000011101110",
12626 => "0000000011101110",
12627 => "0000000011101110",
12628 => "0000000011101110",
12629 => "0000000011101110",
12630 => "0000000011101110",
12631 => "0000000011101110",
12632 => "0000000011101110",
12633 => "0000000011101110",
12634 => "0000000011101110",
12635 => "0000000011101110",
12636 => "0000000011101110",
12637 => "0000000011101110",
12638 => "0000000011101110",
12639 => "0000000011101110",
12640 => "0000000011101110",
12641 => "0000000011101110",
12642 => "0000000011101111",
12643 => "0000000011101111",
12644 => "0000000011101111",
12645 => "0000000011101111",
12646 => "0000000011101111",
12647 => "0000000011101111",
12648 => "0000000011101111",
12649 => "0000000011101111",
12650 => "0000000011101111",
12651 => "0000000011101111",
12652 => "0000000011101111",
12653 => "0000000011101111",
12654 => "0000000011101111",
12655 => "0000000011101111",
12656 => "0000000011101111",
12657 => "0000000011101111",
12658 => "0000000011101111",
12659 => "0000000011110000",
12660 => "0000000011110000",
12661 => "0000000011110000",
12662 => "0000000011110000",
12663 => "0000000011110000",
12664 => "0000000011110000",
12665 => "0000000011110000",
12666 => "0000000011110000",
12667 => "0000000011110000",
12668 => "0000000011110000",
12669 => "0000000011110000",
12670 => "0000000011110000",
12671 => "0000000011110000",
12672 => "0000000011110000",
12673 => "0000000011110000",
12674 => "0000000011110000",
12675 => "0000000011110000",
12676 => "0000000011110001",
12677 => "0000000011110001",
12678 => "0000000011110001",
12679 => "0000000011110001",
12680 => "0000000011110001",
12681 => "0000000011110001",
12682 => "0000000011110001",
12683 => "0000000011110001",
12684 => "0000000011110001",
12685 => "0000000011110001",
12686 => "0000000011110001",
12687 => "0000000011110001",
12688 => "0000000011110001",
12689 => "0000000011110001",
12690 => "0000000011110001",
12691 => "0000000011110001",
12692 => "0000000011110001",
12693 => "0000000011110010",
12694 => "0000000011110010",
12695 => "0000000011110010",
12696 => "0000000011110010",
12697 => "0000000011110010",
12698 => "0000000011110010",
12699 => "0000000011110010",
12700 => "0000000011110010",
12701 => "0000000011110010",
12702 => "0000000011110010",
12703 => "0000000011110010",
12704 => "0000000011110010",
12705 => "0000000011110010",
12706 => "0000000011110010",
12707 => "0000000011110010",
12708 => "0000000011110010",
12709 => "0000000011110010",
12710 => "0000000011110011",
12711 => "0000000011110011",
12712 => "0000000011110011",
12713 => "0000000011110011",
12714 => "0000000011110011",
12715 => "0000000011110011",
12716 => "0000000011110011",
12717 => "0000000011110011",
12718 => "0000000011110011",
12719 => "0000000011110011",
12720 => "0000000011110011",
12721 => "0000000011110011",
12722 => "0000000011110011",
12723 => "0000000011110011",
12724 => "0000000011110011",
12725 => "0000000011110011",
12726 => "0000000011110011",
12727 => "0000000011110100",
12728 => "0000000011110100",
12729 => "0000000011110100",
12730 => "0000000011110100",
12731 => "0000000011110100",
12732 => "0000000011110100",
12733 => "0000000011110100",
12734 => "0000000011110100",
12735 => "0000000011110100",
12736 => "0000000011110100",
12737 => "0000000011110100",
12738 => "0000000011110100",
12739 => "0000000011110100",
12740 => "0000000011110100",
12741 => "0000000011110100",
12742 => "0000000011110100",
12743 => "0000000011110100",
12744 => "0000000011110101",
12745 => "0000000011110101",
12746 => "0000000011110101",
12747 => "0000000011110101",
12748 => "0000000011110101",
12749 => "0000000011110101",
12750 => "0000000011110101",
12751 => "0000000011110101",
12752 => "0000000011110101",
12753 => "0000000011110101",
12754 => "0000000011110101",
12755 => "0000000011110101",
12756 => "0000000011110101",
12757 => "0000000011110101",
12758 => "0000000011110101",
12759 => "0000000011110101",
12760 => "0000000011110101",
12761 => "0000000011110110",
12762 => "0000000011110110",
12763 => "0000000011110110",
12764 => "0000000011110110",
12765 => "0000000011110110",
12766 => "0000000011110110",
12767 => "0000000011110110",
12768 => "0000000011110110",
12769 => "0000000011110110",
12770 => "0000000011110110",
12771 => "0000000011110110",
12772 => "0000000011110110",
12773 => "0000000011110110",
12774 => "0000000011110110",
12775 => "0000000011110110",
12776 => "0000000011110110",
12777 => "0000000011110110",
12778 => "0000000011110111",
12779 => "0000000011110111",
12780 => "0000000011110111",
12781 => "0000000011110111",
12782 => "0000000011110111",
12783 => "0000000011110111",
12784 => "0000000011110111",
12785 => "0000000011110111",
12786 => "0000000011110111",
12787 => "0000000011110111",
12788 => "0000000011110111",
12789 => "0000000011110111",
12790 => "0000000011110111",
12791 => "0000000011110111",
12792 => "0000000011110111",
12793 => "0000000011110111",
12794 => "0000000011111000",
12795 => "0000000011111000",
12796 => "0000000011111000",
12797 => "0000000011111000",
12798 => "0000000011111000",
12799 => "0000000011111000",
12800 => "0000000011111000",
12801 => "0000000011111000",
12802 => "0000000011111000",
12803 => "0000000011111000",
12804 => "0000000011111000",
12805 => "0000000011111000",
12806 => "0000000011111000",
12807 => "0000000011111000",
12808 => "0000000011111000",
12809 => "0000000011111000",
12810 => "0000000011111000",
12811 => "0000000011111001",
12812 => "0000000011111001",
12813 => "0000000011111001",
12814 => "0000000011111001",
12815 => "0000000011111001",
12816 => "0000000011111001",
12817 => "0000000011111001",
12818 => "0000000011111001",
12819 => "0000000011111001",
12820 => "0000000011111001",
12821 => "0000000011111001",
12822 => "0000000011111001",
12823 => "0000000011111001",
12824 => "0000000011111001",
12825 => "0000000011111001",
12826 => "0000000011111001",
12827 => "0000000011111001",
12828 => "0000000011111010",
12829 => "0000000011111010",
12830 => "0000000011111010",
12831 => "0000000011111010",
12832 => "0000000011111010",
12833 => "0000000011111010",
12834 => "0000000011111010",
12835 => "0000000011111010",
12836 => "0000000011111010",
12837 => "0000000011111010",
12838 => "0000000011111010",
12839 => "0000000011111010",
12840 => "0000000011111010",
12841 => "0000000011111010",
12842 => "0000000011111010",
12843 => "0000000011111010",
12844 => "0000000011111011",
12845 => "0000000011111011",
12846 => "0000000011111011",
12847 => "0000000011111011",
12848 => "0000000011111011",
12849 => "0000000011111011",
12850 => "0000000011111011",
12851 => "0000000011111011",
12852 => "0000000011111011",
12853 => "0000000011111011",
12854 => "0000000011111011",
12855 => "0000000011111011",
12856 => "0000000011111011",
12857 => "0000000011111011",
12858 => "0000000011111011",
12859 => "0000000011111011",
12860 => "0000000011111100",
12861 => "0000000011111100",
12862 => "0000000011111100",
12863 => "0000000011111100",
12864 => "0000000011111100",
12865 => "0000000011111100",
12866 => "0000000011111100",
12867 => "0000000011111100",
12868 => "0000000011111100",
12869 => "0000000011111100",
12870 => "0000000011111100",
12871 => "0000000011111100",
12872 => "0000000011111100",
12873 => "0000000011111100",
12874 => "0000000011111100",
12875 => "0000000011111100",
12876 => "0000000011111100",
12877 => "0000000011111101",
12878 => "0000000011111101",
12879 => "0000000011111101",
12880 => "0000000011111101",
12881 => "0000000011111101",
12882 => "0000000011111101",
12883 => "0000000011111101",
12884 => "0000000011111101",
12885 => "0000000011111101",
12886 => "0000000011111101",
12887 => "0000000011111101",
12888 => "0000000011111101",
12889 => "0000000011111101",
12890 => "0000000011111101",
12891 => "0000000011111101",
12892 => "0000000011111101",
12893 => "0000000011111110",
12894 => "0000000011111110",
12895 => "0000000011111110",
12896 => "0000000011111110",
12897 => "0000000011111110",
12898 => "0000000011111110",
12899 => "0000000011111110",
12900 => "0000000011111110",
12901 => "0000000011111110",
12902 => "0000000011111110",
12903 => "0000000011111110",
12904 => "0000000011111110",
12905 => "0000000011111110",
12906 => "0000000011111110",
12907 => "0000000011111110",
12908 => "0000000011111110",
12909 => "0000000011111111",
12910 => "0000000011111111",
12911 => "0000000011111111",
12912 => "0000000011111111",
12913 => "0000000011111111",
12914 => "0000000011111111",
12915 => "0000000011111111",
12916 => "0000000011111111",
12917 => "0000000011111111",
12918 => "0000000011111111",
12919 => "0000000011111111",
12920 => "0000000011111111",
12921 => "0000000011111111",
12922 => "0000000011111111",
12923 => "0000000011111111",
12924 => "0000000011111111",
12925 => "0000000011111111",
12926 => "0000000100000000",
12927 => "0000000100000000",
12928 => "0000000100000000",
12929 => "0000000100000000",
12930 => "0000000100000000",
12931 => "0000000100000000",
12932 => "0000000100000000",
12933 => "0000000100000000",
12934 => "0000000100000000",
12935 => "0000000100000000",
12936 => "0000000100000000",
12937 => "0000000100000000",
12938 => "0000000100000000",
12939 => "0000000100000000",
12940 => "0000000100000000",
12941 => "0000000100000001",
12942 => "0000000100000001",
12943 => "0000000100000001",
12944 => "0000000100000001",
12945 => "0000000100000001",
12946 => "0000000100000001",
12947 => "0000000100000001",
12948 => "0000000100000001",
12949 => "0000000100000001",
12950 => "0000000100000001",
12951 => "0000000100000001",
12952 => "0000000100000001",
12953 => "0000000100000001",
12954 => "0000000100000001",
12955 => "0000000100000001",
12956 => "0000000100000001",
12957 => "0000000100000010",
12958 => "0000000100000010",
12959 => "0000000100000010",
12960 => "0000000100000010",
12961 => "0000000100000010",
12962 => "0000000100000010",
12963 => "0000000100000010",
12964 => "0000000100000010",
12965 => "0000000100000010",
12966 => "0000000100000010",
12967 => "0000000100000010",
12968 => "0000000100000010",
12969 => "0000000100000010",
12970 => "0000000100000010",
12971 => "0000000100000010",
12972 => "0000000100000010",
12973 => "0000000100000011",
12974 => "0000000100000011",
12975 => "0000000100000011",
12976 => "0000000100000011",
12977 => "0000000100000011",
12978 => "0000000100000011",
12979 => "0000000100000011",
12980 => "0000000100000011",
12981 => "0000000100000011",
12982 => "0000000100000011",
12983 => "0000000100000011",
12984 => "0000000100000011",
12985 => "0000000100000011",
12986 => "0000000100000011",
12987 => "0000000100000011",
12988 => "0000000100000011",
12989 => "0000000100000100",
12990 => "0000000100000100",
12991 => "0000000100000100",
12992 => "0000000100000100",
12993 => "0000000100000100",
12994 => "0000000100000100",
12995 => "0000000100000100",
12996 => "0000000100000100",
12997 => "0000000100000100",
12998 => "0000000100000100",
12999 => "0000000100000100",
13000 => "0000000100000100",
13001 => "0000000100000100",
13002 => "0000000100000100",
13003 => "0000000100000100",
13004 => "0000000100000101",
13005 => "0000000100000101",
13006 => "0000000100000101",
13007 => "0000000100000101",
13008 => "0000000100000101",
13009 => "0000000100000101",
13010 => "0000000100000101",
13011 => "0000000100000101",
13012 => "0000000100000101",
13013 => "0000000100000101",
13014 => "0000000100000101",
13015 => "0000000100000101",
13016 => "0000000100000101",
13017 => "0000000100000101",
13018 => "0000000100000101",
13019 => "0000000100000101",
13020 => "0000000100000110",
13021 => "0000000100000110",
13022 => "0000000100000110",
13023 => "0000000100000110",
13024 => "0000000100000110",
13025 => "0000000100000110",
13026 => "0000000100000110",
13027 => "0000000100000110",
13028 => "0000000100000110",
13029 => "0000000100000110",
13030 => "0000000100000110",
13031 => "0000000100000110",
13032 => "0000000100000110",
13033 => "0000000100000110",
13034 => "0000000100000110",
13035 => "0000000100000110",
13036 => "0000000100000111",
13037 => "0000000100000111",
13038 => "0000000100000111",
13039 => "0000000100000111",
13040 => "0000000100000111",
13041 => "0000000100000111",
13042 => "0000000100000111",
13043 => "0000000100000111",
13044 => "0000000100000111",
13045 => "0000000100000111",
13046 => "0000000100000111",
13047 => "0000000100000111",
13048 => "0000000100000111",
13049 => "0000000100000111",
13050 => "0000000100000111",
13051 => "0000000100000111",
13052 => "0000000100001000",
13053 => "0000000100001000",
13054 => "0000000100001000",
13055 => "0000000100001000",
13056 => "0000000100001000",
13057 => "0000000100001000",
13058 => "0000000100001000",
13059 => "0000000100001000",
13060 => "0000000100001000",
13061 => "0000000100001000",
13062 => "0000000100001000",
13063 => "0000000100001000",
13064 => "0000000100001000",
13065 => "0000000100001000",
13066 => "0000000100001000",
13067 => "0000000100001001",
13068 => "0000000100001001",
13069 => "0000000100001001",
13070 => "0000000100001001",
13071 => "0000000100001001",
13072 => "0000000100001001",
13073 => "0000000100001001",
13074 => "0000000100001001",
13075 => "0000000100001001",
13076 => "0000000100001001",
13077 => "0000000100001001",
13078 => "0000000100001001",
13079 => "0000000100001001",
13080 => "0000000100001001",
13081 => "0000000100001001",
13082 => "0000000100001001",
13083 => "0000000100001010",
13084 => "0000000100001010",
13085 => "0000000100001010",
13086 => "0000000100001010",
13087 => "0000000100001010",
13088 => "0000000100001010",
13089 => "0000000100001010",
13090 => "0000000100001010",
13091 => "0000000100001010",
13092 => "0000000100001010",
13093 => "0000000100001010",
13094 => "0000000100001010",
13095 => "0000000100001010",
13096 => "0000000100001010",
13097 => "0000000100001010",
13098 => "0000000100001011",
13099 => "0000000100001011",
13100 => "0000000100001011",
13101 => "0000000100001011",
13102 => "0000000100001011",
13103 => "0000000100001011",
13104 => "0000000100001011",
13105 => "0000000100001011",
13106 => "0000000100001011",
13107 => "0000000100001011",
13108 => "0000000100001011",
13109 => "0000000100001011",
13110 => "0000000100001011",
13111 => "0000000100001011",
13112 => "0000000100001011",
13113 => "0000000100001011",
13114 => "0000000100001100",
13115 => "0000000100001100",
13116 => "0000000100001100",
13117 => "0000000100001100",
13118 => "0000000100001100",
13119 => "0000000100001100",
13120 => "0000000100001100",
13121 => "0000000100001100",
13122 => "0000000100001100",
13123 => "0000000100001100",
13124 => "0000000100001100",
13125 => "0000000100001100",
13126 => "0000000100001100",
13127 => "0000000100001100",
13128 => "0000000100001100",
13129 => "0000000100001101",
13130 => "0000000100001101",
13131 => "0000000100001101",
13132 => "0000000100001101",
13133 => "0000000100001101",
13134 => "0000000100001101",
13135 => "0000000100001101",
13136 => "0000000100001101",
13137 => "0000000100001101",
13138 => "0000000100001101",
13139 => "0000000100001101",
13140 => "0000000100001101",
13141 => "0000000100001101",
13142 => "0000000100001101",
13143 => "0000000100001101",
13144 => "0000000100001110",
13145 => "0000000100001110",
13146 => "0000000100001110",
13147 => "0000000100001110",
13148 => "0000000100001110",
13149 => "0000000100001110",
13150 => "0000000100001110",
13151 => "0000000100001110",
13152 => "0000000100001110",
13153 => "0000000100001110",
13154 => "0000000100001110",
13155 => "0000000100001110",
13156 => "0000000100001110",
13157 => "0000000100001110",
13158 => "0000000100001110",
13159 => "0000000100001110",
13160 => "0000000100001111",
13161 => "0000000100001111",
13162 => "0000000100001111",
13163 => "0000000100001111",
13164 => "0000000100001111",
13165 => "0000000100001111",
13166 => "0000000100001111",
13167 => "0000000100001111",
13168 => "0000000100001111",
13169 => "0000000100001111",
13170 => "0000000100001111",
13171 => "0000000100001111",
13172 => "0000000100001111",
13173 => "0000000100001111",
13174 => "0000000100001111",
13175 => "0000000100010000",
13176 => "0000000100010000",
13177 => "0000000100010000",
13178 => "0000000100010000",
13179 => "0000000100010000",
13180 => "0000000100010000",
13181 => "0000000100010000",
13182 => "0000000100010000",
13183 => "0000000100010000",
13184 => "0000000100010000",
13185 => "0000000100010000",
13186 => "0000000100010000",
13187 => "0000000100010000",
13188 => "0000000100010000",
13189 => "0000000100010000",
13190 => "0000000100010001",
13191 => "0000000100010001",
13192 => "0000000100010001",
13193 => "0000000100010001",
13194 => "0000000100010001",
13195 => "0000000100010001",
13196 => "0000000100010001",
13197 => "0000000100010001",
13198 => "0000000100010001",
13199 => "0000000100010001",
13200 => "0000000100010001",
13201 => "0000000100010001",
13202 => "0000000100010001",
13203 => "0000000100010001",
13204 => "0000000100010001",
13205 => "0000000100010010",
13206 => "0000000100010010",
13207 => "0000000100010010",
13208 => "0000000100010010",
13209 => "0000000100010010",
13210 => "0000000100010010",
13211 => "0000000100010010",
13212 => "0000000100010010",
13213 => "0000000100010010",
13214 => "0000000100010010",
13215 => "0000000100010010",
13216 => "0000000100010010",
13217 => "0000000100010010",
13218 => "0000000100010010",
13219 => "0000000100010010",
13220 => "0000000100010011",
13221 => "0000000100010011",
13222 => "0000000100010011",
13223 => "0000000100010011",
13224 => "0000000100010011",
13225 => "0000000100010011",
13226 => "0000000100010011",
13227 => "0000000100010011",
13228 => "0000000100010011",
13229 => "0000000100010011",
13230 => "0000000100010011",
13231 => "0000000100010011",
13232 => "0000000100010011",
13233 => "0000000100010011",
13234 => "0000000100010011",
13235 => "0000000100010100",
13236 => "0000000100010100",
13237 => "0000000100010100",
13238 => "0000000100010100",
13239 => "0000000100010100",
13240 => "0000000100010100",
13241 => "0000000100010100",
13242 => "0000000100010100",
13243 => "0000000100010100",
13244 => "0000000100010100",
13245 => "0000000100010100",
13246 => "0000000100010100",
13247 => "0000000100010100",
13248 => "0000000100010100",
13249 => "0000000100010100",
13250 => "0000000100010101",
13251 => "0000000100010101",
13252 => "0000000100010101",
13253 => "0000000100010101",
13254 => "0000000100010101",
13255 => "0000000100010101",
13256 => "0000000100010101",
13257 => "0000000100010101",
13258 => "0000000100010101",
13259 => "0000000100010101",
13260 => "0000000100010101",
13261 => "0000000100010101",
13262 => "0000000100010101",
13263 => "0000000100010101",
13264 => "0000000100010101",
13265 => "0000000100010110",
13266 => "0000000100010110",
13267 => "0000000100010110",
13268 => "0000000100010110",
13269 => "0000000100010110",
13270 => "0000000100010110",
13271 => "0000000100010110",
13272 => "0000000100010110",
13273 => "0000000100010110",
13274 => "0000000100010110",
13275 => "0000000100010110",
13276 => "0000000100010110",
13277 => "0000000100010110",
13278 => "0000000100010110",
13279 => "0000000100010110",
13280 => "0000000100010111",
13281 => "0000000100010111",
13282 => "0000000100010111",
13283 => "0000000100010111",
13284 => "0000000100010111",
13285 => "0000000100010111",
13286 => "0000000100010111",
13287 => "0000000100010111",
13288 => "0000000100010111",
13289 => "0000000100010111",
13290 => "0000000100010111",
13291 => "0000000100010111",
13292 => "0000000100010111",
13293 => "0000000100010111",
13294 => "0000000100010111",
13295 => "0000000100011000",
13296 => "0000000100011000",
13297 => "0000000100011000",
13298 => "0000000100011000",
13299 => "0000000100011000",
13300 => "0000000100011000",
13301 => "0000000100011000",
13302 => "0000000100011000",
13303 => "0000000100011000",
13304 => "0000000100011000",
13305 => "0000000100011000",
13306 => "0000000100011000",
13307 => "0000000100011000",
13308 => "0000000100011000",
13309 => "0000000100011001",
13310 => "0000000100011001",
13311 => "0000000100011001",
13312 => "0000000100011001",
13313 => "0000000100011001",
13314 => "0000000100011001",
13315 => "0000000100011001",
13316 => "0000000100011001",
13317 => "0000000100011001",
13318 => "0000000100011001",
13319 => "0000000100011001",
13320 => "0000000100011001",
13321 => "0000000100011001",
13322 => "0000000100011001",
13323 => "0000000100011001",
13324 => "0000000100011010",
13325 => "0000000100011010",
13326 => "0000000100011010",
13327 => "0000000100011010",
13328 => "0000000100011010",
13329 => "0000000100011010",
13330 => "0000000100011010",
13331 => "0000000100011010",
13332 => "0000000100011010",
13333 => "0000000100011010",
13334 => "0000000100011010",
13335 => "0000000100011010",
13336 => "0000000100011010",
13337 => "0000000100011010",
13338 => "0000000100011010",
13339 => "0000000100011011",
13340 => "0000000100011011",
13341 => "0000000100011011",
13342 => "0000000100011011",
13343 => "0000000100011011",
13344 => "0000000100011011",
13345 => "0000000100011011",
13346 => "0000000100011011",
13347 => "0000000100011011",
13348 => "0000000100011011",
13349 => "0000000100011011",
13350 => "0000000100011011",
13351 => "0000000100011011",
13352 => "0000000100011011",
13353 => "0000000100011100",
13354 => "0000000100011100",
13355 => "0000000100011100",
13356 => "0000000100011100",
13357 => "0000000100011100",
13358 => "0000000100011100",
13359 => "0000000100011100",
13360 => "0000000100011100",
13361 => "0000000100011100",
13362 => "0000000100011100",
13363 => "0000000100011100",
13364 => "0000000100011100",
13365 => "0000000100011100",
13366 => "0000000100011100",
13367 => "0000000100011100",
13368 => "0000000100011101",
13369 => "0000000100011101",
13370 => "0000000100011101",
13371 => "0000000100011101",
13372 => "0000000100011101",
13373 => "0000000100011101",
13374 => "0000000100011101",
13375 => "0000000100011101",
13376 => "0000000100011101",
13377 => "0000000100011101",
13378 => "0000000100011101",
13379 => "0000000100011101",
13380 => "0000000100011101",
13381 => "0000000100011101",
13382 => "0000000100011110",
13383 => "0000000100011110",
13384 => "0000000100011110",
13385 => "0000000100011110",
13386 => "0000000100011110",
13387 => "0000000100011110",
13388 => "0000000100011110",
13389 => "0000000100011110",
13390 => "0000000100011110",
13391 => "0000000100011110",
13392 => "0000000100011110",
13393 => "0000000100011110",
13394 => "0000000100011110",
13395 => "0000000100011110",
13396 => "0000000100011110",
13397 => "0000000100011111",
13398 => "0000000100011111",
13399 => "0000000100011111",
13400 => "0000000100011111",
13401 => "0000000100011111",
13402 => "0000000100011111",
13403 => "0000000100011111",
13404 => "0000000100011111",
13405 => "0000000100011111",
13406 => "0000000100011111",
13407 => "0000000100011111",
13408 => "0000000100011111",
13409 => "0000000100011111",
13410 => "0000000100011111",
13411 => "0000000100100000",
13412 => "0000000100100000",
13413 => "0000000100100000",
13414 => "0000000100100000",
13415 => "0000000100100000",
13416 => "0000000100100000",
13417 => "0000000100100000",
13418 => "0000000100100000",
13419 => "0000000100100000",
13420 => "0000000100100000",
13421 => "0000000100100000",
13422 => "0000000100100000",
13423 => "0000000100100000",
13424 => "0000000100100000",
13425 => "0000000100100000",
13426 => "0000000100100001",
13427 => "0000000100100001",
13428 => "0000000100100001",
13429 => "0000000100100001",
13430 => "0000000100100001",
13431 => "0000000100100001",
13432 => "0000000100100001",
13433 => "0000000100100001",
13434 => "0000000100100001",
13435 => "0000000100100001",
13436 => "0000000100100001",
13437 => "0000000100100001",
13438 => "0000000100100001",
13439 => "0000000100100001",
13440 => "0000000100100010",
13441 => "0000000100100010",
13442 => "0000000100100010",
13443 => "0000000100100010",
13444 => "0000000100100010",
13445 => "0000000100100010",
13446 => "0000000100100010",
13447 => "0000000100100010",
13448 => "0000000100100010",
13449 => "0000000100100010",
13450 => "0000000100100010",
13451 => "0000000100100010",
13452 => "0000000100100010",
13453 => "0000000100100010",
13454 => "0000000100100011",
13455 => "0000000100100011",
13456 => "0000000100100011",
13457 => "0000000100100011",
13458 => "0000000100100011",
13459 => "0000000100100011",
13460 => "0000000100100011",
13461 => "0000000100100011",
13462 => "0000000100100011",
13463 => "0000000100100011",
13464 => "0000000100100011",
13465 => "0000000100100011",
13466 => "0000000100100011",
13467 => "0000000100100011",
13468 => "0000000100100100",
13469 => "0000000100100100",
13470 => "0000000100100100",
13471 => "0000000100100100",
13472 => "0000000100100100",
13473 => "0000000100100100",
13474 => "0000000100100100",
13475 => "0000000100100100",
13476 => "0000000100100100",
13477 => "0000000100100100",
13478 => "0000000100100100",
13479 => "0000000100100100",
13480 => "0000000100100100",
13481 => "0000000100100100",
13482 => "0000000100100101",
13483 => "0000000100100101",
13484 => "0000000100100101",
13485 => "0000000100100101",
13486 => "0000000100100101",
13487 => "0000000100100101",
13488 => "0000000100100101",
13489 => "0000000100100101",
13490 => "0000000100100101",
13491 => "0000000100100101",
13492 => "0000000100100101",
13493 => "0000000100100101",
13494 => "0000000100100101",
13495 => "0000000100100101",
13496 => "0000000100100110",
13497 => "0000000100100110",
13498 => "0000000100100110",
13499 => "0000000100100110",
13500 => "0000000100100110",
13501 => "0000000100100110",
13502 => "0000000100100110",
13503 => "0000000100100110",
13504 => "0000000100100110",
13505 => "0000000100100110",
13506 => "0000000100100110",
13507 => "0000000100100110",
13508 => "0000000100100110",
13509 => "0000000100100110",
13510 => "0000000100100111",
13511 => "0000000100100111",
13512 => "0000000100100111",
13513 => "0000000100100111",
13514 => "0000000100100111",
13515 => "0000000100100111",
13516 => "0000000100100111",
13517 => "0000000100100111",
13518 => "0000000100100111",
13519 => "0000000100100111",
13520 => "0000000100100111",
13521 => "0000000100100111",
13522 => "0000000100100111",
13523 => "0000000100100111",
13524 => "0000000100101000",
13525 => "0000000100101000",
13526 => "0000000100101000",
13527 => "0000000100101000",
13528 => "0000000100101000",
13529 => "0000000100101000",
13530 => "0000000100101000",
13531 => "0000000100101000",
13532 => "0000000100101000",
13533 => "0000000100101000",
13534 => "0000000100101000",
13535 => "0000000100101000",
13536 => "0000000100101000",
13537 => "0000000100101000",
13538 => "0000000100101001",
13539 => "0000000100101001",
13540 => "0000000100101001",
13541 => "0000000100101001",
13542 => "0000000100101001",
13543 => "0000000100101001",
13544 => "0000000100101001",
13545 => "0000000100101001",
13546 => "0000000100101001",
13547 => "0000000100101001",
13548 => "0000000100101001",
13549 => "0000000100101001",
13550 => "0000000100101001",
13551 => "0000000100101001",
13552 => "0000000100101010",
13553 => "0000000100101010",
13554 => "0000000100101010",
13555 => "0000000100101010",
13556 => "0000000100101010",
13557 => "0000000100101010",
13558 => "0000000100101010",
13559 => "0000000100101010",
13560 => "0000000100101010",
13561 => "0000000100101010",
13562 => "0000000100101010",
13563 => "0000000100101010",
13564 => "0000000100101010",
13565 => "0000000100101010",
13566 => "0000000100101011",
13567 => "0000000100101011",
13568 => "0000000100101011",
13569 => "0000000100101011",
13570 => "0000000100101011",
13571 => "0000000100101011",
13572 => "0000000100101011",
13573 => "0000000100101011",
13574 => "0000000100101011",
13575 => "0000000100101011",
13576 => "0000000100101011",
13577 => "0000000100101011",
13578 => "0000000100101011",
13579 => "0000000100101011",
13580 => "0000000100101100",
13581 => "0000000100101100",
13582 => "0000000100101100",
13583 => "0000000100101100",
13584 => "0000000100101100",
13585 => "0000000100101100",
13586 => "0000000100101100",
13587 => "0000000100101100",
13588 => "0000000100101100",
13589 => "0000000100101100",
13590 => "0000000100101100",
13591 => "0000000100101100",
13592 => "0000000100101100",
13593 => "0000000100101100",
13594 => "0000000100101101",
13595 => "0000000100101101",
13596 => "0000000100101101",
13597 => "0000000100101101",
13598 => "0000000100101101",
13599 => "0000000100101101",
13600 => "0000000100101101",
13601 => "0000000100101101",
13602 => "0000000100101101",
13603 => "0000000100101101",
13604 => "0000000100101101",
13605 => "0000000100101101",
13606 => "0000000100101101",
13607 => "0000000100101110",
13608 => "0000000100101110",
13609 => "0000000100101110",
13610 => "0000000100101110",
13611 => "0000000100101110",
13612 => "0000000100101110",
13613 => "0000000100101110",
13614 => "0000000100101110",
13615 => "0000000100101110",
13616 => "0000000100101110",
13617 => "0000000100101110",
13618 => "0000000100101110",
13619 => "0000000100101110",
13620 => "0000000100101110",
13621 => "0000000100101111",
13622 => "0000000100101111",
13623 => "0000000100101111",
13624 => "0000000100101111",
13625 => "0000000100101111",
13626 => "0000000100101111",
13627 => "0000000100101111",
13628 => "0000000100101111",
13629 => "0000000100101111",
13630 => "0000000100101111",
13631 => "0000000100101111",
13632 => "0000000100101111",
13633 => "0000000100101111",
13634 => "0000000100101111",
13635 => "0000000100110000",
13636 => "0000000100110000",
13637 => "0000000100110000",
13638 => "0000000100110000",
13639 => "0000000100110000",
13640 => "0000000100110000",
13641 => "0000000100110000",
13642 => "0000000100110000",
13643 => "0000000100110000",
13644 => "0000000100110000",
13645 => "0000000100110000",
13646 => "0000000100110000",
13647 => "0000000100110000",
13648 => "0000000100110001",
13649 => "0000000100110001",
13650 => "0000000100110001",
13651 => "0000000100110001",
13652 => "0000000100110001",
13653 => "0000000100110001",
13654 => "0000000100110001",
13655 => "0000000100110001",
13656 => "0000000100110001",
13657 => "0000000100110001",
13658 => "0000000100110001",
13659 => "0000000100110001",
13660 => "0000000100110001",
13661 => "0000000100110001",
13662 => "0000000100110010",
13663 => "0000000100110010",
13664 => "0000000100110010",
13665 => "0000000100110010",
13666 => "0000000100110010",
13667 => "0000000100110010",
13668 => "0000000100110010",
13669 => "0000000100110010",
13670 => "0000000100110010",
13671 => "0000000100110010",
13672 => "0000000100110010",
13673 => "0000000100110010",
13674 => "0000000100110010",
13675 => "0000000100110011",
13676 => "0000000100110011",
13677 => "0000000100110011",
13678 => "0000000100110011",
13679 => "0000000100110011",
13680 => "0000000100110011",
13681 => "0000000100110011",
13682 => "0000000100110011",
13683 => "0000000100110011",
13684 => "0000000100110011",
13685 => "0000000100110011",
13686 => "0000000100110011",
13687 => "0000000100110011",
13688 => "0000000100110011",
13689 => "0000000100110100",
13690 => "0000000100110100",
13691 => "0000000100110100",
13692 => "0000000100110100",
13693 => "0000000100110100",
13694 => "0000000100110100",
13695 => "0000000100110100",
13696 => "0000000100110100",
13697 => "0000000100110100",
13698 => "0000000100110100",
13699 => "0000000100110100",
13700 => "0000000100110100",
13701 => "0000000100110100",
13702 => "0000000100110101",
13703 => "0000000100110101",
13704 => "0000000100110101",
13705 => "0000000100110101",
13706 => "0000000100110101",
13707 => "0000000100110101",
13708 => "0000000100110101",
13709 => "0000000100110101",
13710 => "0000000100110101",
13711 => "0000000100110101",
13712 => "0000000100110101",
13713 => "0000000100110101",
13714 => "0000000100110101",
13715 => "0000000100110101",
13716 => "0000000100110110",
13717 => "0000000100110110",
13718 => "0000000100110110",
13719 => "0000000100110110",
13720 => "0000000100110110",
13721 => "0000000100110110",
13722 => "0000000100110110",
13723 => "0000000100110110",
13724 => "0000000100110110",
13725 => "0000000100110110",
13726 => "0000000100110110",
13727 => "0000000100110110",
13728 => "0000000100110110",
13729 => "0000000100110111",
13730 => "0000000100110111",
13731 => "0000000100110111",
13732 => "0000000100110111",
13733 => "0000000100110111",
13734 => "0000000100110111",
13735 => "0000000100110111",
13736 => "0000000100110111",
13737 => "0000000100110111",
13738 => "0000000100110111",
13739 => "0000000100110111",
13740 => "0000000100110111",
13741 => "0000000100110111",
13742 => "0000000100111000",
13743 => "0000000100111000",
13744 => "0000000100111000",
13745 => "0000000100111000",
13746 => "0000000100111000",
13747 => "0000000100111000",
13748 => "0000000100111000",
13749 => "0000000100111000",
13750 => "0000000100111000",
13751 => "0000000100111000",
13752 => "0000000100111000",
13753 => "0000000100111000",
13754 => "0000000100111000",
13755 => "0000000100111001",
13756 => "0000000100111001",
13757 => "0000000100111001",
13758 => "0000000100111001",
13759 => "0000000100111001",
13760 => "0000000100111001",
13761 => "0000000100111001",
13762 => "0000000100111001",
13763 => "0000000100111001",
13764 => "0000000100111001",
13765 => "0000000100111001",
13766 => "0000000100111001",
13767 => "0000000100111001",
13768 => "0000000100111001",
13769 => "0000000100111010",
13770 => "0000000100111010",
13771 => "0000000100111010",
13772 => "0000000100111010",
13773 => "0000000100111010",
13774 => "0000000100111010",
13775 => "0000000100111010",
13776 => "0000000100111010",
13777 => "0000000100111010",
13778 => "0000000100111010",
13779 => "0000000100111010",
13780 => "0000000100111010",
13781 => "0000000100111010",
13782 => "0000000100111011",
13783 => "0000000100111011",
13784 => "0000000100111011",
13785 => "0000000100111011",
13786 => "0000000100111011",
13787 => "0000000100111011",
13788 => "0000000100111011",
13789 => "0000000100111011",
13790 => "0000000100111011",
13791 => "0000000100111011",
13792 => "0000000100111011",
13793 => "0000000100111011",
13794 => "0000000100111011",
13795 => "0000000100111100",
13796 => "0000000100111100",
13797 => "0000000100111100",
13798 => "0000000100111100",
13799 => "0000000100111100",
13800 => "0000000100111100",
13801 => "0000000100111100",
13802 => "0000000100111100",
13803 => "0000000100111100",
13804 => "0000000100111100",
13805 => "0000000100111100",
13806 => "0000000100111100",
13807 => "0000000100111100",
13808 => "0000000100111101",
13809 => "0000000100111101",
13810 => "0000000100111101",
13811 => "0000000100111101",
13812 => "0000000100111101",
13813 => "0000000100111101",
13814 => "0000000100111101",
13815 => "0000000100111101",
13816 => "0000000100111101",
13817 => "0000000100111101",
13818 => "0000000100111101",
13819 => "0000000100111101",
13820 => "0000000100111101",
13821 => "0000000100111110",
13822 => "0000000100111110",
13823 => "0000000100111110",
13824 => "0000000100111110",
13825 => "0000000100111110",
13826 => "0000000100111110",
13827 => "0000000100111110",
13828 => "0000000100111110",
13829 => "0000000100111110",
13830 => "0000000100111110",
13831 => "0000000100111110",
13832 => "0000000100111110",
13833 => "0000000100111110",
13834 => "0000000100111111",
13835 => "0000000100111111",
13836 => "0000000100111111",
13837 => "0000000100111111",
13838 => "0000000100111111",
13839 => "0000000100111111",
13840 => "0000000100111111",
13841 => "0000000100111111",
13842 => "0000000100111111",
13843 => "0000000100111111",
13844 => "0000000100111111",
13845 => "0000000100111111",
13846 => "0000000100111111",
13847 => "0000000101000000",
13848 => "0000000101000000",
13849 => "0000000101000000",
13850 => "0000000101000000",
13851 => "0000000101000000",
13852 => "0000000101000000",
13853 => "0000000101000000",
13854 => "0000000101000000",
13855 => "0000000101000000",
13856 => "0000000101000000",
13857 => "0000000101000000",
13858 => "0000000101000000",
13859 => "0000000101000000",
13860 => "0000000101000001",
13861 => "0000000101000001",
13862 => "0000000101000001",
13863 => "0000000101000001",
13864 => "0000000101000001",
13865 => "0000000101000001",
13866 => "0000000101000001",
13867 => "0000000101000001",
13868 => "0000000101000001",
13869 => "0000000101000001",
13870 => "0000000101000001",
13871 => "0000000101000001",
13872 => "0000000101000001",
13873 => "0000000101000010",
13874 => "0000000101000010",
13875 => "0000000101000010",
13876 => "0000000101000010",
13877 => "0000000101000010",
13878 => "0000000101000010",
13879 => "0000000101000010",
13880 => "0000000101000010",
13881 => "0000000101000010",
13882 => "0000000101000010",
13883 => "0000000101000010",
13884 => "0000000101000010",
13885 => "0000000101000010",
13886 => "0000000101000011",
13887 => "0000000101000011",
13888 => "0000000101000011",
13889 => "0000000101000011",
13890 => "0000000101000011",
13891 => "0000000101000011",
13892 => "0000000101000011",
13893 => "0000000101000011",
13894 => "0000000101000011",
13895 => "0000000101000011",
13896 => "0000000101000011",
13897 => "0000000101000011",
13898 => "0000000101000100",
13899 => "0000000101000100",
13900 => "0000000101000100",
13901 => "0000000101000100",
13902 => "0000000101000100",
13903 => "0000000101000100",
13904 => "0000000101000100",
13905 => "0000000101000100",
13906 => "0000000101000100",
13907 => "0000000101000100",
13908 => "0000000101000100",
13909 => "0000000101000100",
13910 => "0000000101000100",
13911 => "0000000101000101",
13912 => "0000000101000101",
13913 => "0000000101000101",
13914 => "0000000101000101",
13915 => "0000000101000101",
13916 => "0000000101000101",
13917 => "0000000101000101",
13918 => "0000000101000101",
13919 => "0000000101000101",
13920 => "0000000101000101",
13921 => "0000000101000101",
13922 => "0000000101000101",
13923 => "0000000101000101",
13924 => "0000000101000110",
13925 => "0000000101000110",
13926 => "0000000101000110",
13927 => "0000000101000110",
13928 => "0000000101000110",
13929 => "0000000101000110",
13930 => "0000000101000110",
13931 => "0000000101000110",
13932 => "0000000101000110",
13933 => "0000000101000110",
13934 => "0000000101000110",
13935 => "0000000101000110",
13936 => "0000000101000111",
13937 => "0000000101000111",
13938 => "0000000101000111",
13939 => "0000000101000111",
13940 => "0000000101000111",
13941 => "0000000101000111",
13942 => "0000000101000111",
13943 => "0000000101000111",
13944 => "0000000101000111",
13945 => "0000000101000111",
13946 => "0000000101000111",
13947 => "0000000101000111",
13948 => "0000000101000111",
13949 => "0000000101001000",
13950 => "0000000101001000",
13951 => "0000000101001000",
13952 => "0000000101001000",
13953 => "0000000101001000",
13954 => "0000000101001000",
13955 => "0000000101001000",
13956 => "0000000101001000",
13957 => "0000000101001000",
13958 => "0000000101001000",
13959 => "0000000101001000",
13960 => "0000000101001000",
13961 => "0000000101001000",
13962 => "0000000101001001",
13963 => "0000000101001001",
13964 => "0000000101001001",
13965 => "0000000101001001",
13966 => "0000000101001001",
13967 => "0000000101001001",
13968 => "0000000101001001",
13969 => "0000000101001001",
13970 => "0000000101001001",
13971 => "0000000101001001",
13972 => "0000000101001001",
13973 => "0000000101001001",
13974 => "0000000101001010",
13975 => "0000000101001010",
13976 => "0000000101001010",
13977 => "0000000101001010",
13978 => "0000000101001010",
13979 => "0000000101001010",
13980 => "0000000101001010",
13981 => "0000000101001010",
13982 => "0000000101001010",
13983 => "0000000101001010",
13984 => "0000000101001010",
13985 => "0000000101001010",
13986 => "0000000101001010",
13987 => "0000000101001011",
13988 => "0000000101001011",
13989 => "0000000101001011",
13990 => "0000000101001011",
13991 => "0000000101001011",
13992 => "0000000101001011",
13993 => "0000000101001011",
13994 => "0000000101001011",
13995 => "0000000101001011",
13996 => "0000000101001011",
13997 => "0000000101001011",
13998 => "0000000101001011",
13999 => "0000000101001100",
14000 => "0000000101001100",
14001 => "0000000101001100",
14002 => "0000000101001100",
14003 => "0000000101001100",
14004 => "0000000101001100",
14005 => "0000000101001100",
14006 => "0000000101001100",
14007 => "0000000101001100",
14008 => "0000000101001100",
14009 => "0000000101001100",
14010 => "0000000101001100",
14011 => "0000000101001100",
14012 => "0000000101001101",
14013 => "0000000101001101",
14014 => "0000000101001101",
14015 => "0000000101001101",
14016 => "0000000101001101",
14017 => "0000000101001101",
14018 => "0000000101001101",
14019 => "0000000101001101",
14020 => "0000000101001101",
14021 => "0000000101001101",
14022 => "0000000101001101",
14023 => "0000000101001101",
14024 => "0000000101001110",
14025 => "0000000101001110",
14026 => "0000000101001110",
14027 => "0000000101001110",
14028 => "0000000101001110",
14029 => "0000000101001110",
14030 => "0000000101001110",
14031 => "0000000101001110",
14032 => "0000000101001110",
14033 => "0000000101001110",
14034 => "0000000101001110",
14035 => "0000000101001110",
14036 => "0000000101001110",
14037 => "0000000101001111",
14038 => "0000000101001111",
14039 => "0000000101001111",
14040 => "0000000101001111",
14041 => "0000000101001111",
14042 => "0000000101001111",
14043 => "0000000101001111",
14044 => "0000000101001111",
14045 => "0000000101001111",
14046 => "0000000101001111",
14047 => "0000000101001111",
14048 => "0000000101001111",
14049 => "0000000101010000",
14050 => "0000000101010000",
14051 => "0000000101010000",
14052 => "0000000101010000",
14053 => "0000000101010000",
14054 => "0000000101010000",
14055 => "0000000101010000",
14056 => "0000000101010000",
14057 => "0000000101010000",
14058 => "0000000101010000",
14059 => "0000000101010000",
14060 => "0000000101010000",
14061 => "0000000101010001",
14062 => "0000000101010001",
14063 => "0000000101010001",
14064 => "0000000101010001",
14065 => "0000000101010001",
14066 => "0000000101010001",
14067 => "0000000101010001",
14068 => "0000000101010001",
14069 => "0000000101010001",
14070 => "0000000101010001",
14071 => "0000000101010001",
14072 => "0000000101010001",
14073 => "0000000101010010",
14074 => "0000000101010010",
14075 => "0000000101010010",
14076 => "0000000101010010",
14077 => "0000000101010010",
14078 => "0000000101010010",
14079 => "0000000101010010",
14080 => "0000000101010010",
14081 => "0000000101010010",
14082 => "0000000101010010",
14083 => "0000000101010010",
14084 => "0000000101010010",
14085 => "0000000101010010",
14086 => "0000000101010011",
14087 => "0000000101010011",
14088 => "0000000101010011",
14089 => "0000000101010011",
14090 => "0000000101010011",
14091 => "0000000101010011",
14092 => "0000000101010011",
14093 => "0000000101010011",
14094 => "0000000101010011",
14095 => "0000000101010011",
14096 => "0000000101010011",
14097 => "0000000101010011",
14098 => "0000000101010100",
14099 => "0000000101010100",
14100 => "0000000101010100",
14101 => "0000000101010100",
14102 => "0000000101010100",
14103 => "0000000101010100",
14104 => "0000000101010100",
14105 => "0000000101010100",
14106 => "0000000101010100",
14107 => "0000000101010100",
14108 => "0000000101010100",
14109 => "0000000101010100",
14110 => "0000000101010101",
14111 => "0000000101010101",
14112 => "0000000101010101",
14113 => "0000000101010101",
14114 => "0000000101010101",
14115 => "0000000101010101",
14116 => "0000000101010101",
14117 => "0000000101010101",
14118 => "0000000101010101",
14119 => "0000000101010101",
14120 => "0000000101010101",
14121 => "0000000101010101",
14122 => "0000000101010110",
14123 => "0000000101010110",
14124 => "0000000101010110",
14125 => "0000000101010110",
14126 => "0000000101010110",
14127 => "0000000101010110",
14128 => "0000000101010110",
14129 => "0000000101010110",
14130 => "0000000101010110",
14131 => "0000000101010110",
14132 => "0000000101010110",
14133 => "0000000101010110",
14134 => "0000000101010111",
14135 => "0000000101010111",
14136 => "0000000101010111",
14137 => "0000000101010111",
14138 => "0000000101010111",
14139 => "0000000101010111",
14140 => "0000000101010111",
14141 => "0000000101010111",
14142 => "0000000101010111",
14143 => "0000000101010111",
14144 => "0000000101010111",
14145 => "0000000101010111",
14146 => "0000000101011000",
14147 => "0000000101011000",
14148 => "0000000101011000",
14149 => "0000000101011000",
14150 => "0000000101011000",
14151 => "0000000101011000",
14152 => "0000000101011000",
14153 => "0000000101011000",
14154 => "0000000101011000",
14155 => "0000000101011000",
14156 => "0000000101011000",
14157 => "0000000101011000",
14158 => "0000000101011001",
14159 => "0000000101011001",
14160 => "0000000101011001",
14161 => "0000000101011001",
14162 => "0000000101011001",
14163 => "0000000101011001",
14164 => "0000000101011001",
14165 => "0000000101011001",
14166 => "0000000101011001",
14167 => "0000000101011001",
14168 => "0000000101011001",
14169 => "0000000101011001",
14170 => "0000000101011010",
14171 => "0000000101011010",
14172 => "0000000101011010",
14173 => "0000000101011010",
14174 => "0000000101011010",
14175 => "0000000101011010",
14176 => "0000000101011010",
14177 => "0000000101011010",
14178 => "0000000101011010",
14179 => "0000000101011010",
14180 => "0000000101011010",
14181 => "0000000101011010",
14182 => "0000000101011011",
14183 => "0000000101011011",
14184 => "0000000101011011",
14185 => "0000000101011011",
14186 => "0000000101011011",
14187 => "0000000101011011",
14188 => "0000000101011011",
14189 => "0000000101011011",
14190 => "0000000101011011",
14191 => "0000000101011011",
14192 => "0000000101011011",
14193 => "0000000101011011",
14194 => "0000000101011100",
14195 => "0000000101011100",
14196 => "0000000101011100",
14197 => "0000000101011100",
14198 => "0000000101011100",
14199 => "0000000101011100",
14200 => "0000000101011100",
14201 => "0000000101011100",
14202 => "0000000101011100",
14203 => "0000000101011100",
14204 => "0000000101011100",
14205 => "0000000101011100",
14206 => "0000000101011101",
14207 => "0000000101011101",
14208 => "0000000101011101",
14209 => "0000000101011101",
14210 => "0000000101011101",
14211 => "0000000101011101",
14212 => "0000000101011101",
14213 => "0000000101011101",
14214 => "0000000101011101",
14215 => "0000000101011101",
14216 => "0000000101011101",
14217 => "0000000101011101",
14218 => "0000000101011110",
14219 => "0000000101011110",
14220 => "0000000101011110",
14221 => "0000000101011110",
14222 => "0000000101011110",
14223 => "0000000101011110",
14224 => "0000000101011110",
14225 => "0000000101011110",
14226 => "0000000101011110",
14227 => "0000000101011110",
14228 => "0000000101011110",
14229 => "0000000101011110",
14230 => "0000000101011111",
14231 => "0000000101011111",
14232 => "0000000101011111",
14233 => "0000000101011111",
14234 => "0000000101011111",
14235 => "0000000101011111",
14236 => "0000000101011111",
14237 => "0000000101011111",
14238 => "0000000101011111",
14239 => "0000000101011111",
14240 => "0000000101011111",
14241 => "0000000101011111",
14242 => "0000000101100000",
14243 => "0000000101100000",
14244 => "0000000101100000",
14245 => "0000000101100000",
14246 => "0000000101100000",
14247 => "0000000101100000",
14248 => "0000000101100000",
14249 => "0000000101100000",
14250 => "0000000101100000",
14251 => "0000000101100000",
14252 => "0000000101100000",
14253 => "0000000101100001",
14254 => "0000000101100001",
14255 => "0000000101100001",
14256 => "0000000101100001",
14257 => "0000000101100001",
14258 => "0000000101100001",
14259 => "0000000101100001",
14260 => "0000000101100001",
14261 => "0000000101100001",
14262 => "0000000101100001",
14263 => "0000000101100001",
14264 => "0000000101100001",
14265 => "0000000101100010",
14266 => "0000000101100010",
14267 => "0000000101100010",
14268 => "0000000101100010",
14269 => "0000000101100010",
14270 => "0000000101100010",
14271 => "0000000101100010",
14272 => "0000000101100010",
14273 => "0000000101100010",
14274 => "0000000101100010",
14275 => "0000000101100010",
14276 => "0000000101100010",
14277 => "0000000101100011",
14278 => "0000000101100011",
14279 => "0000000101100011",
14280 => "0000000101100011",
14281 => "0000000101100011",
14282 => "0000000101100011",
14283 => "0000000101100011",
14284 => "0000000101100011",
14285 => "0000000101100011",
14286 => "0000000101100011",
14287 => "0000000101100011",
14288 => "0000000101100100",
14289 => "0000000101100100",
14290 => "0000000101100100",
14291 => "0000000101100100",
14292 => "0000000101100100",
14293 => "0000000101100100",
14294 => "0000000101100100",
14295 => "0000000101100100",
14296 => "0000000101100100",
14297 => "0000000101100100",
14298 => "0000000101100100",
14299 => "0000000101100100",
14300 => "0000000101100101",
14301 => "0000000101100101",
14302 => "0000000101100101",
14303 => "0000000101100101",
14304 => "0000000101100101",
14305 => "0000000101100101",
14306 => "0000000101100101",
14307 => "0000000101100101",
14308 => "0000000101100101",
14309 => "0000000101100101",
14310 => "0000000101100101",
14311 => "0000000101100101",
14312 => "0000000101100110",
14313 => "0000000101100110",
14314 => "0000000101100110",
14315 => "0000000101100110",
14316 => "0000000101100110",
14317 => "0000000101100110",
14318 => "0000000101100110",
14319 => "0000000101100110",
14320 => "0000000101100110",
14321 => "0000000101100110",
14322 => "0000000101100110",
14323 => "0000000101100111",
14324 => "0000000101100111",
14325 => "0000000101100111",
14326 => "0000000101100111",
14327 => "0000000101100111",
14328 => "0000000101100111",
14329 => "0000000101100111",
14330 => "0000000101100111",
14331 => "0000000101100111",
14332 => "0000000101100111",
14333 => "0000000101100111",
14334 => "0000000101100111",
14335 => "0000000101101000",
14336 => "0000000101101000",
14337 => "0000000101101000",
14338 => "0000000101101000",
14339 => "0000000101101000",
14340 => "0000000101101000",
14341 => "0000000101101000",
14342 => "0000000101101000",
14343 => "0000000101101000",
14344 => "0000000101101000",
14345 => "0000000101101000",
14346 => "0000000101101001",
14347 => "0000000101101001",
14348 => "0000000101101001",
14349 => "0000000101101001",
14350 => "0000000101101001",
14351 => "0000000101101001",
14352 => "0000000101101001",
14353 => "0000000101101001",
14354 => "0000000101101001",
14355 => "0000000101101001",
14356 => "0000000101101001",
14357 => "0000000101101001",
14358 => "0000000101101010",
14359 => "0000000101101010",
14360 => "0000000101101010",
14361 => "0000000101101010",
14362 => "0000000101101010",
14363 => "0000000101101010",
14364 => "0000000101101010",
14365 => "0000000101101010",
14366 => "0000000101101010",
14367 => "0000000101101010",
14368 => "0000000101101010",
14369 => "0000000101101011",
14370 => "0000000101101011",
14371 => "0000000101101011",
14372 => "0000000101101011",
14373 => "0000000101101011",
14374 => "0000000101101011",
14375 => "0000000101101011",
14376 => "0000000101101011",
14377 => "0000000101101011",
14378 => "0000000101101011",
14379 => "0000000101101011",
14380 => "0000000101101100",
14381 => "0000000101101100",
14382 => "0000000101101100",
14383 => "0000000101101100",
14384 => "0000000101101100",
14385 => "0000000101101100",
14386 => "0000000101101100",
14387 => "0000000101101100",
14388 => "0000000101101100",
14389 => "0000000101101100",
14390 => "0000000101101100",
14391 => "0000000101101100",
14392 => "0000000101101101",
14393 => "0000000101101101",
14394 => "0000000101101101",
14395 => "0000000101101101",
14396 => "0000000101101101",
14397 => "0000000101101101",
14398 => "0000000101101101",
14399 => "0000000101101101",
14400 => "0000000101101101",
14401 => "0000000101101101",
14402 => "0000000101101101",
14403 => "0000000101101110",
14404 => "0000000101101110",
14405 => "0000000101101110",
14406 => "0000000101101110",
14407 => "0000000101101110",
14408 => "0000000101101110",
14409 => "0000000101101110",
14410 => "0000000101101110",
14411 => "0000000101101110",
14412 => "0000000101101110",
14413 => "0000000101101110",
14414 => "0000000101101111",
14415 => "0000000101101111",
14416 => "0000000101101111",
14417 => "0000000101101111",
14418 => "0000000101101111",
14419 => "0000000101101111",
14420 => "0000000101101111",
14421 => "0000000101101111",
14422 => "0000000101101111",
14423 => "0000000101101111",
14424 => "0000000101101111",
14425 => "0000000101101111",
14426 => "0000000101110000",
14427 => "0000000101110000",
14428 => "0000000101110000",
14429 => "0000000101110000",
14430 => "0000000101110000",
14431 => "0000000101110000",
14432 => "0000000101110000",
14433 => "0000000101110000",
14434 => "0000000101110000",
14435 => "0000000101110000",
14436 => "0000000101110000",
14437 => "0000000101110001",
14438 => "0000000101110001",
14439 => "0000000101110001",
14440 => "0000000101110001",
14441 => "0000000101110001",
14442 => "0000000101110001",
14443 => "0000000101110001",
14444 => "0000000101110001",
14445 => "0000000101110001",
14446 => "0000000101110001",
14447 => "0000000101110001",
14448 => "0000000101110010",
14449 => "0000000101110010",
14450 => "0000000101110010",
14451 => "0000000101110010",
14452 => "0000000101110010",
14453 => "0000000101110010",
14454 => "0000000101110010",
14455 => "0000000101110010",
14456 => "0000000101110010",
14457 => "0000000101110010",
14458 => "0000000101110010",
14459 => "0000000101110011",
14460 => "0000000101110011",
14461 => "0000000101110011",
14462 => "0000000101110011",
14463 => "0000000101110011",
14464 => "0000000101110011",
14465 => "0000000101110011",
14466 => "0000000101110011",
14467 => "0000000101110011",
14468 => "0000000101110011",
14469 => "0000000101110011",
14470 => "0000000101110100",
14471 => "0000000101110100",
14472 => "0000000101110100",
14473 => "0000000101110100",
14474 => "0000000101110100",
14475 => "0000000101110100",
14476 => "0000000101110100",
14477 => "0000000101110100",
14478 => "0000000101110100",
14479 => "0000000101110100",
14480 => "0000000101110100",
14481 => "0000000101110100",
14482 => "0000000101110101",
14483 => "0000000101110101",
14484 => "0000000101110101",
14485 => "0000000101110101",
14486 => "0000000101110101",
14487 => "0000000101110101",
14488 => "0000000101110101",
14489 => "0000000101110101",
14490 => "0000000101110101",
14491 => "0000000101110101",
14492 => "0000000101110101",
14493 => "0000000101110110",
14494 => "0000000101110110",
14495 => "0000000101110110",
14496 => "0000000101110110",
14497 => "0000000101110110",
14498 => "0000000101110110",
14499 => "0000000101110110",
14500 => "0000000101110110",
14501 => "0000000101110110",
14502 => "0000000101110110",
14503 => "0000000101110110",
14504 => "0000000101110111",
14505 => "0000000101110111",
14506 => "0000000101110111",
14507 => "0000000101110111",
14508 => "0000000101110111",
14509 => "0000000101110111",
14510 => "0000000101110111",
14511 => "0000000101110111",
14512 => "0000000101110111",
14513 => "0000000101110111",
14514 => "0000000101110111",
14515 => "0000000101111000",
14516 => "0000000101111000",
14517 => "0000000101111000",
14518 => "0000000101111000",
14519 => "0000000101111000",
14520 => "0000000101111000",
14521 => "0000000101111000",
14522 => "0000000101111000",
14523 => "0000000101111000",
14524 => "0000000101111000",
14525 => "0000000101111000",
14526 => "0000000101111001",
14527 => "0000000101111001",
14528 => "0000000101111001",
14529 => "0000000101111001",
14530 => "0000000101111001",
14531 => "0000000101111001",
14532 => "0000000101111001",
14533 => "0000000101111001",
14534 => "0000000101111001",
14535 => "0000000101111001",
14536 => "0000000101111001",
14537 => "0000000101111010",
14538 => "0000000101111010",
14539 => "0000000101111010",
14540 => "0000000101111010",
14541 => "0000000101111010",
14542 => "0000000101111010",
14543 => "0000000101111010",
14544 => "0000000101111010",
14545 => "0000000101111010",
14546 => "0000000101111010",
14547 => "0000000101111010",
14548 => "0000000101111011",
14549 => "0000000101111011",
14550 => "0000000101111011",
14551 => "0000000101111011",
14552 => "0000000101111011",
14553 => "0000000101111011",
14554 => "0000000101111011",
14555 => "0000000101111011",
14556 => "0000000101111011",
14557 => "0000000101111011",
14558 => "0000000101111011",
14559 => "0000000101111100",
14560 => "0000000101111100",
14561 => "0000000101111100",
14562 => "0000000101111100",
14563 => "0000000101111100",
14564 => "0000000101111100",
14565 => "0000000101111100",
14566 => "0000000101111100",
14567 => "0000000101111100",
14568 => "0000000101111100",
14569 => "0000000101111100",
14570 => "0000000101111101",
14571 => "0000000101111101",
14572 => "0000000101111101",
14573 => "0000000101111101",
14574 => "0000000101111101",
14575 => "0000000101111101",
14576 => "0000000101111101",
14577 => "0000000101111101",
14578 => "0000000101111101",
14579 => "0000000101111101",
14580 => "0000000101111110",
14581 => "0000000101111110",
14582 => "0000000101111110",
14583 => "0000000101111110",
14584 => "0000000101111110",
14585 => "0000000101111110",
14586 => "0000000101111110",
14587 => "0000000101111110",
14588 => "0000000101111110",
14589 => "0000000101111110",
14590 => "0000000101111110",
14591 => "0000000101111111",
14592 => "0000000101111111",
14593 => "0000000101111111",
14594 => "0000000101111111",
14595 => "0000000101111111",
14596 => "0000000101111111",
14597 => "0000000101111111",
14598 => "0000000101111111",
14599 => "0000000101111111",
14600 => "0000000101111111",
14601 => "0000000101111111",
14602 => "0000000110000000",
14603 => "0000000110000000",
14604 => "0000000110000000",
14605 => "0000000110000000",
14606 => "0000000110000000",
14607 => "0000000110000000",
14608 => "0000000110000000",
14609 => "0000000110000000",
14610 => "0000000110000000",
14611 => "0000000110000000",
14612 => "0000000110000000",
14613 => "0000000110000001",
14614 => "0000000110000001",
14615 => "0000000110000001",
14616 => "0000000110000001",
14617 => "0000000110000001",
14618 => "0000000110000001",
14619 => "0000000110000001",
14620 => "0000000110000001",
14621 => "0000000110000001",
14622 => "0000000110000001",
14623 => "0000000110000001",
14624 => "0000000110000010",
14625 => "0000000110000010",
14626 => "0000000110000010",
14627 => "0000000110000010",
14628 => "0000000110000010",
14629 => "0000000110000010",
14630 => "0000000110000010",
14631 => "0000000110000010",
14632 => "0000000110000010",
14633 => "0000000110000010",
14634 => "0000000110000011",
14635 => "0000000110000011",
14636 => "0000000110000011",
14637 => "0000000110000011",
14638 => "0000000110000011",
14639 => "0000000110000011",
14640 => "0000000110000011",
14641 => "0000000110000011",
14642 => "0000000110000011",
14643 => "0000000110000011",
14644 => "0000000110000011",
14645 => "0000000110000100",
14646 => "0000000110000100",
14647 => "0000000110000100",
14648 => "0000000110000100",
14649 => "0000000110000100",
14650 => "0000000110000100",
14651 => "0000000110000100",
14652 => "0000000110000100",
14653 => "0000000110000100",
14654 => "0000000110000100",
14655 => "0000000110000100",
14656 => "0000000110000101",
14657 => "0000000110000101",
14658 => "0000000110000101",
14659 => "0000000110000101",
14660 => "0000000110000101",
14661 => "0000000110000101",
14662 => "0000000110000101",
14663 => "0000000110000101",
14664 => "0000000110000101",
14665 => "0000000110000101",
14666 => "0000000110000110",
14667 => "0000000110000110",
14668 => "0000000110000110",
14669 => "0000000110000110",
14670 => "0000000110000110",
14671 => "0000000110000110",
14672 => "0000000110000110",
14673 => "0000000110000110",
14674 => "0000000110000110",
14675 => "0000000110000110",
14676 => "0000000110000110",
14677 => "0000000110000111",
14678 => "0000000110000111",
14679 => "0000000110000111",
14680 => "0000000110000111",
14681 => "0000000110000111",
14682 => "0000000110000111",
14683 => "0000000110000111",
14684 => "0000000110000111",
14685 => "0000000110000111",
14686 => "0000000110000111",
14687 => "0000000110000111",
14688 => "0000000110001000",
14689 => "0000000110001000",
14690 => "0000000110001000",
14691 => "0000000110001000",
14692 => "0000000110001000",
14693 => "0000000110001000",
14694 => "0000000110001000",
14695 => "0000000110001000",
14696 => "0000000110001000",
14697 => "0000000110001000",
14698 => "0000000110001001",
14699 => "0000000110001001",
14700 => "0000000110001001",
14701 => "0000000110001001",
14702 => "0000000110001001",
14703 => "0000000110001001",
14704 => "0000000110001001",
14705 => "0000000110001001",
14706 => "0000000110001001",
14707 => "0000000110001001",
14708 => "0000000110001001",
14709 => "0000000110001010",
14710 => "0000000110001010",
14711 => "0000000110001010",
14712 => "0000000110001010",
14713 => "0000000110001010",
14714 => "0000000110001010",
14715 => "0000000110001010",
14716 => "0000000110001010",
14717 => "0000000110001010",
14718 => "0000000110001010",
14719 => "0000000110001011",
14720 => "0000000110001011",
14721 => "0000000110001011",
14722 => "0000000110001011",
14723 => "0000000110001011",
14724 => "0000000110001011",
14725 => "0000000110001011",
14726 => "0000000110001011",
14727 => "0000000110001011",
14728 => "0000000110001011",
14729 => "0000000110001011",
14730 => "0000000110001100",
14731 => "0000000110001100",
14732 => "0000000110001100",
14733 => "0000000110001100",
14734 => "0000000110001100",
14735 => "0000000110001100",
14736 => "0000000110001100",
14737 => "0000000110001100",
14738 => "0000000110001100",
14739 => "0000000110001100",
14740 => "0000000110001101",
14741 => "0000000110001101",
14742 => "0000000110001101",
14743 => "0000000110001101",
14744 => "0000000110001101",
14745 => "0000000110001101",
14746 => "0000000110001101",
14747 => "0000000110001101",
14748 => "0000000110001101",
14749 => "0000000110001101",
14750 => "0000000110001101",
14751 => "0000000110001110",
14752 => "0000000110001110",
14753 => "0000000110001110",
14754 => "0000000110001110",
14755 => "0000000110001110",
14756 => "0000000110001110",
14757 => "0000000110001110",
14758 => "0000000110001110",
14759 => "0000000110001110",
14760 => "0000000110001110",
14761 => "0000000110001111",
14762 => "0000000110001111",
14763 => "0000000110001111",
14764 => "0000000110001111",
14765 => "0000000110001111",
14766 => "0000000110001111",
14767 => "0000000110001111",
14768 => "0000000110001111",
14769 => "0000000110001111",
14770 => "0000000110001111",
14771 => "0000000110010000",
14772 => "0000000110010000",
14773 => "0000000110010000",
14774 => "0000000110010000",
14775 => "0000000110010000",
14776 => "0000000110010000",
14777 => "0000000110010000",
14778 => "0000000110010000",
14779 => "0000000110010000",
14780 => "0000000110010000",
14781 => "0000000110010000",
14782 => "0000000110010001",
14783 => "0000000110010001",
14784 => "0000000110010001",
14785 => "0000000110010001",
14786 => "0000000110010001",
14787 => "0000000110010001",
14788 => "0000000110010001",
14789 => "0000000110010001",
14790 => "0000000110010001",
14791 => "0000000110010001",
14792 => "0000000110010010",
14793 => "0000000110010010",
14794 => "0000000110010010",
14795 => "0000000110010010",
14796 => "0000000110010010",
14797 => "0000000110010010",
14798 => "0000000110010010",
14799 => "0000000110010010",
14800 => "0000000110010010",
14801 => "0000000110010010",
14802 => "0000000110010011",
14803 => "0000000110010011",
14804 => "0000000110010011",
14805 => "0000000110010011",
14806 => "0000000110010011",
14807 => "0000000110010011",
14808 => "0000000110010011",
14809 => "0000000110010011",
14810 => "0000000110010011",
14811 => "0000000110010011",
14812 => "0000000110010011",
14813 => "0000000110010100",
14814 => "0000000110010100",
14815 => "0000000110010100",
14816 => "0000000110010100",
14817 => "0000000110010100",
14818 => "0000000110010100",
14819 => "0000000110010100",
14820 => "0000000110010100",
14821 => "0000000110010100",
14822 => "0000000110010100",
14823 => "0000000110010101",
14824 => "0000000110010101",
14825 => "0000000110010101",
14826 => "0000000110010101",
14827 => "0000000110010101",
14828 => "0000000110010101",
14829 => "0000000110010101",
14830 => "0000000110010101",
14831 => "0000000110010101",
14832 => "0000000110010101",
14833 => "0000000110010110",
14834 => "0000000110010110",
14835 => "0000000110010110",
14836 => "0000000110010110",
14837 => "0000000110010110",
14838 => "0000000110010110",
14839 => "0000000110010110",
14840 => "0000000110010110",
14841 => "0000000110010110",
14842 => "0000000110010110",
14843 => "0000000110010111",
14844 => "0000000110010111",
14845 => "0000000110010111",
14846 => "0000000110010111",
14847 => "0000000110010111",
14848 => "0000000110010111",
14849 => "0000000110010111",
14850 => "0000000110010111",
14851 => "0000000110010111",
14852 => "0000000110010111",
14853 => "0000000110010111",
14854 => "0000000110011000",
14855 => "0000000110011000",
14856 => "0000000110011000",
14857 => "0000000110011000",
14858 => "0000000110011000",
14859 => "0000000110011000",
14860 => "0000000110011000",
14861 => "0000000110011000",
14862 => "0000000110011000",
14863 => "0000000110011000",
14864 => "0000000110011001",
14865 => "0000000110011001",
14866 => "0000000110011001",
14867 => "0000000110011001",
14868 => "0000000110011001",
14869 => "0000000110011001",
14870 => "0000000110011001",
14871 => "0000000110011001",
14872 => "0000000110011001",
14873 => "0000000110011001",
14874 => "0000000110011010",
14875 => "0000000110011010",
14876 => "0000000110011010",
14877 => "0000000110011010",
14878 => "0000000110011010",
14879 => "0000000110011010",
14880 => "0000000110011010",
14881 => "0000000110011010",
14882 => "0000000110011010",
14883 => "0000000110011010",
14884 => "0000000110011011",
14885 => "0000000110011011",
14886 => "0000000110011011",
14887 => "0000000110011011",
14888 => "0000000110011011",
14889 => "0000000110011011",
14890 => "0000000110011011",
14891 => "0000000110011011",
14892 => "0000000110011011",
14893 => "0000000110011011",
14894 => "0000000110011100",
14895 => "0000000110011100",
14896 => "0000000110011100",
14897 => "0000000110011100",
14898 => "0000000110011100",
14899 => "0000000110011100",
14900 => "0000000110011100",
14901 => "0000000110011100",
14902 => "0000000110011100",
14903 => "0000000110011100",
14904 => "0000000110011101",
14905 => "0000000110011101",
14906 => "0000000110011101",
14907 => "0000000110011101",
14908 => "0000000110011101",
14909 => "0000000110011101",
14910 => "0000000110011101",
14911 => "0000000110011101",
14912 => "0000000110011101",
14913 => "0000000110011101",
14914 => "0000000110011110",
14915 => "0000000110011110",
14916 => "0000000110011110",
14917 => "0000000110011110",
14918 => "0000000110011110",
14919 => "0000000110011110",
14920 => "0000000110011110",
14921 => "0000000110011110",
14922 => "0000000110011110",
14923 => "0000000110011110",
14924 => "0000000110011111",
14925 => "0000000110011111",
14926 => "0000000110011111",
14927 => "0000000110011111",
14928 => "0000000110011111",
14929 => "0000000110011111",
14930 => "0000000110011111",
14931 => "0000000110011111",
14932 => "0000000110011111",
14933 => "0000000110011111",
14934 => "0000000110100000",
14935 => "0000000110100000",
14936 => "0000000110100000",
14937 => "0000000110100000",
14938 => "0000000110100000",
14939 => "0000000110100000",
14940 => "0000000110100000",
14941 => "0000000110100000",
14942 => "0000000110100000",
14943 => "0000000110100000",
14944 => "0000000110100001",
14945 => "0000000110100001",
14946 => "0000000110100001",
14947 => "0000000110100001",
14948 => "0000000110100001",
14949 => "0000000110100001",
14950 => "0000000110100001",
14951 => "0000000110100001",
14952 => "0000000110100001",
14953 => "0000000110100001",
14954 => "0000000110100010",
14955 => "0000000110100010",
14956 => "0000000110100010",
14957 => "0000000110100010",
14958 => "0000000110100010",
14959 => "0000000110100010",
14960 => "0000000110100010",
14961 => "0000000110100010",
14962 => "0000000110100010",
14963 => "0000000110100010",
14964 => "0000000110100011",
14965 => "0000000110100011",
14966 => "0000000110100011",
14967 => "0000000110100011",
14968 => "0000000110100011",
14969 => "0000000110100011",
14970 => "0000000110100011",
14971 => "0000000110100011",
14972 => "0000000110100011",
14973 => "0000000110100011",
14974 => "0000000110100100",
14975 => "0000000110100100",
14976 => "0000000110100100",
14977 => "0000000110100100",
14978 => "0000000110100100",
14979 => "0000000110100100",
14980 => "0000000110100100",
14981 => "0000000110100100",
14982 => "0000000110100100",
14983 => "0000000110100100",
14984 => "0000000110100101",
14985 => "0000000110100101",
14986 => "0000000110100101",
14987 => "0000000110100101",
14988 => "0000000110100101",
14989 => "0000000110100101",
14990 => "0000000110100101",
14991 => "0000000110100101",
14992 => "0000000110100101",
14993 => "0000000110100101",
14994 => "0000000110100110",
14995 => "0000000110100110",
14996 => "0000000110100110",
14997 => "0000000110100110",
14998 => "0000000110100110",
14999 => "0000000110100110",
15000 => "0000000110100110",
15001 => "0000000110100110",
15002 => "0000000110100110",
15003 => "0000000110100111",
15004 => "0000000110100111",
15005 => "0000000110100111",
15006 => "0000000110100111",
15007 => "0000000110100111",
15008 => "0000000110100111",
15009 => "0000000110100111",
15010 => "0000000110100111",
15011 => "0000000110100111",
15012 => "0000000110100111",
15013 => "0000000110101000",
15014 => "0000000110101000",
15015 => "0000000110101000",
15016 => "0000000110101000",
15017 => "0000000110101000",
15018 => "0000000110101000",
15019 => "0000000110101000",
15020 => "0000000110101000",
15021 => "0000000110101000",
15022 => "0000000110101000",
15023 => "0000000110101001",
15024 => "0000000110101001",
15025 => "0000000110101001",
15026 => "0000000110101001",
15027 => "0000000110101001",
15028 => "0000000110101001",
15029 => "0000000110101001",
15030 => "0000000110101001",
15031 => "0000000110101001",
15032 => "0000000110101001",
15033 => "0000000110101010",
15034 => "0000000110101010",
15035 => "0000000110101010",
15036 => "0000000110101010",
15037 => "0000000110101010",
15038 => "0000000110101010",
15039 => "0000000110101010",
15040 => "0000000110101010",
15041 => "0000000110101010",
15042 => "0000000110101011",
15043 => "0000000110101011",
15044 => "0000000110101011",
15045 => "0000000110101011",
15046 => "0000000110101011",
15047 => "0000000110101011",
15048 => "0000000110101011",
15049 => "0000000110101011",
15050 => "0000000110101011",
15051 => "0000000110101011",
15052 => "0000000110101100",
15053 => "0000000110101100",
15054 => "0000000110101100",
15055 => "0000000110101100",
15056 => "0000000110101100",
15057 => "0000000110101100",
15058 => "0000000110101100",
15059 => "0000000110101100",
15060 => "0000000110101100",
15061 => "0000000110101100",
15062 => "0000000110101101",
15063 => "0000000110101101",
15064 => "0000000110101101",
15065 => "0000000110101101",
15066 => "0000000110101101",
15067 => "0000000110101101",
15068 => "0000000110101101",
15069 => "0000000110101101",
15070 => "0000000110101101",
15071 => "0000000110101110",
15072 => "0000000110101110",
15073 => "0000000110101110",
15074 => "0000000110101110",
15075 => "0000000110101110",
15076 => "0000000110101110",
15077 => "0000000110101110",
15078 => "0000000110101110",
15079 => "0000000110101110",
15080 => "0000000110101110",
15081 => "0000000110101111",
15082 => "0000000110101111",
15083 => "0000000110101111",
15084 => "0000000110101111",
15085 => "0000000110101111",
15086 => "0000000110101111",
15087 => "0000000110101111",
15088 => "0000000110101111",
15089 => "0000000110101111",
15090 => "0000000110101111",
15091 => "0000000110110000",
15092 => "0000000110110000",
15093 => "0000000110110000",
15094 => "0000000110110000",
15095 => "0000000110110000",
15096 => "0000000110110000",
15097 => "0000000110110000",
15098 => "0000000110110000",
15099 => "0000000110110000",
15100 => "0000000110110001",
15101 => "0000000110110001",
15102 => "0000000110110001",
15103 => "0000000110110001",
15104 => "0000000110110001",
15105 => "0000000110110001",
15106 => "0000000110110001",
15107 => "0000000110110001",
15108 => "0000000110110001",
15109 => "0000000110110001",
15110 => "0000000110110010",
15111 => "0000000110110010",
15112 => "0000000110110010",
15113 => "0000000110110010",
15114 => "0000000110110010",
15115 => "0000000110110010",
15116 => "0000000110110010",
15117 => "0000000110110010",
15118 => "0000000110110010",
15119 => "0000000110110011",
15120 => "0000000110110011",
15121 => "0000000110110011",
15122 => "0000000110110011",
15123 => "0000000110110011",
15124 => "0000000110110011",
15125 => "0000000110110011",
15126 => "0000000110110011",
15127 => "0000000110110011",
15128 => "0000000110110011",
15129 => "0000000110110100",
15130 => "0000000110110100",
15131 => "0000000110110100",
15132 => "0000000110110100",
15133 => "0000000110110100",
15134 => "0000000110110100",
15135 => "0000000110110100",
15136 => "0000000110110100",
15137 => "0000000110110100",
15138 => "0000000110110100",
15139 => "0000000110110101",
15140 => "0000000110110101",
15141 => "0000000110110101",
15142 => "0000000110110101",
15143 => "0000000110110101",
15144 => "0000000110110101",
15145 => "0000000110110101",
15146 => "0000000110110101",
15147 => "0000000110110101",
15148 => "0000000110110110",
15149 => "0000000110110110",
15150 => "0000000110110110",
15151 => "0000000110110110",
15152 => "0000000110110110",
15153 => "0000000110110110",
15154 => "0000000110110110",
15155 => "0000000110110110",
15156 => "0000000110110110",
15157 => "0000000110110111",
15158 => "0000000110110111",
15159 => "0000000110110111",
15160 => "0000000110110111",
15161 => "0000000110110111",
15162 => "0000000110110111",
15163 => "0000000110110111",
15164 => "0000000110110111",
15165 => "0000000110110111",
15166 => "0000000110110111",
15167 => "0000000110111000",
15168 => "0000000110111000",
15169 => "0000000110111000",
15170 => "0000000110111000",
15171 => "0000000110111000",
15172 => "0000000110111000",
15173 => "0000000110111000",
15174 => "0000000110111000",
15175 => "0000000110111000",
15176 => "0000000110111001",
15177 => "0000000110111001",
15178 => "0000000110111001",
15179 => "0000000110111001",
15180 => "0000000110111001",
15181 => "0000000110111001",
15182 => "0000000110111001",
15183 => "0000000110111001",
15184 => "0000000110111001",
15185 => "0000000110111001",
15186 => "0000000110111010",
15187 => "0000000110111010",
15188 => "0000000110111010",
15189 => "0000000110111010",
15190 => "0000000110111010",
15191 => "0000000110111010",
15192 => "0000000110111010",
15193 => "0000000110111010",
15194 => "0000000110111010",
15195 => "0000000110111011",
15196 => "0000000110111011",
15197 => "0000000110111011",
15198 => "0000000110111011",
15199 => "0000000110111011",
15200 => "0000000110111011",
15201 => "0000000110111011",
15202 => "0000000110111011",
15203 => "0000000110111011",
15204 => "0000000110111011",
15205 => "0000000110111100",
15206 => "0000000110111100",
15207 => "0000000110111100",
15208 => "0000000110111100",
15209 => "0000000110111100",
15210 => "0000000110111100",
15211 => "0000000110111100",
15212 => "0000000110111100",
15213 => "0000000110111100",
15214 => "0000000110111101",
15215 => "0000000110111101",
15216 => "0000000110111101",
15217 => "0000000110111101",
15218 => "0000000110111101",
15219 => "0000000110111101",
15220 => "0000000110111101",
15221 => "0000000110111101",
15222 => "0000000110111101",
15223 => "0000000110111110",
15224 => "0000000110111110",
15225 => "0000000110111110",
15226 => "0000000110111110",
15227 => "0000000110111110",
15228 => "0000000110111110",
15229 => "0000000110111110",
15230 => "0000000110111110",
15231 => "0000000110111110",
15232 => "0000000110111111",
15233 => "0000000110111111",
15234 => "0000000110111111",
15235 => "0000000110111111",
15236 => "0000000110111111",
15237 => "0000000110111111",
15238 => "0000000110111111",
15239 => "0000000110111111",
15240 => "0000000110111111",
15241 => "0000000110111111",
15242 => "0000000111000000",
15243 => "0000000111000000",
15244 => "0000000111000000",
15245 => "0000000111000000",
15246 => "0000000111000000",
15247 => "0000000111000000",
15248 => "0000000111000000",
15249 => "0000000111000000",
15250 => "0000000111000000",
15251 => "0000000111000001",
15252 => "0000000111000001",
15253 => "0000000111000001",
15254 => "0000000111000001",
15255 => "0000000111000001",
15256 => "0000000111000001",
15257 => "0000000111000001",
15258 => "0000000111000001",
15259 => "0000000111000001",
15260 => "0000000111000010",
15261 => "0000000111000010",
15262 => "0000000111000010",
15263 => "0000000111000010",
15264 => "0000000111000010",
15265 => "0000000111000010",
15266 => "0000000111000010",
15267 => "0000000111000010",
15268 => "0000000111000010",
15269 => "0000000111000011",
15270 => "0000000111000011",
15271 => "0000000111000011",
15272 => "0000000111000011",
15273 => "0000000111000011",
15274 => "0000000111000011",
15275 => "0000000111000011",
15276 => "0000000111000011",
15277 => "0000000111000011",
15278 => "0000000111000011",
15279 => "0000000111000100",
15280 => "0000000111000100",
15281 => "0000000111000100",
15282 => "0000000111000100",
15283 => "0000000111000100",
15284 => "0000000111000100",
15285 => "0000000111000100",
15286 => "0000000111000100",
15287 => "0000000111000100",
15288 => "0000000111000101",
15289 => "0000000111000101",
15290 => "0000000111000101",
15291 => "0000000111000101",
15292 => "0000000111000101",
15293 => "0000000111000101",
15294 => "0000000111000101",
15295 => "0000000111000101",
15296 => "0000000111000101",
15297 => "0000000111000110",
15298 => "0000000111000110",
15299 => "0000000111000110",
15300 => "0000000111000110",
15301 => "0000000111000110",
15302 => "0000000111000110",
15303 => "0000000111000110",
15304 => "0000000111000110",
15305 => "0000000111000110",
15306 => "0000000111000111",
15307 => "0000000111000111",
15308 => "0000000111000111",
15309 => "0000000111000111",
15310 => "0000000111000111",
15311 => "0000000111000111",
15312 => "0000000111000111",
15313 => "0000000111000111",
15314 => "0000000111000111",
15315 => "0000000111001000",
15316 => "0000000111001000",
15317 => "0000000111001000",
15318 => "0000000111001000",
15319 => "0000000111001000",
15320 => "0000000111001000",
15321 => "0000000111001000",
15322 => "0000000111001000",
15323 => "0000000111001000",
15324 => "0000000111001001",
15325 => "0000000111001001",
15326 => "0000000111001001",
15327 => "0000000111001001",
15328 => "0000000111001001",
15329 => "0000000111001001",
15330 => "0000000111001001",
15331 => "0000000111001001",
15332 => "0000000111001001",
15333 => "0000000111001010",
15334 => "0000000111001010",
15335 => "0000000111001010",
15336 => "0000000111001010",
15337 => "0000000111001010",
15338 => "0000000111001010",
15339 => "0000000111001010",
15340 => "0000000111001010",
15341 => "0000000111001010",
15342 => "0000000111001010",
15343 => "0000000111001011",
15344 => "0000000111001011",
15345 => "0000000111001011",
15346 => "0000000111001011",
15347 => "0000000111001011",
15348 => "0000000111001011",
15349 => "0000000111001011",
15350 => "0000000111001011",
15351 => "0000000111001011",
15352 => "0000000111001100",
15353 => "0000000111001100",
15354 => "0000000111001100",
15355 => "0000000111001100",
15356 => "0000000111001100",
15357 => "0000000111001100",
15358 => "0000000111001100",
15359 => "0000000111001100",
15360 => "0000000111001100",
15361 => "0000000111001101",
15362 => "0000000111001101",
15363 => "0000000111001101",
15364 => "0000000111001101",
15365 => "0000000111001101",
15366 => "0000000111001101",
15367 => "0000000111001101",
15368 => "0000000111001101",
15369 => "0000000111001101",
15370 => "0000000111001110",
15371 => "0000000111001110",
15372 => "0000000111001110",
15373 => "0000000111001110",
15374 => "0000000111001110",
15375 => "0000000111001110",
15376 => "0000000111001110",
15377 => "0000000111001110",
15378 => "0000000111001110",
15379 => "0000000111001111",
15380 => "0000000111001111",
15381 => "0000000111001111",
15382 => "0000000111001111",
15383 => "0000000111001111",
15384 => "0000000111001111",
15385 => "0000000111001111",
15386 => "0000000111001111",
15387 => "0000000111001111",
15388 => "0000000111010000",
15389 => "0000000111010000",
15390 => "0000000111010000",
15391 => "0000000111010000",
15392 => "0000000111010000",
15393 => "0000000111010000",
15394 => "0000000111010000",
15395 => "0000000111010000",
15396 => "0000000111010000",
15397 => "0000000111010001",
15398 => "0000000111010001",
15399 => "0000000111010001",
15400 => "0000000111010001",
15401 => "0000000111010001",
15402 => "0000000111010001",
15403 => "0000000111010001",
15404 => "0000000111010001",
15405 => "0000000111010010",
15406 => "0000000111010010",
15407 => "0000000111010010",
15408 => "0000000111010010",
15409 => "0000000111010010",
15410 => "0000000111010010",
15411 => "0000000111010010",
15412 => "0000000111010010",
15413 => "0000000111010010",
15414 => "0000000111010011",
15415 => "0000000111010011",
15416 => "0000000111010011",
15417 => "0000000111010011",
15418 => "0000000111010011",
15419 => "0000000111010011",
15420 => "0000000111010011",
15421 => "0000000111010011",
15422 => "0000000111010011",
15423 => "0000000111010100",
15424 => "0000000111010100",
15425 => "0000000111010100",
15426 => "0000000111010100",
15427 => "0000000111010100",
15428 => "0000000111010100",
15429 => "0000000111010100",
15430 => "0000000111010100",
15431 => "0000000111010100",
15432 => "0000000111010101",
15433 => "0000000111010101",
15434 => "0000000111010101",
15435 => "0000000111010101",
15436 => "0000000111010101",
15437 => "0000000111010101",
15438 => "0000000111010101",
15439 => "0000000111010101",
15440 => "0000000111010101",
15441 => "0000000111010110",
15442 => "0000000111010110",
15443 => "0000000111010110",
15444 => "0000000111010110",
15445 => "0000000111010110",
15446 => "0000000111010110",
15447 => "0000000111010110",
15448 => "0000000111010110",
15449 => "0000000111010110",
15450 => "0000000111010111",
15451 => "0000000111010111",
15452 => "0000000111010111",
15453 => "0000000111010111",
15454 => "0000000111010111",
15455 => "0000000111010111",
15456 => "0000000111010111",
15457 => "0000000111010111",
15458 => "0000000111010111",
15459 => "0000000111011000",
15460 => "0000000111011000",
15461 => "0000000111011000",
15462 => "0000000111011000",
15463 => "0000000111011000",
15464 => "0000000111011000",
15465 => "0000000111011000",
15466 => "0000000111011000",
15467 => "0000000111011001",
15468 => "0000000111011001",
15469 => "0000000111011001",
15470 => "0000000111011001",
15471 => "0000000111011001",
15472 => "0000000111011001",
15473 => "0000000111011001",
15474 => "0000000111011001",
15475 => "0000000111011001",
15476 => "0000000111011010",
15477 => "0000000111011010",
15478 => "0000000111011010",
15479 => "0000000111011010",
15480 => "0000000111011010",
15481 => "0000000111011010",
15482 => "0000000111011010",
15483 => "0000000111011010",
15484 => "0000000111011010",
15485 => "0000000111011011",
15486 => "0000000111011011",
15487 => "0000000111011011",
15488 => "0000000111011011",
15489 => "0000000111011011",
15490 => "0000000111011011",
15491 => "0000000111011011",
15492 => "0000000111011011",
15493 => "0000000111011011",
15494 => "0000000111011100",
15495 => "0000000111011100",
15496 => "0000000111011100",
15497 => "0000000111011100",
15498 => "0000000111011100",
15499 => "0000000111011100",
15500 => "0000000111011100",
15501 => "0000000111011100",
15502 => "0000000111011101",
15503 => "0000000111011101",
15504 => "0000000111011101",
15505 => "0000000111011101",
15506 => "0000000111011101",
15507 => "0000000111011101",
15508 => "0000000111011101",
15509 => "0000000111011101",
15510 => "0000000111011101",
15511 => "0000000111011110",
15512 => "0000000111011110",
15513 => "0000000111011110",
15514 => "0000000111011110",
15515 => "0000000111011110",
15516 => "0000000111011110",
15517 => "0000000111011110",
15518 => "0000000111011110",
15519 => "0000000111011110",
15520 => "0000000111011111",
15521 => "0000000111011111",
15522 => "0000000111011111",
15523 => "0000000111011111",
15524 => "0000000111011111",
15525 => "0000000111011111",
15526 => "0000000111011111",
15527 => "0000000111011111",
15528 => "0000000111100000",
15529 => "0000000111100000",
15530 => "0000000111100000",
15531 => "0000000111100000",
15532 => "0000000111100000",
15533 => "0000000111100000",
15534 => "0000000111100000",
15535 => "0000000111100000",
15536 => "0000000111100000",
15537 => "0000000111100001",
15538 => "0000000111100001",
15539 => "0000000111100001",
15540 => "0000000111100001",
15541 => "0000000111100001",
15542 => "0000000111100001",
15543 => "0000000111100001",
15544 => "0000000111100001",
15545 => "0000000111100001",
15546 => "0000000111100010",
15547 => "0000000111100010",
15548 => "0000000111100010",
15549 => "0000000111100010",
15550 => "0000000111100010",
15551 => "0000000111100010",
15552 => "0000000111100010",
15553 => "0000000111100010",
15554 => "0000000111100011",
15555 => "0000000111100011",
15556 => "0000000111100011",
15557 => "0000000111100011",
15558 => "0000000111100011",
15559 => "0000000111100011",
15560 => "0000000111100011",
15561 => "0000000111100011",
15562 => "0000000111100011",
15563 => "0000000111100100",
15564 => "0000000111100100",
15565 => "0000000111100100",
15566 => "0000000111100100",
15567 => "0000000111100100",
15568 => "0000000111100100",
15569 => "0000000111100100",
15570 => "0000000111100100",
15571 => "0000000111100100",
15572 => "0000000111100101",
15573 => "0000000111100101",
15574 => "0000000111100101",
15575 => "0000000111100101",
15576 => "0000000111100101",
15577 => "0000000111100101",
15578 => "0000000111100101",
15579 => "0000000111100101",
15580 => "0000000111100110",
15581 => "0000000111100110",
15582 => "0000000111100110",
15583 => "0000000111100110",
15584 => "0000000111100110",
15585 => "0000000111100110",
15586 => "0000000111100110",
15587 => "0000000111100110",
15588 => "0000000111100110",
15589 => "0000000111100111",
15590 => "0000000111100111",
15591 => "0000000111100111",
15592 => "0000000111100111",
15593 => "0000000111100111",
15594 => "0000000111100111",
15595 => "0000000111100111",
15596 => "0000000111100111",
15597 => "0000000111101000",
15598 => "0000000111101000",
15599 => "0000000111101000",
15600 => "0000000111101000",
15601 => "0000000111101000",
15602 => "0000000111101000",
15603 => "0000000111101000",
15604 => "0000000111101000",
15605 => "0000000111101000",
15606 => "0000000111101001",
15607 => "0000000111101001",
15608 => "0000000111101001",
15609 => "0000000111101001",
15610 => "0000000111101001",
15611 => "0000000111101001",
15612 => "0000000111101001",
15613 => "0000000111101001",
15614 => "0000000111101010",
15615 => "0000000111101010",
15616 => "0000000111101010",
15617 => "0000000111101010",
15618 => "0000000111101010",
15619 => "0000000111101010",
15620 => "0000000111101010",
15621 => "0000000111101010",
15622 => "0000000111101010",
15623 => "0000000111101011",
15624 => "0000000111101011",
15625 => "0000000111101011",
15626 => "0000000111101011",
15627 => "0000000111101011",
15628 => "0000000111101011",
15629 => "0000000111101011",
15630 => "0000000111101011",
15631 => "0000000111101100",
15632 => "0000000111101100",
15633 => "0000000111101100",
15634 => "0000000111101100",
15635 => "0000000111101100",
15636 => "0000000111101100",
15637 => "0000000111101100",
15638 => "0000000111101100",
15639 => "0000000111101100",
15640 => "0000000111101101",
15641 => "0000000111101101",
15642 => "0000000111101101",
15643 => "0000000111101101",
15644 => "0000000111101101",
15645 => "0000000111101101",
15646 => "0000000111101101",
15647 => "0000000111101101",
15648 => "0000000111101110",
15649 => "0000000111101110",
15650 => "0000000111101110",
15651 => "0000000111101110",
15652 => "0000000111101110",
15653 => "0000000111101110",
15654 => "0000000111101110",
15655 => "0000000111101110",
15656 => "0000000111101111",
15657 => "0000000111101111",
15658 => "0000000111101111",
15659 => "0000000111101111",
15660 => "0000000111101111",
15661 => "0000000111101111",
15662 => "0000000111101111",
15663 => "0000000111101111",
15664 => "0000000111101111",
15665 => "0000000111110000",
15666 => "0000000111110000",
15667 => "0000000111110000",
15668 => "0000000111110000",
15669 => "0000000111110000",
15670 => "0000000111110000",
15671 => "0000000111110000",
15672 => "0000000111110000",
15673 => "0000000111110001",
15674 => "0000000111110001",
15675 => "0000000111110001",
15676 => "0000000111110001",
15677 => "0000000111110001",
15678 => "0000000111110001",
15679 => "0000000111110001",
15680 => "0000000111110001",
15681 => "0000000111110001",
15682 => "0000000111110010",
15683 => "0000000111110010",
15684 => "0000000111110010",
15685 => "0000000111110010",
15686 => "0000000111110010",
15687 => "0000000111110010",
15688 => "0000000111110010",
15689 => "0000000111110010",
15690 => "0000000111110011",
15691 => "0000000111110011",
15692 => "0000000111110011",
15693 => "0000000111110011",
15694 => "0000000111110011",
15695 => "0000000111110011",
15696 => "0000000111110011",
15697 => "0000000111110011",
15698 => "0000000111110100",
15699 => "0000000111110100",
15700 => "0000000111110100",
15701 => "0000000111110100",
15702 => "0000000111110100",
15703 => "0000000111110100",
15704 => "0000000111110100",
15705 => "0000000111110100",
15706 => "0000000111110100",
15707 => "0000000111110101",
15708 => "0000000111110101",
15709 => "0000000111110101",
15710 => "0000000111110101",
15711 => "0000000111110101",
15712 => "0000000111110101",
15713 => "0000000111110101",
15714 => "0000000111110101",
15715 => "0000000111110110",
15716 => "0000000111110110",
15717 => "0000000111110110",
15718 => "0000000111110110",
15719 => "0000000111110110",
15720 => "0000000111110110",
15721 => "0000000111110110",
15722 => "0000000111110110",
15723 => "0000000111110111",
15724 => "0000000111110111",
15725 => "0000000111110111",
15726 => "0000000111110111",
15727 => "0000000111110111",
15728 => "0000000111110111",
15729 => "0000000111110111",
15730 => "0000000111110111",
15731 => "0000000111111000",
15732 => "0000000111111000",
15733 => "0000000111111000",
15734 => "0000000111111000",
15735 => "0000000111111000",
15736 => "0000000111111000",
15737 => "0000000111111000",
15738 => "0000000111111000",
15739 => "0000000111111000",
15740 => "0000000111111001",
15741 => "0000000111111001",
15742 => "0000000111111001",
15743 => "0000000111111001",
15744 => "0000000111111001",
15745 => "0000000111111001",
15746 => "0000000111111001",
15747 => "0000000111111001",
15748 => "0000000111111010",
15749 => "0000000111111010",
15750 => "0000000111111010",
15751 => "0000000111111010",
15752 => "0000000111111010",
15753 => "0000000111111010",
15754 => "0000000111111010",
15755 => "0000000111111010",
15756 => "0000000111111011",
15757 => "0000000111111011",
15758 => "0000000111111011",
15759 => "0000000111111011",
15760 => "0000000111111011",
15761 => "0000000111111011",
15762 => "0000000111111011",
15763 => "0000000111111011",
15764 => "0000000111111100",
15765 => "0000000111111100",
15766 => "0000000111111100",
15767 => "0000000111111100",
15768 => "0000000111111100",
15769 => "0000000111111100",
15770 => "0000000111111100",
15771 => "0000000111111100",
15772 => "0000000111111100",
15773 => "0000000111111101",
15774 => "0000000111111101",
15775 => "0000000111111101",
15776 => "0000000111111101",
15777 => "0000000111111101",
15778 => "0000000111111101",
15779 => "0000000111111101",
15780 => "0000000111111101",
15781 => "0000000111111110",
15782 => "0000000111111110",
15783 => "0000000111111110",
15784 => "0000000111111110",
15785 => "0000000111111110",
15786 => "0000000111111110",
15787 => "0000000111111110",
15788 => "0000000111111110",
15789 => "0000000111111111",
15790 => "0000000111111111",
15791 => "0000000111111111",
15792 => "0000000111111111",
15793 => "0000000111111111",
15794 => "0000000111111111",
15795 => "0000000111111111",
15796 => "0000000111111111",
15797 => "0000001000000000",
15798 => "0000001000000000",
15799 => "0000001000000000",
15800 => "0000001000000000",
15801 => "0000001000000000",
15802 => "0000001000000000",
15803 => "0000001000000000",
15804 => "0000001000000001",
15805 => "0000001000000001",
15806 => "0000001000000001",
15807 => "0000001000000001",
15808 => "0000001000000001",
15809 => "0000001000000001",
15810 => "0000001000000001",
15811 => "0000001000000001",
15812 => "0000001000000010",
15813 => "0000001000000010",
15814 => "0000001000000010",
15815 => "0000001000000010",
15816 => "0000001000000010",
15817 => "0000001000000010",
15818 => "0000001000000010",
15819 => "0000001000000010",
15820 => "0000001000000011",
15821 => "0000001000000011",
15822 => "0000001000000011",
15823 => "0000001000000011",
15824 => "0000001000000011",
15825 => "0000001000000011",
15826 => "0000001000000011",
15827 => "0000001000000011",
15828 => "0000001000000100",
15829 => "0000001000000100",
15830 => "0000001000000100",
15831 => "0000001000000100",
15832 => "0000001000000100",
15833 => "0000001000000100",
15834 => "0000001000000100",
15835 => "0000001000000100",
15836 => "0000001000000101",
15837 => "0000001000000101",
15838 => "0000001000000101",
15839 => "0000001000000101",
15840 => "0000001000000101",
15841 => "0000001000000101",
15842 => "0000001000000101",
15843 => "0000001000000101",
15844 => "0000001000000110",
15845 => "0000001000000110",
15846 => "0000001000000110",
15847 => "0000001000000110",
15848 => "0000001000000110",
15849 => "0000001000000110",
15850 => "0000001000000110",
15851 => "0000001000000110",
15852 => "0000001000000111",
15853 => "0000001000000111",
15854 => "0000001000000111",
15855 => "0000001000000111",
15856 => "0000001000000111",
15857 => "0000001000000111",
15858 => "0000001000000111",
15859 => "0000001000000111",
15860 => "0000001000001000",
15861 => "0000001000001000",
15862 => "0000001000001000",
15863 => "0000001000001000",
15864 => "0000001000001000",
15865 => "0000001000001000",
15866 => "0000001000001000",
15867 => "0000001000001000",
15868 => "0000001000001001",
15869 => "0000001000001001",
15870 => "0000001000001001",
15871 => "0000001000001001",
15872 => "0000001000001001",
15873 => "0000001000001001",
15874 => "0000001000001001",
15875 => "0000001000001001",
15876 => "0000001000001010",
15877 => "0000001000001010",
15878 => "0000001000001010",
15879 => "0000001000001010",
15880 => "0000001000001010",
15881 => "0000001000001010",
15882 => "0000001000001010",
15883 => "0000001000001010",
15884 => "0000001000001011",
15885 => "0000001000001011",
15886 => "0000001000001011",
15887 => "0000001000001011",
15888 => "0000001000001011",
15889 => "0000001000001011",
15890 => "0000001000001011",
15891 => "0000001000001011",
15892 => "0000001000001100",
15893 => "0000001000001100",
15894 => "0000001000001100",
15895 => "0000001000001100",
15896 => "0000001000001100",
15897 => "0000001000001100",
15898 => "0000001000001100",
15899 => "0000001000001100",
15900 => "0000001000001101",
15901 => "0000001000001101",
15902 => "0000001000001101",
15903 => "0000001000001101",
15904 => "0000001000001101",
15905 => "0000001000001101",
15906 => "0000001000001101",
15907 => "0000001000001101",
15908 => "0000001000001110",
15909 => "0000001000001110",
15910 => "0000001000001110",
15911 => "0000001000001110",
15912 => "0000001000001110",
15913 => "0000001000001110",
15914 => "0000001000001110",
15915 => "0000001000001110",
15916 => "0000001000001111",
15917 => "0000001000001111",
15918 => "0000001000001111",
15919 => "0000001000001111",
15920 => "0000001000001111",
15921 => "0000001000001111",
15922 => "0000001000001111",
15923 => "0000001000001111",
15924 => "0000001000010000",
15925 => "0000001000010000",
15926 => "0000001000010000",
15927 => "0000001000010000",
15928 => "0000001000010000",
15929 => "0000001000010000",
15930 => "0000001000010000",
15931 => "0000001000010000",
15932 => "0000001000010001",
15933 => "0000001000010001",
15934 => "0000001000010001",
15935 => "0000001000010001",
15936 => "0000001000010001",
15937 => "0000001000010001",
15938 => "0000001000010001",
15939 => "0000001000010001",
15940 => "0000001000010010",
15941 => "0000001000010010",
15942 => "0000001000010010",
15943 => "0000001000010010",
15944 => "0000001000010010",
15945 => "0000001000010010",
15946 => "0000001000010010",
15947 => "0000001000010010",
15948 => "0000001000010011",
15949 => "0000001000010011",
15950 => "0000001000010011",
15951 => "0000001000010011",
15952 => "0000001000010011",
15953 => "0000001000010011",
15954 => "0000001000010011",
15955 => "0000001000010011",
15956 => "0000001000010100",
15957 => "0000001000010100",
15958 => "0000001000010100",
15959 => "0000001000010100",
15960 => "0000001000010100",
15961 => "0000001000010100",
15962 => "0000001000010100",
15963 => "0000001000010101",
15964 => "0000001000010101",
15965 => "0000001000010101",
15966 => "0000001000010101",
15967 => "0000001000010101",
15968 => "0000001000010101",
15969 => "0000001000010101",
15970 => "0000001000010101",
15971 => "0000001000010110",
15972 => "0000001000010110",
15973 => "0000001000010110",
15974 => "0000001000010110",
15975 => "0000001000010110",
15976 => "0000001000010110",
15977 => "0000001000010110",
15978 => "0000001000010110",
15979 => "0000001000010111",
15980 => "0000001000010111",
15981 => "0000001000010111",
15982 => "0000001000010111",
15983 => "0000001000010111",
15984 => "0000001000010111",
15985 => "0000001000010111",
15986 => "0000001000010111",
15987 => "0000001000011000",
15988 => "0000001000011000",
15989 => "0000001000011000",
15990 => "0000001000011000",
15991 => "0000001000011000",
15992 => "0000001000011000",
15993 => "0000001000011000",
15994 => "0000001000011001",
15995 => "0000001000011001",
15996 => "0000001000011001",
15997 => "0000001000011001",
15998 => "0000001000011001",
15999 => "0000001000011001",
16000 => "0000001000011001",
16001 => "0000001000011001",
16002 => "0000001000011010",
16003 => "0000001000011010",
16004 => "0000001000011010",
16005 => "0000001000011010",
16006 => "0000001000011010",
16007 => "0000001000011010",
16008 => "0000001000011010",
16009 => "0000001000011010",
16010 => "0000001000011011",
16011 => "0000001000011011",
16012 => "0000001000011011",
16013 => "0000001000011011",
16014 => "0000001000011011",
16015 => "0000001000011011",
16016 => "0000001000011011",
16017 => "0000001000011011",
16018 => "0000001000011100",
16019 => "0000001000011100",
16020 => "0000001000011100",
16021 => "0000001000011100",
16022 => "0000001000011100",
16023 => "0000001000011100",
16024 => "0000001000011100",
16025 => "0000001000011101",
16026 => "0000001000011101",
16027 => "0000001000011101",
16028 => "0000001000011101",
16029 => "0000001000011101",
16030 => "0000001000011101",
16031 => "0000001000011101",
16032 => "0000001000011101",
16033 => "0000001000011110",
16034 => "0000001000011110",
16035 => "0000001000011110",
16036 => "0000001000011110",
16037 => "0000001000011110",
16038 => "0000001000011110",
16039 => "0000001000011110",
16040 => "0000001000011110",
16041 => "0000001000011111",
16042 => "0000001000011111",
16043 => "0000001000011111",
16044 => "0000001000011111",
16045 => "0000001000011111",
16046 => "0000001000011111",
16047 => "0000001000011111",
16048 => "0000001000100000",
16049 => "0000001000100000",
16050 => "0000001000100000",
16051 => "0000001000100000",
16052 => "0000001000100000",
16053 => "0000001000100000",
16054 => "0000001000100000",
16055 => "0000001000100000",
16056 => "0000001000100001",
16057 => "0000001000100001",
16058 => "0000001000100001",
16059 => "0000001000100001",
16060 => "0000001000100001",
16061 => "0000001000100001",
16062 => "0000001000100001",
16063 => "0000001000100001",
16064 => "0000001000100010",
16065 => "0000001000100010",
16066 => "0000001000100010",
16067 => "0000001000100010",
16068 => "0000001000100010",
16069 => "0000001000100010",
16070 => "0000001000100010",
16071 => "0000001000100011",
16072 => "0000001000100011",
16073 => "0000001000100011",
16074 => "0000001000100011",
16075 => "0000001000100011",
16076 => "0000001000100011",
16077 => "0000001000100011",
16078 => "0000001000100011",
16079 => "0000001000100100",
16080 => "0000001000100100",
16081 => "0000001000100100",
16082 => "0000001000100100",
16083 => "0000001000100100",
16084 => "0000001000100100",
16085 => "0000001000100100",
16086 => "0000001000100100",
16087 => "0000001000100101",
16088 => "0000001000100101",
16089 => "0000001000100101",
16090 => "0000001000100101",
16091 => "0000001000100101",
16092 => "0000001000100101",
16093 => "0000001000100101",
16094 => "0000001000100110",
16095 => "0000001000100110",
16096 => "0000001000100110",
16097 => "0000001000100110",
16098 => "0000001000100110",
16099 => "0000001000100110",
16100 => "0000001000100110",
16101 => "0000001000100110",
16102 => "0000001000100111",
16103 => "0000001000100111",
16104 => "0000001000100111",
16105 => "0000001000100111",
16106 => "0000001000100111",
16107 => "0000001000100111",
16108 => "0000001000100111",
16109 => "0000001000101000",
16110 => "0000001000101000",
16111 => "0000001000101000",
16112 => "0000001000101000",
16113 => "0000001000101000",
16114 => "0000001000101000",
16115 => "0000001000101000",
16116 => "0000001000101000",
16117 => "0000001000101001",
16118 => "0000001000101001",
16119 => "0000001000101001",
16120 => "0000001000101001",
16121 => "0000001000101001",
16122 => "0000001000101001",
16123 => "0000001000101001",
16124 => "0000001000101010",
16125 => "0000001000101010",
16126 => "0000001000101010",
16127 => "0000001000101010",
16128 => "0000001000101010",
16129 => "0000001000101010",
16130 => "0000001000101010",
16131 => "0000001000101010",
16132 => "0000001000101011",
16133 => "0000001000101011",
16134 => "0000001000101011",
16135 => "0000001000101011",
16136 => "0000001000101011",
16137 => "0000001000101011",
16138 => "0000001000101011",
16139 => "0000001000101100",
16140 => "0000001000101100",
16141 => "0000001000101100",
16142 => "0000001000101100",
16143 => "0000001000101100",
16144 => "0000001000101100",
16145 => "0000001000101100",
16146 => "0000001000101100",
16147 => "0000001000101101",
16148 => "0000001000101101",
16149 => "0000001000101101",
16150 => "0000001000101101",
16151 => "0000001000101101",
16152 => "0000001000101101",
16153 => "0000001000101101",
16154 => "0000001000101110",
16155 => "0000001000101110",
16156 => "0000001000101110",
16157 => "0000001000101110",
16158 => "0000001000101110",
16159 => "0000001000101110",
16160 => "0000001000101110",
16161 => "0000001000101110",
16162 => "0000001000101111",
16163 => "0000001000101111",
16164 => "0000001000101111",
16165 => "0000001000101111",
16166 => "0000001000101111",
16167 => "0000001000101111",
16168 => "0000001000101111",
16169 => "0000001000110000",
16170 => "0000001000110000",
16171 => "0000001000110000",
16172 => "0000001000110000",
16173 => "0000001000110000",
16174 => "0000001000110000",
16175 => "0000001000110000",
16176 => "0000001000110000",
16177 => "0000001000110001",
16178 => "0000001000110001",
16179 => "0000001000110001",
16180 => "0000001000110001",
16181 => "0000001000110001",
16182 => "0000001000110001",
16183 => "0000001000110001",
16184 => "0000001000110010",
16185 => "0000001000110010",
16186 => "0000001000110010",
16187 => "0000001000110010",
16188 => "0000001000110010",
16189 => "0000001000110010",
16190 => "0000001000110010",
16191 => "0000001000110010",
16192 => "0000001000110011",
16193 => "0000001000110011",
16194 => "0000001000110011",
16195 => "0000001000110011",
16196 => "0000001000110011",
16197 => "0000001000110011",
16198 => "0000001000110011",
16199 => "0000001000110100",
16200 => "0000001000110100",
16201 => "0000001000110100",
16202 => "0000001000110100",
16203 => "0000001000110100",
16204 => "0000001000110100",
16205 => "0000001000110100",
16206 => "0000001000110101",
16207 => "0000001000110101",
16208 => "0000001000110101",
16209 => "0000001000110101",
16210 => "0000001000110101",
16211 => "0000001000110101",
16212 => "0000001000110101",
16213 => "0000001000110101",
16214 => "0000001000110110",
16215 => "0000001000110110",
16216 => "0000001000110110",
16217 => "0000001000110110",
16218 => "0000001000110110",
16219 => "0000001000110110",
16220 => "0000001000110110",
16221 => "0000001000110111",
16222 => "0000001000110111",
16223 => "0000001000110111",
16224 => "0000001000110111",
16225 => "0000001000110111",
16226 => "0000001000110111",
16227 => "0000001000110111",
16228 => "0000001000111000",
16229 => "0000001000111000",
16230 => "0000001000111000",
16231 => "0000001000111000",
16232 => "0000001000111000",
16233 => "0000001000111000",
16234 => "0000001000111000",
16235 => "0000001000111000",
16236 => "0000001000111001",
16237 => "0000001000111001",
16238 => "0000001000111001",
16239 => "0000001000111001",
16240 => "0000001000111001",
16241 => "0000001000111001",
16242 => "0000001000111001",
16243 => "0000001000111010",
16244 => "0000001000111010",
16245 => "0000001000111010",
16246 => "0000001000111010",
16247 => "0000001000111010",
16248 => "0000001000111010",
16249 => "0000001000111010",
16250 => "0000001000111011",
16251 => "0000001000111011",
16252 => "0000001000111011",
16253 => "0000001000111011",
16254 => "0000001000111011",
16255 => "0000001000111011",
16256 => "0000001000111011",
16257 => "0000001000111011",
16258 => "0000001000111100",
16259 => "0000001000111100",
16260 => "0000001000111100",
16261 => "0000001000111100",
16262 => "0000001000111100",
16263 => "0000001000111100",
16264 => "0000001000111100",
16265 => "0000001000111101",
16266 => "0000001000111101",
16267 => "0000001000111101",
16268 => "0000001000111101",
16269 => "0000001000111101",
16270 => "0000001000111101",
16271 => "0000001000111101",
16272 => "0000001000111110",
16273 => "0000001000111110",
16274 => "0000001000111110",
16275 => "0000001000111110",
16276 => "0000001000111110",
16277 => "0000001000111110",
16278 => "0000001000111110",
16279 => "0000001000111111",
16280 => "0000001000111111",
16281 => "0000001000111111",
16282 => "0000001000111111",
16283 => "0000001000111111",
16284 => "0000001000111111",
16285 => "0000001000111111",
16286 => "0000001000111111",
16287 => "0000001001000000",
16288 => "0000001001000000",
16289 => "0000001001000000",
16290 => "0000001001000000",
16291 => "0000001001000000",
16292 => "0000001001000000",
16293 => "0000001001000000",
16294 => "0000001001000001",
16295 => "0000001001000001",
16296 => "0000001001000001",
16297 => "0000001001000001",
16298 => "0000001001000001",
16299 => "0000001001000001",
16300 => "0000001001000001",
16301 => "0000001001000010",
16302 => "0000001001000010",
16303 => "0000001001000010",
16304 => "0000001001000010",
16305 => "0000001001000010",
16306 => "0000001001000010",
16307 => "0000001001000010",
16308 => "0000001001000011",
16309 => "0000001001000011",
16310 => "0000001001000011",
16311 => "0000001001000011",
16312 => "0000001001000011",
16313 => "0000001001000011",
16314 => "0000001001000011",
16315 => "0000001001000011",
16316 => "0000001001000100",
16317 => "0000001001000100",
16318 => "0000001001000100",
16319 => "0000001001000100",
16320 => "0000001001000100",
16321 => "0000001001000100",
16322 => "0000001001000100",
16323 => "0000001001000101",
16324 => "0000001001000101",
16325 => "0000001001000101",
16326 => "0000001001000101",
16327 => "0000001001000101",
16328 => "0000001001000101",
16329 => "0000001001000101",
16330 => "0000001001000110",
16331 => "0000001001000110",
16332 => "0000001001000110",
16333 => "0000001001000110",
16334 => "0000001001000110",
16335 => "0000001001000110",
16336 => "0000001001000110",
16337 => "0000001001000111",
16338 => "0000001001000111",
16339 => "0000001001000111",
16340 => "0000001001000111",
16341 => "0000001001000111",
16342 => "0000001001000111",
16343 => "0000001001000111",
16344 => "0000001001001000",
16345 => "0000001001001000",
16346 => "0000001001001000",
16347 => "0000001001001000",
16348 => "0000001001001000",
16349 => "0000001001001000",
16350 => "0000001001001000",
16351 => "0000001001001001",
16352 => "0000001001001001",
16353 => "0000001001001001",
16354 => "0000001001001001",
16355 => "0000001001001001",
16356 => "0000001001001001",
16357 => "0000001001001001",
16358 => "0000001001001001",
16359 => "0000001001001010",
16360 => "0000001001001010",
16361 => "0000001001001010",
16362 => "0000001001001010",
16363 => "0000001001001010",
16364 => "0000001001001010",
16365 => "0000001001001010",
16366 => "0000001001001011",
16367 => "0000001001001011",
16368 => "0000001001001011",
16369 => "0000001001001011",
16370 => "0000001001001011",
16371 => "0000001001001011",
16372 => "0000001001001011",
16373 => "0000001001001100",
16374 => "0000001001001100",
16375 => "0000001001001100",
16376 => "0000001001001100",
16377 => "0000001001001100",
16378 => "0000001001001100",
16379 => "0000001001001100",
16380 => "0000001001001101",
16381 => "0000001001001101",
16382 => "0000001001001101",
16383 => "0000001001001101",
16384 => "0000001001001101",
16385 => "0000001001001101",
16386 => "0000001001001101",
16387 => "0000001001001110",
16388 => "0000001001001110",
16389 => "0000001001001110",
16390 => "0000001001001110",
16391 => "0000001001001110",
16392 => "0000001001001110",
16393 => "0000001001001110",
16394 => "0000001001001111",
16395 => "0000001001001111",
16396 => "0000001001001111",
16397 => "0000001001001111",
16398 => "0000001001001111",
16399 => "0000001001001111",
16400 => "0000001001001111",
16401 => "0000001001010000",
16402 => "0000001001010000",
16403 => "0000001001010000",
16404 => "0000001001010000",
16405 => "0000001001010000",
16406 => "0000001001010000",
16407 => "0000001001010000",
16408 => "0000001001010001",
16409 => "0000001001010001",
16410 => "0000001001010001",
16411 => "0000001001010001",
16412 => "0000001001010001",
16413 => "0000001001010001",
16414 => "0000001001010001",
16415 => "0000001001010010",
16416 => "0000001001010010",
16417 => "0000001001010010",
16418 => "0000001001010010",
16419 => "0000001001010010",
16420 => "0000001001010010",
16421 => "0000001001010010",
16422 => "0000001001010011",
16423 => "0000001001010011",
16424 => "0000001001010011",
16425 => "0000001001010011",
16426 => "0000001001010011",
16427 => "0000001001010011",
16428 => "0000001001010011",
16429 => "0000001001010100",
16430 => "0000001001010100",
16431 => "0000001001010100",
16432 => "0000001001010100",
16433 => "0000001001010100",
16434 => "0000001001010100",
16435 => "0000001001010100",
16436 => "0000001001010101",
16437 => "0000001001010101",
16438 => "0000001001010101",
16439 => "0000001001010101",
16440 => "0000001001010101",
16441 => "0000001001010101",
16442 => "0000001001010101",
16443 => "0000001001010110",
16444 => "0000001001010110",
16445 => "0000001001010110",
16446 => "0000001001010110",
16447 => "0000001001010110",
16448 => "0000001001010110",
16449 => "0000001001010110",
16450 => "0000001001010111",
16451 => "0000001001010111",
16452 => "0000001001010111",
16453 => "0000001001010111",
16454 => "0000001001010111",
16455 => "0000001001010111",
16456 => "0000001001010111",
16457 => "0000001001011000",
16458 => "0000001001011000",
16459 => "0000001001011000",
16460 => "0000001001011000",
16461 => "0000001001011000",
16462 => "0000001001011000",
16463 => "0000001001011000",
16464 => "0000001001011001",
16465 => "0000001001011001",
16466 => "0000001001011001",
16467 => "0000001001011001",
16468 => "0000001001011001",
16469 => "0000001001011001",
16470 => "0000001001011001",
16471 => "0000001001011010",
16472 => "0000001001011010",
16473 => "0000001001011010",
16474 => "0000001001011010",
16475 => "0000001001011010",
16476 => "0000001001011010",
16477 => "0000001001011010",
16478 => "0000001001011011",
16479 => "0000001001011011",
16480 => "0000001001011011",
16481 => "0000001001011011",
16482 => "0000001001011011",
16483 => "0000001001011011",
16484 => "0000001001011011",
16485 => "0000001001011100",
16486 => "0000001001011100",
16487 => "0000001001011100",
16488 => "0000001001011100",
16489 => "0000001001011100",
16490 => "0000001001011100",
16491 => "0000001001011100",
16492 => "0000001001011101",
16493 => "0000001001011101",
16494 => "0000001001011101",
16495 => "0000001001011101",
16496 => "0000001001011101",
16497 => "0000001001011101",
16498 => "0000001001011101",
16499 => "0000001001011110",
16500 => "0000001001011110",
16501 => "0000001001011110",
16502 => "0000001001011110",
16503 => "0000001001011110",
16504 => "0000001001011110",
16505 => "0000001001011111",
16506 => "0000001001011111",
16507 => "0000001001011111",
16508 => "0000001001011111",
16509 => "0000001001011111",
16510 => "0000001001011111",
16511 => "0000001001011111",
16512 => "0000001001100000",
16513 => "0000001001100000",
16514 => "0000001001100000",
16515 => "0000001001100000",
16516 => "0000001001100000",
16517 => "0000001001100000",
16518 => "0000001001100000",
16519 => "0000001001100001",
16520 => "0000001001100001",
16521 => "0000001001100001",
16522 => "0000001001100001",
16523 => "0000001001100001",
16524 => "0000001001100001",
16525 => "0000001001100001",
16526 => "0000001001100010",
16527 => "0000001001100010",
16528 => "0000001001100010",
16529 => "0000001001100010",
16530 => "0000001001100010",
16531 => "0000001001100010",
16532 => "0000001001100010",
16533 => "0000001001100011",
16534 => "0000001001100011",
16535 => "0000001001100011",
16536 => "0000001001100011",
16537 => "0000001001100011",
16538 => "0000001001100011",
16539 => "0000001001100011",
16540 => "0000001001100100",
16541 => "0000001001100100",
16542 => "0000001001100100",
16543 => "0000001001100100",
16544 => "0000001001100100",
16545 => "0000001001100100",
16546 => "0000001001100100",
16547 => "0000001001100101",
16548 => "0000001001100101",
16549 => "0000001001100101",
16550 => "0000001001100101",
16551 => "0000001001100101",
16552 => "0000001001100101",
16553 => "0000001001100110",
16554 => "0000001001100110",
16555 => "0000001001100110",
16556 => "0000001001100110",
16557 => "0000001001100110",
16558 => "0000001001100110",
16559 => "0000001001100110",
16560 => "0000001001100111",
16561 => "0000001001100111",
16562 => "0000001001100111",
16563 => "0000001001100111",
16564 => "0000001001100111",
16565 => "0000001001100111",
16566 => "0000001001100111",
16567 => "0000001001101000",
16568 => "0000001001101000",
16569 => "0000001001101000",
16570 => "0000001001101000",
16571 => "0000001001101000",
16572 => "0000001001101000",
16573 => "0000001001101000",
16574 => "0000001001101001",
16575 => "0000001001101001",
16576 => "0000001001101001",
16577 => "0000001001101001",
16578 => "0000001001101001",
16579 => "0000001001101001",
16580 => "0000001001101010",
16581 => "0000001001101010",
16582 => "0000001001101010",
16583 => "0000001001101010",
16584 => "0000001001101010",
16585 => "0000001001101010",
16586 => "0000001001101010",
16587 => "0000001001101011",
16588 => "0000001001101011",
16589 => "0000001001101011",
16590 => "0000001001101011",
16591 => "0000001001101011",
16592 => "0000001001101011",
16593 => "0000001001101011",
16594 => "0000001001101100",
16595 => "0000001001101100",
16596 => "0000001001101100",
16597 => "0000001001101100",
16598 => "0000001001101100",
16599 => "0000001001101100",
16600 => "0000001001101100",
16601 => "0000001001101101",
16602 => "0000001001101101",
16603 => "0000001001101101",
16604 => "0000001001101101",
16605 => "0000001001101101",
16606 => "0000001001101101",
16607 => "0000001001101110",
16608 => "0000001001101110",
16609 => "0000001001101110",
16610 => "0000001001101110",
16611 => "0000001001101110",
16612 => "0000001001101110",
16613 => "0000001001101110",
16614 => "0000001001101111",
16615 => "0000001001101111",
16616 => "0000001001101111",
16617 => "0000001001101111",
16618 => "0000001001101111",
16619 => "0000001001101111",
16620 => "0000001001101111",
16621 => "0000001001110000",
16622 => "0000001001110000",
16623 => "0000001001110000",
16624 => "0000001001110000",
16625 => "0000001001110000",
16626 => "0000001001110000",
16627 => "0000001001110000",
16628 => "0000001001110001",
16629 => "0000001001110001",
16630 => "0000001001110001",
16631 => "0000001001110001",
16632 => "0000001001110001",
16633 => "0000001001110001",
16634 => "0000001001110010",
16635 => "0000001001110010",
16636 => "0000001001110010",
16637 => "0000001001110010",
16638 => "0000001001110010",
16639 => "0000001001110010",
16640 => "0000001001110010",
16641 => "0000001001110011",
16642 => "0000001001110011",
16643 => "0000001001110011",
16644 => "0000001001110011",
16645 => "0000001001110011",
16646 => "0000001001110011",
16647 => "0000001001110011",
16648 => "0000001001110100",
16649 => "0000001001110100",
16650 => "0000001001110100",
16651 => "0000001001110100",
16652 => "0000001001110100",
16653 => "0000001001110100",
16654 => "0000001001110101",
16655 => "0000001001110101",
16656 => "0000001001110101",
16657 => "0000001001110101",
16658 => "0000001001110101",
16659 => "0000001001110101",
16660 => "0000001001110101",
16661 => "0000001001110110",
16662 => "0000001001110110",
16663 => "0000001001110110",
16664 => "0000001001110110",
16665 => "0000001001110110",
16666 => "0000001001110110",
16667 => "0000001001110111",
16668 => "0000001001110111",
16669 => "0000001001110111",
16670 => "0000001001110111",
16671 => "0000001001110111",
16672 => "0000001001110111",
16673 => "0000001001110111",
16674 => "0000001001111000",
16675 => "0000001001111000",
16676 => "0000001001111000",
16677 => "0000001001111000",
16678 => "0000001001111000",
16679 => "0000001001111000",
16680 => "0000001001111000",
16681 => "0000001001111001",
16682 => "0000001001111001",
16683 => "0000001001111001",
16684 => "0000001001111001",
16685 => "0000001001111001",
16686 => "0000001001111001",
16687 => "0000001001111010",
16688 => "0000001001111010",
16689 => "0000001001111010",
16690 => "0000001001111010",
16691 => "0000001001111010",
16692 => "0000001001111010",
16693 => "0000001001111010",
16694 => "0000001001111011",
16695 => "0000001001111011",
16696 => "0000001001111011",
16697 => "0000001001111011",
16698 => "0000001001111011",
16699 => "0000001001111011",
16700 => "0000001001111100",
16701 => "0000001001111100",
16702 => "0000001001111100",
16703 => "0000001001111100",
16704 => "0000001001111100",
16705 => "0000001001111100",
16706 => "0000001001111100",
16707 => "0000001001111101",
16708 => "0000001001111101",
16709 => "0000001001111101",
16710 => "0000001001111101",
16711 => "0000001001111101",
16712 => "0000001001111101",
16713 => "0000001001111101",
16714 => "0000001001111110",
16715 => "0000001001111110",
16716 => "0000001001111110",
16717 => "0000001001111110",
16718 => "0000001001111110",
16719 => "0000001001111110",
16720 => "0000001001111111",
16721 => "0000001001111111",
16722 => "0000001001111111",
16723 => "0000001001111111",
16724 => "0000001001111111",
16725 => "0000001001111111",
16726 => "0000001001111111",
16727 => "0000001010000000",
16728 => "0000001010000000",
16729 => "0000001010000000",
16730 => "0000001010000000",
16731 => "0000001010000000",
16732 => "0000001010000000",
16733 => "0000001010000001",
16734 => "0000001010000001",
16735 => "0000001010000001",
16736 => "0000001010000001",
16737 => "0000001010000001",
16738 => "0000001010000001",
16739 => "0000001010000001",
16740 => "0000001010000010",
16741 => "0000001010000010",
16742 => "0000001010000010",
16743 => "0000001010000010",
16744 => "0000001010000010",
16745 => "0000001010000010",
16746 => "0000001010000011",
16747 => "0000001010000011",
16748 => "0000001010000011",
16749 => "0000001010000011",
16750 => "0000001010000011",
16751 => "0000001010000011",
16752 => "0000001010000011",
16753 => "0000001010000100",
16754 => "0000001010000100",
16755 => "0000001010000100",
16756 => "0000001010000100",
16757 => "0000001010000100",
16758 => "0000001010000100",
16759 => "0000001010000101",
16760 => "0000001010000101",
16761 => "0000001010000101",
16762 => "0000001010000101",
16763 => "0000001010000101",
16764 => "0000001010000101",
16765 => "0000001010000101",
16766 => "0000001010000110",
16767 => "0000001010000110",
16768 => "0000001010000110",
16769 => "0000001010000110",
16770 => "0000001010000110",
16771 => "0000001010000110",
16772 => "0000001010000111",
16773 => "0000001010000111",
16774 => "0000001010000111",
16775 => "0000001010000111",
16776 => "0000001010000111",
16777 => "0000001010000111",
16778 => "0000001010000111",
16779 => "0000001010001000",
16780 => "0000001010001000",
16781 => "0000001010001000",
16782 => "0000001010001000",
16783 => "0000001010001000",
16784 => "0000001010001000",
16785 => "0000001010001001",
16786 => "0000001010001001",
16787 => "0000001010001001",
16788 => "0000001010001001",
16789 => "0000001010001001",
16790 => "0000001010001001",
16791 => "0000001010001010",
16792 => "0000001010001010",
16793 => "0000001010001010",
16794 => "0000001010001010",
16795 => "0000001010001010",
16796 => "0000001010001010",
16797 => "0000001010001010",
16798 => "0000001010001011",
16799 => "0000001010001011",
16800 => "0000001010001011",
16801 => "0000001010001011",
16802 => "0000001010001011",
16803 => "0000001010001011",
16804 => "0000001010001100",
16805 => "0000001010001100",
16806 => "0000001010001100",
16807 => "0000001010001100",
16808 => "0000001010001100",
16809 => "0000001010001100",
16810 => "0000001010001100",
16811 => "0000001010001101",
16812 => "0000001010001101",
16813 => "0000001010001101",
16814 => "0000001010001101",
16815 => "0000001010001101",
16816 => "0000001010001101",
16817 => "0000001010001110",
16818 => "0000001010001110",
16819 => "0000001010001110",
16820 => "0000001010001110",
16821 => "0000001010001110",
16822 => "0000001010001110",
16823 => "0000001010001111",
16824 => "0000001010001111",
16825 => "0000001010001111",
16826 => "0000001010001111",
16827 => "0000001010001111",
16828 => "0000001010001111",
16829 => "0000001010001111",
16830 => "0000001010010000",
16831 => "0000001010010000",
16832 => "0000001010010000",
16833 => "0000001010010000",
16834 => "0000001010010000",
16835 => "0000001010010000",
16836 => "0000001010010001",
16837 => "0000001010010001",
16838 => "0000001010010001",
16839 => "0000001010010001",
16840 => "0000001010010001",
16841 => "0000001010010001",
16842 => "0000001010010001",
16843 => "0000001010010010",
16844 => "0000001010010010",
16845 => "0000001010010010",
16846 => "0000001010010010",
16847 => "0000001010010010",
16848 => "0000001010010010",
16849 => "0000001010010011",
16850 => "0000001010010011",
16851 => "0000001010010011",
16852 => "0000001010010011",
16853 => "0000001010010011",
16854 => "0000001010010011",
16855 => "0000001010010100",
16856 => "0000001010010100",
16857 => "0000001010010100",
16858 => "0000001010010100",
16859 => "0000001010010100",
16860 => "0000001010010100",
16861 => "0000001010010100",
16862 => "0000001010010101",
16863 => "0000001010010101",
16864 => "0000001010010101",
16865 => "0000001010010101",
16866 => "0000001010010101",
16867 => "0000001010010101",
16868 => "0000001010010110",
16869 => "0000001010010110",
16870 => "0000001010010110",
16871 => "0000001010010110",
16872 => "0000001010010110",
16873 => "0000001010010110",
16874 => "0000001010010111",
16875 => "0000001010010111",
16876 => "0000001010010111",
16877 => "0000001010010111",
16878 => "0000001010010111",
16879 => "0000001010010111",
16880 => "0000001010010111",
16881 => "0000001010011000",
16882 => "0000001010011000",
16883 => "0000001010011000",
16884 => "0000001010011000",
16885 => "0000001010011000",
16886 => "0000001010011000",
16887 => "0000001010011001",
16888 => "0000001010011001",
16889 => "0000001010011001",
16890 => "0000001010011001",
16891 => "0000001010011001",
16892 => "0000001010011001",
16893 => "0000001010011010",
16894 => "0000001010011010",
16895 => "0000001010011010",
16896 => "0000001010011010",
16897 => "0000001010011010",
16898 => "0000001010011010",
16899 => "0000001010011011",
16900 => "0000001010011011",
16901 => "0000001010011011",
16902 => "0000001010011011",
16903 => "0000001010011011",
16904 => "0000001010011011",
16905 => "0000001010011011",
16906 => "0000001010011100",
16907 => "0000001010011100",
16908 => "0000001010011100",
16909 => "0000001010011100",
16910 => "0000001010011100",
16911 => "0000001010011100",
16912 => "0000001010011101",
16913 => "0000001010011101",
16914 => "0000001010011101",
16915 => "0000001010011101",
16916 => "0000001010011101",
16917 => "0000001010011101",
16918 => "0000001010011110",
16919 => "0000001010011110",
16920 => "0000001010011110",
16921 => "0000001010011110",
16922 => "0000001010011110",
16923 => "0000001010011110",
16924 => "0000001010011111",
16925 => "0000001010011111",
16926 => "0000001010011111",
16927 => "0000001010011111",
16928 => "0000001010011111",
16929 => "0000001010011111",
16930 => "0000001010011111",
16931 => "0000001010100000",
16932 => "0000001010100000",
16933 => "0000001010100000",
16934 => "0000001010100000",
16935 => "0000001010100000",
16936 => "0000001010100000",
16937 => "0000001010100001",
16938 => "0000001010100001",
16939 => "0000001010100001",
16940 => "0000001010100001",
16941 => "0000001010100001",
16942 => "0000001010100001",
16943 => "0000001010100010",
16944 => "0000001010100010",
16945 => "0000001010100010",
16946 => "0000001010100010",
16947 => "0000001010100010",
16948 => "0000001010100010",
16949 => "0000001010100011",
16950 => "0000001010100011",
16951 => "0000001010100011",
16952 => "0000001010100011",
16953 => "0000001010100011",
16954 => "0000001010100011",
16955 => "0000001010100100",
16956 => "0000001010100100",
16957 => "0000001010100100",
16958 => "0000001010100100",
16959 => "0000001010100100",
16960 => "0000001010100100",
16961 => "0000001010100100",
16962 => "0000001010100101",
16963 => "0000001010100101",
16964 => "0000001010100101",
16965 => "0000001010100101",
16966 => "0000001010100101",
16967 => "0000001010100101",
16968 => "0000001010100110",
16969 => "0000001010100110",
16970 => "0000001010100110",
16971 => "0000001010100110",
16972 => "0000001010100110",
16973 => "0000001010100110",
16974 => "0000001010100111",
16975 => "0000001010100111",
16976 => "0000001010100111",
16977 => "0000001010100111",
16978 => "0000001010100111",
16979 => "0000001010100111",
16980 => "0000001010101000",
16981 => "0000001010101000",
16982 => "0000001010101000",
16983 => "0000001010101000",
16984 => "0000001010101000",
16985 => "0000001010101000",
16986 => "0000001010101001",
16987 => "0000001010101001",
16988 => "0000001010101001",
16989 => "0000001010101001",
16990 => "0000001010101001",
16991 => "0000001010101001",
16992 => "0000001010101010",
16993 => "0000001010101010",
16994 => "0000001010101010",
16995 => "0000001010101010",
16996 => "0000001010101010",
16997 => "0000001010101010",
16998 => "0000001010101010",
16999 => "0000001010101011",
17000 => "0000001010101011",
17001 => "0000001010101011",
17002 => "0000001010101011",
17003 => "0000001010101011",
17004 => "0000001010101011",
17005 => "0000001010101100",
17006 => "0000001010101100",
17007 => "0000001010101100",
17008 => "0000001010101100",
17009 => "0000001010101100",
17010 => "0000001010101100",
17011 => "0000001010101101",
17012 => "0000001010101101",
17013 => "0000001010101101",
17014 => "0000001010101101",
17015 => "0000001010101101",
17016 => "0000001010101101",
17017 => "0000001010101110",
17018 => "0000001010101110",
17019 => "0000001010101110",
17020 => "0000001010101110",
17021 => "0000001010101110",
17022 => "0000001010101110",
17023 => "0000001010101111",
17024 => "0000001010101111",
17025 => "0000001010101111",
17026 => "0000001010101111",
17027 => "0000001010101111",
17028 => "0000001010101111",
17029 => "0000001010110000",
17030 => "0000001010110000",
17031 => "0000001010110000",
17032 => "0000001010110000",
17033 => "0000001010110000",
17034 => "0000001010110000",
17035 => "0000001010110001",
17036 => "0000001010110001",
17037 => "0000001010110001",
17038 => "0000001010110001",
17039 => "0000001010110001",
17040 => "0000001010110001",
17041 => "0000001010110010",
17042 => "0000001010110010",
17043 => "0000001010110010",
17044 => "0000001010110010",
17045 => "0000001010110010",
17046 => "0000001010110010",
17047 => "0000001010110011",
17048 => "0000001010110011",
17049 => "0000001010110011",
17050 => "0000001010110011",
17051 => "0000001010110011",
17052 => "0000001010110011",
17053 => "0000001010110100",
17054 => "0000001010110100",
17055 => "0000001010110100",
17056 => "0000001010110100",
17057 => "0000001010110100",
17058 => "0000001010110100",
17059 => "0000001010110101",
17060 => "0000001010110101",
17061 => "0000001010110101",
17062 => "0000001010110101",
17063 => "0000001010110101",
17064 => "0000001010110101",
17065 => "0000001010110110",
17066 => "0000001010110110",
17067 => "0000001010110110",
17068 => "0000001010110110",
17069 => "0000001010110110",
17070 => "0000001010110110",
17071 => "0000001010110111",
17072 => "0000001010110111",
17073 => "0000001010110111",
17074 => "0000001010110111",
17075 => "0000001010110111",
17076 => "0000001010110111",
17077 => "0000001010111000",
17078 => "0000001010111000",
17079 => "0000001010111000",
17080 => "0000001010111000",
17081 => "0000001010111000",
17082 => "0000001010111000",
17083 => "0000001010111001",
17084 => "0000001010111001",
17085 => "0000001010111001",
17086 => "0000001010111001",
17087 => "0000001010111001",
17088 => "0000001010111001",
17089 => "0000001010111010",
17090 => "0000001010111010",
17091 => "0000001010111010",
17092 => "0000001010111010",
17093 => "0000001010111010",
17094 => "0000001010111010",
17095 => "0000001010111011",
17096 => "0000001010111011",
17097 => "0000001010111011",
17098 => "0000001010111011",
17099 => "0000001010111011",
17100 => "0000001010111011",
17101 => "0000001010111100",
17102 => "0000001010111100",
17103 => "0000001010111100",
17104 => "0000001010111100",
17105 => "0000001010111100",
17106 => "0000001010111100",
17107 => "0000001010111101",
17108 => "0000001010111101",
17109 => "0000001010111101",
17110 => "0000001010111101",
17111 => "0000001010111101",
17112 => "0000001010111101",
17113 => "0000001010111110",
17114 => "0000001010111110",
17115 => "0000001010111110",
17116 => "0000001010111110",
17117 => "0000001010111110",
17118 => "0000001010111110",
17119 => "0000001010111111",
17120 => "0000001010111111",
17121 => "0000001010111111",
17122 => "0000001010111111",
17123 => "0000001010111111",
17124 => "0000001010111111",
17125 => "0000001011000000",
17126 => "0000001011000000",
17127 => "0000001011000000",
17128 => "0000001011000000",
17129 => "0000001011000000",
17130 => "0000001011000000",
17131 => "0000001011000001",
17132 => "0000001011000001",
17133 => "0000001011000001",
17134 => "0000001011000001",
17135 => "0000001011000001",
17136 => "0000001011000001",
17137 => "0000001011000010",
17138 => "0000001011000010",
17139 => "0000001011000010",
17140 => "0000001011000010",
17141 => "0000001011000010",
17142 => "0000001011000010",
17143 => "0000001011000011",
17144 => "0000001011000011",
17145 => "0000001011000011",
17146 => "0000001011000011",
17147 => "0000001011000011",
17148 => "0000001011000011",
17149 => "0000001011000100",
17150 => "0000001011000100",
17151 => "0000001011000100",
17152 => "0000001011000100",
17153 => "0000001011000100",
17154 => "0000001011000100",
17155 => "0000001011000101",
17156 => "0000001011000101",
17157 => "0000001011000101",
17158 => "0000001011000101",
17159 => "0000001011000101",
17160 => "0000001011000101",
17161 => "0000001011000110",
17162 => "0000001011000110",
17163 => "0000001011000110",
17164 => "0000001011000110",
17165 => "0000001011000110",
17166 => "0000001011000110",
17167 => "0000001011000111",
17168 => "0000001011000111",
17169 => "0000001011000111",
17170 => "0000001011000111",
17171 => "0000001011000111",
17172 => "0000001011000111",
17173 => "0000001011001000",
17174 => "0000001011001000",
17175 => "0000001011001000",
17176 => "0000001011001000",
17177 => "0000001011001000",
17178 => "0000001011001000",
17179 => "0000001011001001",
17180 => "0000001011001001",
17181 => "0000001011001001",
17182 => "0000001011001001",
17183 => "0000001011001001",
17184 => "0000001011001010",
17185 => "0000001011001010",
17186 => "0000001011001010",
17187 => "0000001011001010",
17188 => "0000001011001010",
17189 => "0000001011001010",
17190 => "0000001011001011",
17191 => "0000001011001011",
17192 => "0000001011001011",
17193 => "0000001011001011",
17194 => "0000001011001011",
17195 => "0000001011001011",
17196 => "0000001011001100",
17197 => "0000001011001100",
17198 => "0000001011001100",
17199 => "0000001011001100",
17200 => "0000001011001100",
17201 => "0000001011001100",
17202 => "0000001011001101",
17203 => "0000001011001101",
17204 => "0000001011001101",
17205 => "0000001011001101",
17206 => "0000001011001101",
17207 => "0000001011001101",
17208 => "0000001011001110",
17209 => "0000001011001110",
17210 => "0000001011001110",
17211 => "0000001011001110",
17212 => "0000001011001110",
17213 => "0000001011001110",
17214 => "0000001011001111",
17215 => "0000001011001111",
17216 => "0000001011001111",
17217 => "0000001011001111",
17218 => "0000001011001111",
17219 => "0000001011010000",
17220 => "0000001011010000",
17221 => "0000001011010000",
17222 => "0000001011010000",
17223 => "0000001011010000",
17224 => "0000001011010000",
17225 => "0000001011010001",
17226 => "0000001011010001",
17227 => "0000001011010001",
17228 => "0000001011010001",
17229 => "0000001011010001",
17230 => "0000001011010001",
17231 => "0000001011010010",
17232 => "0000001011010010",
17233 => "0000001011010010",
17234 => "0000001011010010",
17235 => "0000001011010010",
17236 => "0000001011010010",
17237 => "0000001011010011",
17238 => "0000001011010011",
17239 => "0000001011010011",
17240 => "0000001011010011",
17241 => "0000001011010011",
17242 => "0000001011010011",
17243 => "0000001011010100",
17244 => "0000001011010100",
17245 => "0000001011010100",
17246 => "0000001011010100",
17247 => "0000001011010100",
17248 => "0000001011010101",
17249 => "0000001011010101",
17250 => "0000001011010101",
17251 => "0000001011010101",
17252 => "0000001011010101",
17253 => "0000001011010101",
17254 => "0000001011010110",
17255 => "0000001011010110",
17256 => "0000001011010110",
17257 => "0000001011010110",
17258 => "0000001011010110",
17259 => "0000001011010110",
17260 => "0000001011010111",
17261 => "0000001011010111",
17262 => "0000001011010111",
17263 => "0000001011010111",
17264 => "0000001011010111",
17265 => "0000001011010111",
17266 => "0000001011011000",
17267 => "0000001011011000",
17268 => "0000001011011000",
17269 => "0000001011011000",
17270 => "0000001011011000",
17271 => "0000001011011001",
17272 => "0000001011011001",
17273 => "0000001011011001",
17274 => "0000001011011001",
17275 => "0000001011011001",
17276 => "0000001011011001",
17277 => "0000001011011010",
17278 => "0000001011011010",
17279 => "0000001011011010",
17280 => "0000001011011010",
17281 => "0000001011011010",
17282 => "0000001011011010",
17283 => "0000001011011011",
17284 => "0000001011011011",
17285 => "0000001011011011",
17286 => "0000001011011011",
17287 => "0000001011011011",
17288 => "0000001011011011",
17289 => "0000001011011100",
17290 => "0000001011011100",
17291 => "0000001011011100",
17292 => "0000001011011100",
17293 => "0000001011011100",
17294 => "0000001011011101",
17295 => "0000001011011101",
17296 => "0000001011011101",
17297 => "0000001011011101",
17298 => "0000001011011101",
17299 => "0000001011011101",
17300 => "0000001011011110",
17301 => "0000001011011110",
17302 => "0000001011011110",
17303 => "0000001011011110",
17304 => "0000001011011110",
17305 => "0000001011011110",
17306 => "0000001011011111",
17307 => "0000001011011111",
17308 => "0000001011011111",
17309 => "0000001011011111",
17310 => "0000001011011111",
17311 => "0000001011011111",
17312 => "0000001011100000",
17313 => "0000001011100000",
17314 => "0000001011100000",
17315 => "0000001011100000",
17316 => "0000001011100000",
17317 => "0000001011100001",
17318 => "0000001011100001",
17319 => "0000001011100001",
17320 => "0000001011100001",
17321 => "0000001011100001",
17322 => "0000001011100001",
17323 => "0000001011100010",
17324 => "0000001011100010",
17325 => "0000001011100010",
17326 => "0000001011100010",
17327 => "0000001011100010",
17328 => "0000001011100010",
17329 => "0000001011100011",
17330 => "0000001011100011",
17331 => "0000001011100011",
17332 => "0000001011100011",
17333 => "0000001011100011",
17334 => "0000001011100100",
17335 => "0000001011100100",
17336 => "0000001011100100",
17337 => "0000001011100100",
17338 => "0000001011100100",
17339 => "0000001011100100",
17340 => "0000001011100101",
17341 => "0000001011100101",
17342 => "0000001011100101",
17343 => "0000001011100101",
17344 => "0000001011100101",
17345 => "0000001011100101",
17346 => "0000001011100110",
17347 => "0000001011100110",
17348 => "0000001011100110",
17349 => "0000001011100110",
17350 => "0000001011100110",
17351 => "0000001011100111",
17352 => "0000001011100111",
17353 => "0000001011100111",
17354 => "0000001011100111",
17355 => "0000001011100111",
17356 => "0000001011100111",
17357 => "0000001011101000",
17358 => "0000001011101000",
17359 => "0000001011101000",
17360 => "0000001011101000",
17361 => "0000001011101000",
17362 => "0000001011101001",
17363 => "0000001011101001",
17364 => "0000001011101001",
17365 => "0000001011101001",
17366 => "0000001011101001",
17367 => "0000001011101001",
17368 => "0000001011101010",
17369 => "0000001011101010",
17370 => "0000001011101010",
17371 => "0000001011101010",
17372 => "0000001011101010",
17373 => "0000001011101010",
17374 => "0000001011101011",
17375 => "0000001011101011",
17376 => "0000001011101011",
17377 => "0000001011101011",
17378 => "0000001011101011",
17379 => "0000001011101100",
17380 => "0000001011101100",
17381 => "0000001011101100",
17382 => "0000001011101100",
17383 => "0000001011101100",
17384 => "0000001011101100",
17385 => "0000001011101101",
17386 => "0000001011101101",
17387 => "0000001011101101",
17388 => "0000001011101101",
17389 => "0000001011101101",
17390 => "0000001011101101",
17391 => "0000001011101110",
17392 => "0000001011101110",
17393 => "0000001011101110",
17394 => "0000001011101110",
17395 => "0000001011101110",
17396 => "0000001011101111",
17397 => "0000001011101111",
17398 => "0000001011101111",
17399 => "0000001011101111",
17400 => "0000001011101111",
17401 => "0000001011101111",
17402 => "0000001011110000",
17403 => "0000001011110000",
17404 => "0000001011110000",
17405 => "0000001011110000",
17406 => "0000001011110000",
17407 => "0000001011110001",
17408 => "0000001011110001",
17409 => "0000001011110001",
17410 => "0000001011110001",
17411 => "0000001011110001",
17412 => "0000001011110001",
17413 => "0000001011110010",
17414 => "0000001011110010",
17415 => "0000001011110010",
17416 => "0000001011110010",
17417 => "0000001011110010",
17418 => "0000001011110011",
17419 => "0000001011110011",
17420 => "0000001011110011",
17421 => "0000001011110011",
17422 => "0000001011110011",
17423 => "0000001011110011",
17424 => "0000001011110100",
17425 => "0000001011110100",
17426 => "0000001011110100",
17427 => "0000001011110100",
17428 => "0000001011110100",
17429 => "0000001011110101",
17430 => "0000001011110101",
17431 => "0000001011110101",
17432 => "0000001011110101",
17433 => "0000001011110101",
17434 => "0000001011110101",
17435 => "0000001011110110",
17436 => "0000001011110110",
17437 => "0000001011110110",
17438 => "0000001011110110",
17439 => "0000001011110110",
17440 => "0000001011110110",
17441 => "0000001011110111",
17442 => "0000001011110111",
17443 => "0000001011110111",
17444 => "0000001011110111",
17445 => "0000001011110111",
17446 => "0000001011111000",
17447 => "0000001011111000",
17448 => "0000001011111000",
17449 => "0000001011111000",
17450 => "0000001011111000",
17451 => "0000001011111000",
17452 => "0000001011111001",
17453 => "0000001011111001",
17454 => "0000001011111001",
17455 => "0000001011111001",
17456 => "0000001011111001",
17457 => "0000001011111010",
17458 => "0000001011111010",
17459 => "0000001011111010",
17460 => "0000001011111010",
17461 => "0000001011111010",
17462 => "0000001011111010",
17463 => "0000001011111011",
17464 => "0000001011111011",
17465 => "0000001011111011",
17466 => "0000001011111011",
17467 => "0000001011111011",
17468 => "0000001011111100",
17469 => "0000001011111100",
17470 => "0000001011111100",
17471 => "0000001011111100",
17472 => "0000001011111100",
17473 => "0000001011111100",
17474 => "0000001011111101",
17475 => "0000001011111101",
17476 => "0000001011111101",
17477 => "0000001011111101",
17478 => "0000001011111101",
17479 => "0000001011111110",
17480 => "0000001011111110",
17481 => "0000001011111110",
17482 => "0000001011111110",
17483 => "0000001011111110",
17484 => "0000001011111110",
17485 => "0000001011111111",
17486 => "0000001011111111",
17487 => "0000001011111111",
17488 => "0000001011111111",
17489 => "0000001011111111",
17490 => "0000001100000000",
17491 => "0000001100000000",
17492 => "0000001100000000",
17493 => "0000001100000000",
17494 => "0000001100000000",
17495 => "0000001100000001",
17496 => "0000001100000001",
17497 => "0000001100000001",
17498 => "0000001100000001",
17499 => "0000001100000001",
17500 => "0000001100000001",
17501 => "0000001100000010",
17502 => "0000001100000010",
17503 => "0000001100000010",
17504 => "0000001100000010",
17505 => "0000001100000010",
17506 => "0000001100000011",
17507 => "0000001100000011",
17508 => "0000001100000011",
17509 => "0000001100000011",
17510 => "0000001100000011",
17511 => "0000001100000011",
17512 => "0000001100000100",
17513 => "0000001100000100",
17514 => "0000001100000100",
17515 => "0000001100000100",
17516 => "0000001100000100",
17517 => "0000001100000101",
17518 => "0000001100000101",
17519 => "0000001100000101",
17520 => "0000001100000101",
17521 => "0000001100000101",
17522 => "0000001100000101",
17523 => "0000001100000110",
17524 => "0000001100000110",
17525 => "0000001100000110",
17526 => "0000001100000110",
17527 => "0000001100000110",
17528 => "0000001100000111",
17529 => "0000001100000111",
17530 => "0000001100000111",
17531 => "0000001100000111",
17532 => "0000001100000111",
17533 => "0000001100001000",
17534 => "0000001100001000",
17535 => "0000001100001000",
17536 => "0000001100001000",
17537 => "0000001100001000",
17538 => "0000001100001000",
17539 => "0000001100001001",
17540 => "0000001100001001",
17541 => "0000001100001001",
17542 => "0000001100001001",
17543 => "0000001100001001",
17544 => "0000001100001010",
17545 => "0000001100001010",
17546 => "0000001100001010",
17547 => "0000001100001010",
17548 => "0000001100001010",
17549 => "0000001100001010",
17550 => "0000001100001011",
17551 => "0000001100001011",
17552 => "0000001100001011",
17553 => "0000001100001011",
17554 => "0000001100001011",
17555 => "0000001100001100",
17556 => "0000001100001100",
17557 => "0000001100001100",
17558 => "0000001100001100",
17559 => "0000001100001100",
17560 => "0000001100001101",
17561 => "0000001100001101",
17562 => "0000001100001101",
17563 => "0000001100001101",
17564 => "0000001100001101",
17565 => "0000001100001101",
17566 => "0000001100001110",
17567 => "0000001100001110",
17568 => "0000001100001110",
17569 => "0000001100001110",
17570 => "0000001100001110",
17571 => "0000001100001111",
17572 => "0000001100001111",
17573 => "0000001100001111",
17574 => "0000001100001111",
17575 => "0000001100001111",
17576 => "0000001100001111",
17577 => "0000001100010000",
17578 => "0000001100010000",
17579 => "0000001100010000",
17580 => "0000001100010000",
17581 => "0000001100010000",
17582 => "0000001100010001",
17583 => "0000001100010001",
17584 => "0000001100010001",
17585 => "0000001100010001",
17586 => "0000001100010001",
17587 => "0000001100010010",
17588 => "0000001100010010",
17589 => "0000001100010010",
17590 => "0000001100010010",
17591 => "0000001100010010",
17592 => "0000001100010010",
17593 => "0000001100010011",
17594 => "0000001100010011",
17595 => "0000001100010011",
17596 => "0000001100010011",
17597 => "0000001100010011",
17598 => "0000001100010100",
17599 => "0000001100010100",
17600 => "0000001100010100",
17601 => "0000001100010100",
17602 => "0000001100010100",
17603 => "0000001100010101",
17604 => "0000001100010101",
17605 => "0000001100010101",
17606 => "0000001100010101",
17607 => "0000001100010101",
17608 => "0000001100010101",
17609 => "0000001100010110",
17610 => "0000001100010110",
17611 => "0000001100010110",
17612 => "0000001100010110",
17613 => "0000001100010110",
17614 => "0000001100010111",
17615 => "0000001100010111",
17616 => "0000001100010111",
17617 => "0000001100010111",
17618 => "0000001100010111",
17619 => "0000001100011000",
17620 => "0000001100011000",
17621 => "0000001100011000",
17622 => "0000001100011000",
17623 => "0000001100011000",
17624 => "0000001100011001",
17625 => "0000001100011001",
17626 => "0000001100011001",
17627 => "0000001100011001",
17628 => "0000001100011001",
17629 => "0000001100011001",
17630 => "0000001100011010",
17631 => "0000001100011010",
17632 => "0000001100011010",
17633 => "0000001100011010",
17634 => "0000001100011010",
17635 => "0000001100011011",
17636 => "0000001100011011",
17637 => "0000001100011011",
17638 => "0000001100011011",
17639 => "0000001100011011",
17640 => "0000001100011100",
17641 => "0000001100011100",
17642 => "0000001100011100",
17643 => "0000001100011100",
17644 => "0000001100011100",
17645 => "0000001100011100",
17646 => "0000001100011101",
17647 => "0000001100011101",
17648 => "0000001100011101",
17649 => "0000001100011101",
17650 => "0000001100011101",
17651 => "0000001100011110",
17652 => "0000001100011110",
17653 => "0000001100011110",
17654 => "0000001100011110",
17655 => "0000001100011110",
17656 => "0000001100011111",
17657 => "0000001100011111",
17658 => "0000001100011111",
17659 => "0000001100011111",
17660 => "0000001100011111",
17661 => "0000001100100000",
17662 => "0000001100100000",
17663 => "0000001100100000",
17664 => "0000001100100000",
17665 => "0000001100100000",
17666 => "0000001100100000",
17667 => "0000001100100001",
17668 => "0000001100100001",
17669 => "0000001100100001",
17670 => "0000001100100001",
17671 => "0000001100100001",
17672 => "0000001100100010",
17673 => "0000001100100010",
17674 => "0000001100100010",
17675 => "0000001100100010",
17676 => "0000001100100010",
17677 => "0000001100100011",
17678 => "0000001100100011",
17679 => "0000001100100011",
17680 => "0000001100100011",
17681 => "0000001100100011",
17682 => "0000001100100100",
17683 => "0000001100100100",
17684 => "0000001100100100",
17685 => "0000001100100100",
17686 => "0000001100100100",
17687 => "0000001100100100",
17688 => "0000001100100101",
17689 => "0000001100100101",
17690 => "0000001100100101",
17691 => "0000001100100101",
17692 => "0000001100100101",
17693 => "0000001100100110",
17694 => "0000001100100110",
17695 => "0000001100100110",
17696 => "0000001100100110",
17697 => "0000001100100110",
17698 => "0000001100100111",
17699 => "0000001100100111",
17700 => "0000001100100111",
17701 => "0000001100100111",
17702 => "0000001100100111",
17703 => "0000001100101000",
17704 => "0000001100101000",
17705 => "0000001100101000",
17706 => "0000001100101000",
17707 => "0000001100101000",
17708 => "0000001100101001",
17709 => "0000001100101001",
17710 => "0000001100101001",
17711 => "0000001100101001",
17712 => "0000001100101001",
17713 => "0000001100101001",
17714 => "0000001100101010",
17715 => "0000001100101010",
17716 => "0000001100101010",
17717 => "0000001100101010",
17718 => "0000001100101010",
17719 => "0000001100101011",
17720 => "0000001100101011",
17721 => "0000001100101011",
17722 => "0000001100101011",
17723 => "0000001100101011",
17724 => "0000001100101100",
17725 => "0000001100101100",
17726 => "0000001100101100",
17727 => "0000001100101100",
17728 => "0000001100101100",
17729 => "0000001100101101",
17730 => "0000001100101101",
17731 => "0000001100101101",
17732 => "0000001100101101",
17733 => "0000001100101101",
17734 => "0000001100101110",
17735 => "0000001100101110",
17736 => "0000001100101110",
17737 => "0000001100101110",
17738 => "0000001100101110",
17739 => "0000001100101111",
17740 => "0000001100101111",
17741 => "0000001100101111",
17742 => "0000001100101111",
17743 => "0000001100101111",
17744 => "0000001100101111",
17745 => "0000001100110000",
17746 => "0000001100110000",
17747 => "0000001100110000",
17748 => "0000001100110000",
17749 => "0000001100110000",
17750 => "0000001100110001",
17751 => "0000001100110001",
17752 => "0000001100110001",
17753 => "0000001100110001",
17754 => "0000001100110001",
17755 => "0000001100110010",
17756 => "0000001100110010",
17757 => "0000001100110010",
17758 => "0000001100110010",
17759 => "0000001100110010",
17760 => "0000001100110011",
17761 => "0000001100110011",
17762 => "0000001100110011",
17763 => "0000001100110011",
17764 => "0000001100110011",
17765 => "0000001100110100",
17766 => "0000001100110100",
17767 => "0000001100110100",
17768 => "0000001100110100",
17769 => "0000001100110100",
17770 => "0000001100110101",
17771 => "0000001100110101",
17772 => "0000001100110101",
17773 => "0000001100110101",
17774 => "0000001100110101",
17775 => "0000001100110110",
17776 => "0000001100110110",
17777 => "0000001100110110",
17778 => "0000001100110110",
17779 => "0000001100110110",
17780 => "0000001100110111",
17781 => "0000001100110111",
17782 => "0000001100110111",
17783 => "0000001100110111",
17784 => "0000001100110111",
17785 => "0000001100110111",
17786 => "0000001100111000",
17787 => "0000001100111000",
17788 => "0000001100111000",
17789 => "0000001100111000",
17790 => "0000001100111000",
17791 => "0000001100111001",
17792 => "0000001100111001",
17793 => "0000001100111001",
17794 => "0000001100111001",
17795 => "0000001100111001",
17796 => "0000001100111010",
17797 => "0000001100111010",
17798 => "0000001100111010",
17799 => "0000001100111010",
17800 => "0000001100111010",
17801 => "0000001100111011",
17802 => "0000001100111011",
17803 => "0000001100111011",
17804 => "0000001100111011",
17805 => "0000001100111011",
17806 => "0000001100111100",
17807 => "0000001100111100",
17808 => "0000001100111100",
17809 => "0000001100111100",
17810 => "0000001100111100",
17811 => "0000001100111101",
17812 => "0000001100111101",
17813 => "0000001100111101",
17814 => "0000001100111101",
17815 => "0000001100111101",
17816 => "0000001100111110",
17817 => "0000001100111110",
17818 => "0000001100111110",
17819 => "0000001100111110",
17820 => "0000001100111110",
17821 => "0000001100111111",
17822 => "0000001100111111",
17823 => "0000001100111111",
17824 => "0000001100111111",
17825 => "0000001100111111",
17826 => "0000001101000000",
17827 => "0000001101000000",
17828 => "0000001101000000",
17829 => "0000001101000000",
17830 => "0000001101000000",
17831 => "0000001101000001",
17832 => "0000001101000001",
17833 => "0000001101000001",
17834 => "0000001101000001",
17835 => "0000001101000001",
17836 => "0000001101000010",
17837 => "0000001101000010",
17838 => "0000001101000010",
17839 => "0000001101000010",
17840 => "0000001101000010",
17841 => "0000001101000011",
17842 => "0000001101000011",
17843 => "0000001101000011",
17844 => "0000001101000011",
17845 => "0000001101000011",
17846 => "0000001101000100",
17847 => "0000001101000100",
17848 => "0000001101000100",
17849 => "0000001101000100",
17850 => "0000001101000100",
17851 => "0000001101000101",
17852 => "0000001101000101",
17853 => "0000001101000101",
17854 => "0000001101000101",
17855 => "0000001101000101",
17856 => "0000001101000110",
17857 => "0000001101000110",
17858 => "0000001101000110",
17859 => "0000001101000110",
17860 => "0000001101000110",
17861 => "0000001101000111",
17862 => "0000001101000111",
17863 => "0000001101000111",
17864 => "0000001101000111",
17865 => "0000001101000111",
17866 => "0000001101001000",
17867 => "0000001101001000",
17868 => "0000001101001000",
17869 => "0000001101001000",
17870 => "0000001101001000",
17871 => "0000001101001001",
17872 => "0000001101001001",
17873 => "0000001101001001",
17874 => "0000001101001001",
17875 => "0000001101001001",
17876 => "0000001101001010",
17877 => "0000001101001010",
17878 => "0000001101001010",
17879 => "0000001101001010",
17880 => "0000001101001010",
17881 => "0000001101001011",
17882 => "0000001101001011",
17883 => "0000001101001011",
17884 => "0000001101001011",
17885 => "0000001101001011",
17886 => "0000001101001100",
17887 => "0000001101001100",
17888 => "0000001101001100",
17889 => "0000001101001100",
17890 => "0000001101001100",
17891 => "0000001101001101",
17892 => "0000001101001101",
17893 => "0000001101001101",
17894 => "0000001101001101",
17895 => "0000001101001101",
17896 => "0000001101001110",
17897 => "0000001101001110",
17898 => "0000001101001110",
17899 => "0000001101001110",
17900 => "0000001101001110",
17901 => "0000001101001111",
17902 => "0000001101001111",
17903 => "0000001101001111",
17904 => "0000001101001111",
17905 => "0000001101001111",
17906 => "0000001101010000",
17907 => "0000001101010000",
17908 => "0000001101010000",
17909 => "0000001101010000",
17910 => "0000001101010000",
17911 => "0000001101010001",
17912 => "0000001101010001",
17913 => "0000001101010001",
17914 => "0000001101010001",
17915 => "0000001101010001",
17916 => "0000001101010010",
17917 => "0000001101010010",
17918 => "0000001101010010",
17919 => "0000001101010010",
17920 => "0000001101010010",
17921 => "0000001101010011",
17922 => "0000001101010011",
17923 => "0000001101010011",
17924 => "0000001101010011",
17925 => "0000001101010011",
17926 => "0000001101010100",
17927 => "0000001101010100",
17928 => "0000001101010100",
17929 => "0000001101010100",
17930 => "0000001101010100",
17931 => "0000001101010101",
17932 => "0000001101010101",
17933 => "0000001101010101",
17934 => "0000001101010101",
17935 => "0000001101010101",
17936 => "0000001101010110",
17937 => "0000001101010110",
17938 => "0000001101010110",
17939 => "0000001101010110",
17940 => "0000001101010110",
17941 => "0000001101010111",
17942 => "0000001101010111",
17943 => "0000001101010111",
17944 => "0000001101010111",
17945 => "0000001101010111",
17946 => "0000001101011000",
17947 => "0000001101011000",
17948 => "0000001101011000",
17949 => "0000001101011000",
17950 => "0000001101011000",
17951 => "0000001101011001",
17952 => "0000001101011001",
17953 => "0000001101011001",
17954 => "0000001101011001",
17955 => "0000001101011001",
17956 => "0000001101011010",
17957 => "0000001101011010",
17958 => "0000001101011010",
17959 => "0000001101011010",
17960 => "0000001101011011",
17961 => "0000001101011011",
17962 => "0000001101011011",
17963 => "0000001101011011",
17964 => "0000001101011011",
17965 => "0000001101011100",
17966 => "0000001101011100",
17967 => "0000001101011100",
17968 => "0000001101011100",
17969 => "0000001101011100",
17970 => "0000001101011101",
17971 => "0000001101011101",
17972 => "0000001101011101",
17973 => "0000001101011101",
17974 => "0000001101011101",
17975 => "0000001101011110",
17976 => "0000001101011110",
17977 => "0000001101011110",
17978 => "0000001101011110",
17979 => "0000001101011110",
17980 => "0000001101011111",
17981 => "0000001101011111",
17982 => "0000001101011111",
17983 => "0000001101011111",
17984 => "0000001101011111",
17985 => "0000001101100000",
17986 => "0000001101100000",
17987 => "0000001101100000",
17988 => "0000001101100000",
17989 => "0000001101100000",
17990 => "0000001101100001",
17991 => "0000001101100001",
17992 => "0000001101100001",
17993 => "0000001101100001",
17994 => "0000001101100001",
17995 => "0000001101100010",
17996 => "0000001101100010",
17997 => "0000001101100010",
17998 => "0000001101100010",
17999 => "0000001101100011",
18000 => "0000001101100011",
18001 => "0000001101100011",
18002 => "0000001101100011",
18003 => "0000001101100011",
18004 => "0000001101100100",
18005 => "0000001101100100",
18006 => "0000001101100100",
18007 => "0000001101100100",
18008 => "0000001101100100",
18009 => "0000001101100101",
18010 => "0000001101100101",
18011 => "0000001101100101",
18012 => "0000001101100101",
18013 => "0000001101100101",
18014 => "0000001101100110",
18015 => "0000001101100110",
18016 => "0000001101100110",
18017 => "0000001101100110",
18018 => "0000001101100110",
18019 => "0000001101100111",
18020 => "0000001101100111",
18021 => "0000001101100111",
18022 => "0000001101100111",
18023 => "0000001101100111",
18024 => "0000001101101000",
18025 => "0000001101101000",
18026 => "0000001101101000",
18027 => "0000001101101000",
18028 => "0000001101101000",
18029 => "0000001101101001",
18030 => "0000001101101001",
18031 => "0000001101101001",
18032 => "0000001101101001",
18033 => "0000001101101010",
18034 => "0000001101101010",
18035 => "0000001101101010",
18036 => "0000001101101010",
18037 => "0000001101101010",
18038 => "0000001101101011",
18039 => "0000001101101011",
18040 => "0000001101101011",
18041 => "0000001101101011",
18042 => "0000001101101011",
18043 => "0000001101101100",
18044 => "0000001101101100",
18045 => "0000001101101100",
18046 => "0000001101101100",
18047 => "0000001101101100",
18048 => "0000001101101101",
18049 => "0000001101101101",
18050 => "0000001101101101",
18051 => "0000001101101101",
18052 => "0000001101101101",
18053 => "0000001101101110",
18054 => "0000001101101110",
18055 => "0000001101101110",
18056 => "0000001101101110",
18057 => "0000001101101111",
18058 => "0000001101101111",
18059 => "0000001101101111",
18060 => "0000001101101111",
18061 => "0000001101101111",
18062 => "0000001101110000",
18063 => "0000001101110000",
18064 => "0000001101110000",
18065 => "0000001101110000",
18066 => "0000001101110000",
18067 => "0000001101110001",
18068 => "0000001101110001",
18069 => "0000001101110001",
18070 => "0000001101110001",
18071 => "0000001101110001",
18072 => "0000001101110010",
18073 => "0000001101110010",
18074 => "0000001101110010",
18075 => "0000001101110010",
18076 => "0000001101110011",
18077 => "0000001101110011",
18078 => "0000001101110011",
18079 => "0000001101110011",
18080 => "0000001101110011",
18081 => "0000001101110100",
18082 => "0000001101110100",
18083 => "0000001101110100",
18084 => "0000001101110100",
18085 => "0000001101110100",
18086 => "0000001101110101",
18087 => "0000001101110101",
18088 => "0000001101110101",
18089 => "0000001101110101",
18090 => "0000001101110101",
18091 => "0000001101110110",
18092 => "0000001101110110",
18093 => "0000001101110110",
18094 => "0000001101110110",
18095 => "0000001101110111",
18096 => "0000001101110111",
18097 => "0000001101110111",
18098 => "0000001101110111",
18099 => "0000001101110111",
18100 => "0000001101111000",
18101 => "0000001101111000",
18102 => "0000001101111000",
18103 => "0000001101111000",
18104 => "0000001101111000",
18105 => "0000001101111001",
18106 => "0000001101111001",
18107 => "0000001101111001",
18108 => "0000001101111001",
18109 => "0000001101111001",
18110 => "0000001101111010",
18111 => "0000001101111010",
18112 => "0000001101111010",
18113 => "0000001101111010",
18114 => "0000001101111011",
18115 => "0000001101111011",
18116 => "0000001101111011",
18117 => "0000001101111011",
18118 => "0000001101111011",
18119 => "0000001101111100",
18120 => "0000001101111100",
18121 => "0000001101111100",
18122 => "0000001101111100",
18123 => "0000001101111100",
18124 => "0000001101111101",
18125 => "0000001101111101",
18126 => "0000001101111101",
18127 => "0000001101111101",
18128 => "0000001101111101",
18129 => "0000001101111110",
18130 => "0000001101111110",
18131 => "0000001101111110",
18132 => "0000001101111110",
18133 => "0000001101111111",
18134 => "0000001101111111",
18135 => "0000001101111111",
18136 => "0000001101111111",
18137 => "0000001101111111",
18138 => "0000001110000000",
18139 => "0000001110000000",
18140 => "0000001110000000",
18141 => "0000001110000000",
18142 => "0000001110000000",
18143 => "0000001110000001",
18144 => "0000001110000001",
18145 => "0000001110000001",
18146 => "0000001110000001",
18147 => "0000001110000010",
18148 => "0000001110000010",
18149 => "0000001110000010",
18150 => "0000001110000010",
18151 => "0000001110000010",
18152 => "0000001110000011",
18153 => "0000001110000011",
18154 => "0000001110000011",
18155 => "0000001110000011",
18156 => "0000001110000011",
18157 => "0000001110000100",
18158 => "0000001110000100",
18159 => "0000001110000100",
18160 => "0000001110000100",
18161 => "0000001110000101",
18162 => "0000001110000101",
18163 => "0000001110000101",
18164 => "0000001110000101",
18165 => "0000001110000101",
18166 => "0000001110000110",
18167 => "0000001110000110",
18168 => "0000001110000110",
18169 => "0000001110000110",
18170 => "0000001110000110",
18171 => "0000001110000111",
18172 => "0000001110000111",
18173 => "0000001110000111",
18174 => "0000001110000111",
18175 => "0000001110001000",
18176 => "0000001110001000",
18177 => "0000001110001000",
18178 => "0000001110001000",
18179 => "0000001110001000",
18180 => "0000001110001001",
18181 => "0000001110001001",
18182 => "0000001110001001",
18183 => "0000001110001001",
18184 => "0000001110001001",
18185 => "0000001110001010",
18186 => "0000001110001010",
18187 => "0000001110001010",
18188 => "0000001110001010",
18189 => "0000001110001011",
18190 => "0000001110001011",
18191 => "0000001110001011",
18192 => "0000001110001011",
18193 => "0000001110001011",
18194 => "0000001110001100",
18195 => "0000001110001100",
18196 => "0000001110001100",
18197 => "0000001110001100",
18198 => "0000001110001100",
18199 => "0000001110001101",
18200 => "0000001110001101",
18201 => "0000001110001101",
18202 => "0000001110001101",
18203 => "0000001110001110",
18204 => "0000001110001110",
18205 => "0000001110001110",
18206 => "0000001110001110",
18207 => "0000001110001110",
18208 => "0000001110001111",
18209 => "0000001110001111",
18210 => "0000001110001111",
18211 => "0000001110001111",
18212 => "0000001110001111",
18213 => "0000001110010000",
18214 => "0000001110010000",
18215 => "0000001110010000",
18216 => "0000001110010000",
18217 => "0000001110010001",
18218 => "0000001110010001",
18219 => "0000001110010001",
18220 => "0000001110010001",
18221 => "0000001110010001",
18222 => "0000001110010010",
18223 => "0000001110010010",
18224 => "0000001110010010",
18225 => "0000001110010010",
18226 => "0000001110010011",
18227 => "0000001110010011",
18228 => "0000001110010011",
18229 => "0000001110010011",
18230 => "0000001110010011",
18231 => "0000001110010100",
18232 => "0000001110010100",
18233 => "0000001110010100",
18234 => "0000001110010100",
18235 => "0000001110010100",
18236 => "0000001110010101",
18237 => "0000001110010101",
18238 => "0000001110010101",
18239 => "0000001110010101",
18240 => "0000001110010110",
18241 => "0000001110010110",
18242 => "0000001110010110",
18243 => "0000001110010110",
18244 => "0000001110010110",
18245 => "0000001110010111",
18246 => "0000001110010111",
18247 => "0000001110010111",
18248 => "0000001110010111",
18249 => "0000001110011000",
18250 => "0000001110011000",
18251 => "0000001110011000",
18252 => "0000001110011000",
18253 => "0000001110011000",
18254 => "0000001110011001",
18255 => "0000001110011001",
18256 => "0000001110011001",
18257 => "0000001110011001",
18258 => "0000001110011001",
18259 => "0000001110011010",
18260 => "0000001110011010",
18261 => "0000001110011010",
18262 => "0000001110011010",
18263 => "0000001110011011",
18264 => "0000001110011011",
18265 => "0000001110011011",
18266 => "0000001110011011",
18267 => "0000001110011011",
18268 => "0000001110011100",
18269 => "0000001110011100",
18270 => "0000001110011100",
18271 => "0000001110011100",
18272 => "0000001110011101",
18273 => "0000001110011101",
18274 => "0000001110011101",
18275 => "0000001110011101",
18276 => "0000001110011101",
18277 => "0000001110011110",
18278 => "0000001110011110",
18279 => "0000001110011110",
18280 => "0000001110011110",
18281 => "0000001110011111",
18282 => "0000001110011111",
18283 => "0000001110011111",
18284 => "0000001110011111",
18285 => "0000001110011111",
18286 => "0000001110100000",
18287 => "0000001110100000",
18288 => "0000001110100000",
18289 => "0000001110100000",
18290 => "0000001110100001",
18291 => "0000001110100001",
18292 => "0000001110100001",
18293 => "0000001110100001",
18294 => "0000001110100001",
18295 => "0000001110100010",
18296 => "0000001110100010",
18297 => "0000001110100010",
18298 => "0000001110100010",
18299 => "0000001110100010",
18300 => "0000001110100011",
18301 => "0000001110100011",
18302 => "0000001110100011",
18303 => "0000001110100011",
18304 => "0000001110100100",
18305 => "0000001110100100",
18306 => "0000001110100100",
18307 => "0000001110100100",
18308 => "0000001110100100",
18309 => "0000001110100101",
18310 => "0000001110100101",
18311 => "0000001110100101",
18312 => "0000001110100101",
18313 => "0000001110100110",
18314 => "0000001110100110",
18315 => "0000001110100110",
18316 => "0000001110100110",
18317 => "0000001110100110",
18318 => "0000001110100111",
18319 => "0000001110100111",
18320 => "0000001110100111",
18321 => "0000001110100111",
18322 => "0000001110101000",
18323 => "0000001110101000",
18324 => "0000001110101000",
18325 => "0000001110101000",
18326 => "0000001110101000",
18327 => "0000001110101001",
18328 => "0000001110101001",
18329 => "0000001110101001",
18330 => "0000001110101001",
18331 => "0000001110101010",
18332 => "0000001110101010",
18333 => "0000001110101010",
18334 => "0000001110101010",
18335 => "0000001110101010",
18336 => "0000001110101011",
18337 => "0000001110101011",
18338 => "0000001110101011",
18339 => "0000001110101011",
18340 => "0000001110101100",
18341 => "0000001110101100",
18342 => "0000001110101100",
18343 => "0000001110101100",
18344 => "0000001110101100",
18345 => "0000001110101101",
18346 => "0000001110101101",
18347 => "0000001110101101",
18348 => "0000001110101101",
18349 => "0000001110101110",
18350 => "0000001110101110",
18351 => "0000001110101110",
18352 => "0000001110101110",
18353 => "0000001110101110",
18354 => "0000001110101111",
18355 => "0000001110101111",
18356 => "0000001110101111",
18357 => "0000001110101111",
18358 => "0000001110110000",
18359 => "0000001110110000",
18360 => "0000001110110000",
18361 => "0000001110110000",
18362 => "0000001110110001",
18363 => "0000001110110001",
18364 => "0000001110110001",
18365 => "0000001110110001",
18366 => "0000001110110001",
18367 => "0000001110110010",
18368 => "0000001110110010",
18369 => "0000001110110010",
18370 => "0000001110110010",
18371 => "0000001110110011",
18372 => "0000001110110011",
18373 => "0000001110110011",
18374 => "0000001110110011",
18375 => "0000001110110011",
18376 => "0000001110110100",
18377 => "0000001110110100",
18378 => "0000001110110100",
18379 => "0000001110110100",
18380 => "0000001110110101",
18381 => "0000001110110101",
18382 => "0000001110110101",
18383 => "0000001110110101",
18384 => "0000001110110101",
18385 => "0000001110110110",
18386 => "0000001110110110",
18387 => "0000001110110110",
18388 => "0000001110110110",
18389 => "0000001110110111",
18390 => "0000001110110111",
18391 => "0000001110110111",
18392 => "0000001110110111",
18393 => "0000001110110111",
18394 => "0000001110111000",
18395 => "0000001110111000",
18396 => "0000001110111000",
18397 => "0000001110111000",
18398 => "0000001110111001",
18399 => "0000001110111001",
18400 => "0000001110111001",
18401 => "0000001110111001",
18402 => "0000001110111010",
18403 => "0000001110111010",
18404 => "0000001110111010",
18405 => "0000001110111010",
18406 => "0000001110111010",
18407 => "0000001110111011",
18408 => "0000001110111011",
18409 => "0000001110111011",
18410 => "0000001110111011",
18411 => "0000001110111100",
18412 => "0000001110111100",
18413 => "0000001110111100",
18414 => "0000001110111100",
18415 => "0000001110111100",
18416 => "0000001110111101",
18417 => "0000001110111101",
18418 => "0000001110111101",
18419 => "0000001110111101",
18420 => "0000001110111110",
18421 => "0000001110111110",
18422 => "0000001110111110",
18423 => "0000001110111110",
18424 => "0000001110111110",
18425 => "0000001110111111",
18426 => "0000001110111111",
18427 => "0000001110111111",
18428 => "0000001110111111",
18429 => "0000001111000000",
18430 => "0000001111000000",
18431 => "0000001111000000",
18432 => "0000001111000000",
18433 => "0000001111000001",
18434 => "0000001111000001",
18435 => "0000001111000001",
18436 => "0000001111000001",
18437 => "0000001111000001",
18438 => "0000001111000010",
18439 => "0000001111000010",
18440 => "0000001111000010",
18441 => "0000001111000010",
18442 => "0000001111000011",
18443 => "0000001111000011",
18444 => "0000001111000011",
18445 => "0000001111000011",
18446 => "0000001111000100",
18447 => "0000001111000100",
18448 => "0000001111000100",
18449 => "0000001111000100",
18450 => "0000001111000100",
18451 => "0000001111000101",
18452 => "0000001111000101",
18453 => "0000001111000101",
18454 => "0000001111000101",
18455 => "0000001111000110",
18456 => "0000001111000110",
18457 => "0000001111000110",
18458 => "0000001111000110",
18459 => "0000001111000110",
18460 => "0000001111000111",
18461 => "0000001111000111",
18462 => "0000001111000111",
18463 => "0000001111000111",
18464 => "0000001111001000",
18465 => "0000001111001000",
18466 => "0000001111001000",
18467 => "0000001111001000",
18468 => "0000001111001001",
18469 => "0000001111001001",
18470 => "0000001111001001",
18471 => "0000001111001001",
18472 => "0000001111001001",
18473 => "0000001111001010",
18474 => "0000001111001010",
18475 => "0000001111001010",
18476 => "0000001111001010",
18477 => "0000001111001011",
18478 => "0000001111001011",
18479 => "0000001111001011",
18480 => "0000001111001011",
18481 => "0000001111001100",
18482 => "0000001111001100",
18483 => "0000001111001100",
18484 => "0000001111001100",
18485 => "0000001111001100",
18486 => "0000001111001101",
18487 => "0000001111001101",
18488 => "0000001111001101",
18489 => "0000001111001101",
18490 => "0000001111001110",
18491 => "0000001111001110",
18492 => "0000001111001110",
18493 => "0000001111001110",
18494 => "0000001111001111",
18495 => "0000001111001111",
18496 => "0000001111001111",
18497 => "0000001111001111",
18498 => "0000001111001111",
18499 => "0000001111010000",
18500 => "0000001111010000",
18501 => "0000001111010000",
18502 => "0000001111010000",
18503 => "0000001111010001",
18504 => "0000001111010001",
18505 => "0000001111010001",
18506 => "0000001111010001",
18507 => "0000001111010010",
18508 => "0000001111010010",
18509 => "0000001111010010",
18510 => "0000001111010010",
18511 => "0000001111010010",
18512 => "0000001111010011",
18513 => "0000001111010011",
18514 => "0000001111010011",
18515 => "0000001111010011",
18516 => "0000001111010100",
18517 => "0000001111010100",
18518 => "0000001111010100",
18519 => "0000001111010100",
18520 => "0000001111010101",
18521 => "0000001111010101",
18522 => "0000001111010101",
18523 => "0000001111010101",
18524 => "0000001111010101",
18525 => "0000001111010110",
18526 => "0000001111010110",
18527 => "0000001111010110",
18528 => "0000001111010110",
18529 => "0000001111010111",
18530 => "0000001111010111",
18531 => "0000001111010111",
18532 => "0000001111010111",
18533 => "0000001111011000",
18534 => "0000001111011000",
18535 => "0000001111011000",
18536 => "0000001111011000",
18537 => "0000001111011001",
18538 => "0000001111011001",
18539 => "0000001111011001",
18540 => "0000001111011001",
18541 => "0000001111011001",
18542 => "0000001111011010",
18543 => "0000001111011010",
18544 => "0000001111011010",
18545 => "0000001111011010",
18546 => "0000001111011011",
18547 => "0000001111011011",
18548 => "0000001111011011",
18549 => "0000001111011011",
18550 => "0000001111011100",
18551 => "0000001111011100",
18552 => "0000001111011100",
18553 => "0000001111011100",
18554 => "0000001111011100",
18555 => "0000001111011101",
18556 => "0000001111011101",
18557 => "0000001111011101",
18558 => "0000001111011101",
18559 => "0000001111011110",
18560 => "0000001111011110",
18561 => "0000001111011110",
18562 => "0000001111011110",
18563 => "0000001111011111",
18564 => "0000001111011111",
18565 => "0000001111011111",
18566 => "0000001111011111",
18567 => "0000001111100000",
18568 => "0000001111100000",
18569 => "0000001111100000",
18570 => "0000001111100000",
18571 => "0000001111100000",
18572 => "0000001111100001",
18573 => "0000001111100001",
18574 => "0000001111100001",
18575 => "0000001111100001",
18576 => "0000001111100010",
18577 => "0000001111100010",
18578 => "0000001111100010",
18579 => "0000001111100010",
18580 => "0000001111100011",
18581 => "0000001111100011",
18582 => "0000001111100011",
18583 => "0000001111100011",
18584 => "0000001111100100",
18585 => "0000001111100100",
18586 => "0000001111100100",
18587 => "0000001111100100",
18588 => "0000001111100100",
18589 => "0000001111100101",
18590 => "0000001111100101",
18591 => "0000001111100101",
18592 => "0000001111100101",
18593 => "0000001111100110",
18594 => "0000001111100110",
18595 => "0000001111100110",
18596 => "0000001111100110",
18597 => "0000001111100111",
18598 => "0000001111100111",
18599 => "0000001111100111",
18600 => "0000001111100111",
18601 => "0000001111101000",
18602 => "0000001111101000",
18603 => "0000001111101000",
18604 => "0000001111101000",
18605 => "0000001111101000",
18606 => "0000001111101001",
18607 => "0000001111101001",
18608 => "0000001111101001",
18609 => "0000001111101001",
18610 => "0000001111101010",
18611 => "0000001111101010",
18612 => "0000001111101010",
18613 => "0000001111101010",
18614 => "0000001111101011",
18615 => "0000001111101011",
18616 => "0000001111101011",
18617 => "0000001111101011",
18618 => "0000001111101100",
18619 => "0000001111101100",
18620 => "0000001111101100",
18621 => "0000001111101100",
18622 => "0000001111101101",
18623 => "0000001111101101",
18624 => "0000001111101101",
18625 => "0000001111101101",
18626 => "0000001111101101",
18627 => "0000001111101110",
18628 => "0000001111101110",
18629 => "0000001111101110",
18630 => "0000001111101110",
18631 => "0000001111101111",
18632 => "0000001111101111",
18633 => "0000001111101111",
18634 => "0000001111101111",
18635 => "0000001111110000",
18636 => "0000001111110000",
18637 => "0000001111110000",
18638 => "0000001111110000",
18639 => "0000001111110001",
18640 => "0000001111110001",
18641 => "0000001111110001",
18642 => "0000001111110001",
18643 => "0000001111110010",
18644 => "0000001111110010",
18645 => "0000001111110010",
18646 => "0000001111110010",
18647 => "0000001111110010",
18648 => "0000001111110011",
18649 => "0000001111110011",
18650 => "0000001111110011",
18651 => "0000001111110011",
18652 => "0000001111110100",
18653 => "0000001111110100",
18654 => "0000001111110100",
18655 => "0000001111110100",
18656 => "0000001111110101",
18657 => "0000001111110101",
18658 => "0000001111110101",
18659 => "0000001111110101",
18660 => "0000001111110110",
18661 => "0000001111110110",
18662 => "0000001111110110",
18663 => "0000001111110110",
18664 => "0000001111110111",
18665 => "0000001111110111",
18666 => "0000001111110111",
18667 => "0000001111110111",
18668 => "0000001111111000",
18669 => "0000001111111000",
18670 => "0000001111111000",
18671 => "0000001111111000",
18672 => "0000001111111000",
18673 => "0000001111111001",
18674 => "0000001111111001",
18675 => "0000001111111001",
18676 => "0000001111111001",
18677 => "0000001111111010",
18678 => "0000001111111010",
18679 => "0000001111111010",
18680 => "0000001111111010",
18681 => "0000001111111011",
18682 => "0000001111111011",
18683 => "0000001111111011",
18684 => "0000001111111011",
18685 => "0000001111111100",
18686 => "0000001111111100",
18687 => "0000001111111100",
18688 => "0000001111111100",
18689 => "0000001111111101",
18690 => "0000001111111101",
18691 => "0000001111111101",
18692 => "0000001111111101",
18693 => "0000001111111110",
18694 => "0000001111111110",
18695 => "0000001111111110",
18696 => "0000001111111110",
18697 => "0000001111111111",
18698 => "0000001111111111",
18699 => "0000001111111111",
18700 => "0000001111111111",
18701 => "0000001111111111",
18702 => "0000010000000000",
18703 => "0000010000000000",
18704 => "0000010000000000",
18705 => "0000010000000001",
18706 => "0000010000000001",
18707 => "0000010000000001",
18708 => "0000010000000001",
18709 => "0000010000000010",
18710 => "0000010000000010",
18711 => "0000010000000010",
18712 => "0000010000000010",
18713 => "0000010000000011",
18714 => "0000010000000011",
18715 => "0000010000000011",
18716 => "0000010000000011",
18717 => "0000010000000100",
18718 => "0000010000000100",
18719 => "0000010000000100",
18720 => "0000010000000100",
18721 => "0000010000000101",
18722 => "0000010000000101",
18723 => "0000010000000101",
18724 => "0000010000000101",
18725 => "0000010000000110",
18726 => "0000010000000110",
18727 => "0000010000000110",
18728 => "0000010000000110",
18729 => "0000010000000111",
18730 => "0000010000000111",
18731 => "0000010000000111",
18732 => "0000010000000111",
18733 => "0000010000001000",
18734 => "0000010000001000",
18735 => "0000010000001000",
18736 => "0000010000001000",
18737 => "0000010000001000",
18738 => "0000010000001001",
18739 => "0000010000001001",
18740 => "0000010000001001",
18741 => "0000010000001001",
18742 => "0000010000001010",
18743 => "0000010000001010",
18744 => "0000010000001010",
18745 => "0000010000001010",
18746 => "0000010000001011",
18747 => "0000010000001011",
18748 => "0000010000001011",
18749 => "0000010000001011",
18750 => "0000010000001100",
18751 => "0000010000001100",
18752 => "0000010000001100",
18753 => "0000010000001100",
18754 => "0000010000001101",
18755 => "0000010000001101",
18756 => "0000010000001101",
18757 => "0000010000001101",
18758 => "0000010000001110",
18759 => "0000010000001110",
18760 => "0000010000001110",
18761 => "0000010000001110",
18762 => "0000010000001111",
18763 => "0000010000001111",
18764 => "0000010000001111",
18765 => "0000010000001111",
18766 => "0000010000010000",
18767 => "0000010000010000",
18768 => "0000010000010000",
18769 => "0000010000010000",
18770 => "0000010000010001",
18771 => "0000010000010001",
18772 => "0000010000010001",
18773 => "0000010000010001",
18774 => "0000010000010010",
18775 => "0000010000010010",
18776 => "0000010000010010",
18777 => "0000010000010010",
18778 => "0000010000010011",
18779 => "0000010000010011",
18780 => "0000010000010011",
18781 => "0000010000010011",
18782 => "0000010000010100",
18783 => "0000010000010100",
18784 => "0000010000010100",
18785 => "0000010000010100",
18786 => "0000010000010101",
18787 => "0000010000010101",
18788 => "0000010000010101",
18789 => "0000010000010101",
18790 => "0000010000010110",
18791 => "0000010000010110",
18792 => "0000010000010110",
18793 => "0000010000010110",
18794 => "0000010000010110",
18795 => "0000010000010111",
18796 => "0000010000010111",
18797 => "0000010000010111",
18798 => "0000010000010111",
18799 => "0000010000011000",
18800 => "0000010000011000",
18801 => "0000010000011000",
18802 => "0000010000011000",
18803 => "0000010000011001",
18804 => "0000010000011001",
18805 => "0000010000011001",
18806 => "0000010000011001",
18807 => "0000010000011010",
18808 => "0000010000011010",
18809 => "0000010000011010",
18810 => "0000010000011010",
18811 => "0000010000011011",
18812 => "0000010000011011",
18813 => "0000010000011011",
18814 => "0000010000011011",
18815 => "0000010000011100",
18816 => "0000010000011100",
18817 => "0000010000011100",
18818 => "0000010000011100",
18819 => "0000010000011101",
18820 => "0000010000011101",
18821 => "0000010000011101",
18822 => "0000010000011101",
18823 => "0000010000011110",
18824 => "0000010000011110",
18825 => "0000010000011110",
18826 => "0000010000011110",
18827 => "0000010000011111",
18828 => "0000010000011111",
18829 => "0000010000011111",
18830 => "0000010000011111",
18831 => "0000010000100000",
18832 => "0000010000100000",
18833 => "0000010000100000",
18834 => "0000010000100000",
18835 => "0000010000100001",
18836 => "0000010000100001",
18837 => "0000010000100001",
18838 => "0000010000100001",
18839 => "0000010000100010",
18840 => "0000010000100010",
18841 => "0000010000100010",
18842 => "0000010000100010",
18843 => "0000010000100011",
18844 => "0000010000100011",
18845 => "0000010000100011",
18846 => "0000010000100011",
18847 => "0000010000100100",
18848 => "0000010000100100",
18849 => "0000010000100100",
18850 => "0000010000100100",
18851 => "0000010000100101",
18852 => "0000010000100101",
18853 => "0000010000100101",
18854 => "0000010000100101",
18855 => "0000010000100110",
18856 => "0000010000100110",
18857 => "0000010000100110",
18858 => "0000010000100110",
18859 => "0000010000100111",
18860 => "0000010000100111",
18861 => "0000010000100111",
18862 => "0000010000100111",
18863 => "0000010000101000",
18864 => "0000010000101000",
18865 => "0000010000101000",
18866 => "0000010000101000",
18867 => "0000010000101001",
18868 => "0000010000101001",
18869 => "0000010000101001",
18870 => "0000010000101001",
18871 => "0000010000101010",
18872 => "0000010000101010",
18873 => "0000010000101010",
18874 => "0000010000101010",
18875 => "0000010000101011",
18876 => "0000010000101011",
18877 => "0000010000101011",
18878 => "0000010000101011",
18879 => "0000010000101100",
18880 => "0000010000101100",
18881 => "0000010000101100",
18882 => "0000010000101100",
18883 => "0000010000101101",
18884 => "0000010000101101",
18885 => "0000010000101101",
18886 => "0000010000101101",
18887 => "0000010000101110",
18888 => "0000010000101110",
18889 => "0000010000101110",
18890 => "0000010000101110",
18891 => "0000010000101111",
18892 => "0000010000101111",
18893 => "0000010000101111",
18894 => "0000010000110000",
18895 => "0000010000110000",
18896 => "0000010000110000",
18897 => "0000010000110000",
18898 => "0000010000110001",
18899 => "0000010000110001",
18900 => "0000010000110001",
18901 => "0000010000110001",
18902 => "0000010000110010",
18903 => "0000010000110010",
18904 => "0000010000110010",
18905 => "0000010000110010",
18906 => "0000010000110011",
18907 => "0000010000110011",
18908 => "0000010000110011",
18909 => "0000010000110011",
18910 => "0000010000110100",
18911 => "0000010000110100",
18912 => "0000010000110100",
18913 => "0000010000110100",
18914 => "0000010000110101",
18915 => "0000010000110101",
18916 => "0000010000110101",
18917 => "0000010000110101",
18918 => "0000010000110110",
18919 => "0000010000110110",
18920 => "0000010000110110",
18921 => "0000010000110110",
18922 => "0000010000110111",
18923 => "0000010000110111",
18924 => "0000010000110111",
18925 => "0000010000110111",
18926 => "0000010000111000",
18927 => "0000010000111000",
18928 => "0000010000111000",
18929 => "0000010000111000",
18930 => "0000010000111001",
18931 => "0000010000111001",
18932 => "0000010000111001",
18933 => "0000010000111001",
18934 => "0000010000111010",
18935 => "0000010000111010",
18936 => "0000010000111010",
18937 => "0000010000111010",
18938 => "0000010000111011",
18939 => "0000010000111011",
18940 => "0000010000111011",
18941 => "0000010000111011",
18942 => "0000010000111100",
18943 => "0000010000111100",
18944 => "0000010000111100",
18945 => "0000010000111100",
18946 => "0000010000111101",
18947 => "0000010000111101",
18948 => "0000010000111101",
18949 => "0000010000111110",
18950 => "0000010000111110",
18951 => "0000010000111110",
18952 => "0000010000111110",
18953 => "0000010000111111",
18954 => "0000010000111111",
18955 => "0000010000111111",
18956 => "0000010000111111",
18957 => "0000010001000000",
18958 => "0000010001000000",
18959 => "0000010001000000",
18960 => "0000010001000000",
18961 => "0000010001000001",
18962 => "0000010001000001",
18963 => "0000010001000001",
18964 => "0000010001000001",
18965 => "0000010001000010",
18966 => "0000010001000010",
18967 => "0000010001000010",
18968 => "0000010001000010",
18969 => "0000010001000011",
18970 => "0000010001000011",
18971 => "0000010001000011",
18972 => "0000010001000011",
18973 => "0000010001000100",
18974 => "0000010001000100",
18975 => "0000010001000100",
18976 => "0000010001000100",
18977 => "0000010001000101",
18978 => "0000010001000101",
18979 => "0000010001000101",
18980 => "0000010001000101",
18981 => "0000010001000110",
18982 => "0000010001000110",
18983 => "0000010001000110",
18984 => "0000010001000111",
18985 => "0000010001000111",
18986 => "0000010001000111",
18987 => "0000010001000111",
18988 => "0000010001001000",
18989 => "0000010001001000",
18990 => "0000010001001000",
18991 => "0000010001001000",
18992 => "0000010001001001",
18993 => "0000010001001001",
18994 => "0000010001001001",
18995 => "0000010001001001",
18996 => "0000010001001010",
18997 => "0000010001001010",
18998 => "0000010001001010",
18999 => "0000010001001010",
19000 => "0000010001001011",
19001 => "0000010001001011",
19002 => "0000010001001011",
19003 => "0000010001001011",
19004 => "0000010001001100",
19005 => "0000010001001100",
19006 => "0000010001001100",
19007 => "0000010001001100",
19008 => "0000010001001101",
19009 => "0000010001001101",
19010 => "0000010001001101",
19011 => "0000010001001110",
19012 => "0000010001001110",
19013 => "0000010001001110",
19014 => "0000010001001110",
19015 => "0000010001001111",
19016 => "0000010001001111",
19017 => "0000010001001111",
19018 => "0000010001001111",
19019 => "0000010001010000",
19020 => "0000010001010000",
19021 => "0000010001010000",
19022 => "0000010001010000",
19023 => "0000010001010001",
19024 => "0000010001010001",
19025 => "0000010001010001",
19026 => "0000010001010001",
19027 => "0000010001010010",
19028 => "0000010001010010",
19029 => "0000010001010010",
19030 => "0000010001010010",
19031 => "0000010001010011",
19032 => "0000010001010011",
19033 => "0000010001010011",
19034 => "0000010001010100",
19035 => "0000010001010100",
19036 => "0000010001010100",
19037 => "0000010001010100",
19038 => "0000010001010101",
19039 => "0000010001010101",
19040 => "0000010001010101",
19041 => "0000010001010101",
19042 => "0000010001010110",
19043 => "0000010001010110",
19044 => "0000010001010110",
19045 => "0000010001010110",
19046 => "0000010001010111",
19047 => "0000010001010111",
19048 => "0000010001010111",
19049 => "0000010001010111",
19050 => "0000010001011000",
19051 => "0000010001011000",
19052 => "0000010001011000",
19053 => "0000010001011000",
19054 => "0000010001011001",
19055 => "0000010001011001",
19056 => "0000010001011001",
19057 => "0000010001011010",
19058 => "0000010001011010",
19059 => "0000010001011010",
19060 => "0000010001011010",
19061 => "0000010001011011",
19062 => "0000010001011011",
19063 => "0000010001011011",
19064 => "0000010001011011",
19065 => "0000010001011100",
19066 => "0000010001011100",
19067 => "0000010001011100",
19068 => "0000010001011100",
19069 => "0000010001011101",
19070 => "0000010001011101",
19071 => "0000010001011101",
19072 => "0000010001011101",
19073 => "0000010001011110",
19074 => "0000010001011110",
19075 => "0000010001011110",
19076 => "0000010001011111",
19077 => "0000010001011111",
19078 => "0000010001011111",
19079 => "0000010001011111",
19080 => "0000010001100000",
19081 => "0000010001100000",
19082 => "0000010001100000",
19083 => "0000010001100000",
19084 => "0000010001100001",
19085 => "0000010001100001",
19086 => "0000010001100001",
19087 => "0000010001100001",
19088 => "0000010001100010",
19089 => "0000010001100010",
19090 => "0000010001100010",
19091 => "0000010001100010",
19092 => "0000010001100011",
19093 => "0000010001100011",
19094 => "0000010001100011",
19095 => "0000010001100100",
19096 => "0000010001100100",
19097 => "0000010001100100",
19098 => "0000010001100100",
19099 => "0000010001100101",
19100 => "0000010001100101",
19101 => "0000010001100101",
19102 => "0000010001100101",
19103 => "0000010001100110",
19104 => "0000010001100110",
19105 => "0000010001100110",
19106 => "0000010001100110",
19107 => "0000010001100111",
19108 => "0000010001100111",
19109 => "0000010001100111",
19110 => "0000010001101000",
19111 => "0000010001101000",
19112 => "0000010001101000",
19113 => "0000010001101000",
19114 => "0000010001101001",
19115 => "0000010001101001",
19116 => "0000010001101001",
19117 => "0000010001101001",
19118 => "0000010001101010",
19119 => "0000010001101010",
19120 => "0000010001101010",
19121 => "0000010001101010",
19122 => "0000010001101011",
19123 => "0000010001101011",
19124 => "0000010001101011",
19125 => "0000010001101100",
19126 => "0000010001101100",
19127 => "0000010001101100",
19128 => "0000010001101100",
19129 => "0000010001101101",
19130 => "0000010001101101",
19131 => "0000010001101101",
19132 => "0000010001101101",
19133 => "0000010001101110",
19134 => "0000010001101110",
19135 => "0000010001101110",
19136 => "0000010001101110",
19137 => "0000010001101111",
19138 => "0000010001101111",
19139 => "0000010001101111",
19140 => "0000010001110000",
19141 => "0000010001110000",
19142 => "0000010001110000",
19143 => "0000010001110000",
19144 => "0000010001110001",
19145 => "0000010001110001",
19146 => "0000010001110001",
19147 => "0000010001110001",
19148 => "0000010001110010",
19149 => "0000010001110010",
19150 => "0000010001110010",
19151 => "0000010001110010",
19152 => "0000010001110011",
19153 => "0000010001110011",
19154 => "0000010001110011",
19155 => "0000010001110100",
19156 => "0000010001110100",
19157 => "0000010001110100",
19158 => "0000010001110100",
19159 => "0000010001110101",
19160 => "0000010001110101",
19161 => "0000010001110101",
19162 => "0000010001110101",
19163 => "0000010001110110",
19164 => "0000010001110110",
19165 => "0000010001110110",
19166 => "0000010001110111",
19167 => "0000010001110111",
19168 => "0000010001110111",
19169 => "0000010001110111",
19170 => "0000010001111000",
19171 => "0000010001111000",
19172 => "0000010001111000",
19173 => "0000010001111000",
19174 => "0000010001111001",
19175 => "0000010001111001",
19176 => "0000010001111001",
19177 => "0000010001111001",
19178 => "0000010001111010",
19179 => "0000010001111010",
19180 => "0000010001111010",
19181 => "0000010001111011",
19182 => "0000010001111011",
19183 => "0000010001111011",
19184 => "0000010001111011",
19185 => "0000010001111100",
19186 => "0000010001111100",
19187 => "0000010001111100",
19188 => "0000010001111100",
19189 => "0000010001111101",
19190 => "0000010001111101",
19191 => "0000010001111101",
19192 => "0000010001111110",
19193 => "0000010001111110",
19194 => "0000010001111110",
19195 => "0000010001111110",
19196 => "0000010001111111",
19197 => "0000010001111111",
19198 => "0000010001111111",
19199 => "0000010001111111",
19200 => "0000010010000000",
19201 => "0000010010000000",
19202 => "0000010010000000",
19203 => "0000010010000001",
19204 => "0000010010000001",
19205 => "0000010010000001",
19206 => "0000010010000001",
19207 => "0000010010000010",
19208 => "0000010010000010",
19209 => "0000010010000010",
19210 => "0000010010000010",
19211 => "0000010010000011",
19212 => "0000010010000011",
19213 => "0000010010000011",
19214 => "0000010010000100",
19215 => "0000010010000100",
19216 => "0000010010000100",
19217 => "0000010010000100",
19218 => "0000010010000101",
19219 => "0000010010000101",
19220 => "0000010010000101",
19221 => "0000010010000101",
19222 => "0000010010000110",
19223 => "0000010010000110",
19224 => "0000010010000110",
19225 => "0000010010000111",
19226 => "0000010010000111",
19227 => "0000010010000111",
19228 => "0000010010000111",
19229 => "0000010010001000",
19230 => "0000010010001000",
19231 => "0000010010001000",
19232 => "0000010010001000",
19233 => "0000010010001001",
19234 => "0000010010001001",
19235 => "0000010010001001",
19236 => "0000010010001010",
19237 => "0000010010001010",
19238 => "0000010010001010",
19239 => "0000010010001010",
19240 => "0000010010001011",
19241 => "0000010010001011",
19242 => "0000010010001011",
19243 => "0000010010001011",
19244 => "0000010010001100",
19245 => "0000010010001100",
19246 => "0000010010001100",
19247 => "0000010010001101",
19248 => "0000010010001101",
19249 => "0000010010001101",
19250 => "0000010010001101",
19251 => "0000010010001110",
19252 => "0000010010001110",
19253 => "0000010010001110",
19254 => "0000010010001110",
19255 => "0000010010001111",
19256 => "0000010010001111",
19257 => "0000010010001111",
19258 => "0000010010010000",
19259 => "0000010010010000",
19260 => "0000010010010000",
19261 => "0000010010010000",
19262 => "0000010010010001",
19263 => "0000010010010001",
19264 => "0000010010010001",
19265 => "0000010010010001",
19266 => "0000010010010010",
19267 => "0000010010010010",
19268 => "0000010010010010",
19269 => "0000010010010011",
19270 => "0000010010010011",
19271 => "0000010010010011",
19272 => "0000010010010011",
19273 => "0000010010010100",
19274 => "0000010010010100",
19275 => "0000010010010100",
19276 => "0000010010010101",
19277 => "0000010010010101",
19278 => "0000010010010101",
19279 => "0000010010010101",
19280 => "0000010010010110",
19281 => "0000010010010110",
19282 => "0000010010010110",
19283 => "0000010010010110",
19284 => "0000010010010111",
19285 => "0000010010010111",
19286 => "0000010010010111",
19287 => "0000010010011000",
19288 => "0000010010011000",
19289 => "0000010010011000",
19290 => "0000010010011000",
19291 => "0000010010011001",
19292 => "0000010010011001",
19293 => "0000010010011001",
19294 => "0000010010011001",
19295 => "0000010010011010",
19296 => "0000010010011010",
19297 => "0000010010011010",
19298 => "0000010010011011",
19299 => "0000010010011011",
19300 => "0000010010011011",
19301 => "0000010010011011",
19302 => "0000010010011100",
19303 => "0000010010011100",
19304 => "0000010010011100",
19305 => "0000010010011101",
19306 => "0000010010011101",
19307 => "0000010010011101",
19308 => "0000010010011101",
19309 => "0000010010011110",
19310 => "0000010010011110",
19311 => "0000010010011110",
19312 => "0000010010011110",
19313 => "0000010010011111",
19314 => "0000010010011111",
19315 => "0000010010011111",
19316 => "0000010010100000",
19317 => "0000010010100000",
19318 => "0000010010100000",
19319 => "0000010010100000",
19320 => "0000010010100001",
19321 => "0000010010100001",
19322 => "0000010010100001",
19323 => "0000010010100010",
19324 => "0000010010100010",
19325 => "0000010010100010",
19326 => "0000010010100010",
19327 => "0000010010100011",
19328 => "0000010010100011",
19329 => "0000010010100011",
19330 => "0000010010100011",
19331 => "0000010010100100",
19332 => "0000010010100100",
19333 => "0000010010100100",
19334 => "0000010010100101",
19335 => "0000010010100101",
19336 => "0000010010100101",
19337 => "0000010010100101",
19338 => "0000010010100110",
19339 => "0000010010100110",
19340 => "0000010010100110",
19341 => "0000010010100111",
19342 => "0000010010100111",
19343 => "0000010010100111",
19344 => "0000010010100111",
19345 => "0000010010101000",
19346 => "0000010010101000",
19347 => "0000010010101000",
19348 => "0000010010101001",
19349 => "0000010010101001",
19350 => "0000010010101001",
19351 => "0000010010101001",
19352 => "0000010010101010",
19353 => "0000010010101010",
19354 => "0000010010101010",
19355 => "0000010010101011",
19356 => "0000010010101011",
19357 => "0000010010101011",
19358 => "0000010010101011",
19359 => "0000010010101100",
19360 => "0000010010101100",
19361 => "0000010010101100",
19362 => "0000010010101100",
19363 => "0000010010101101",
19364 => "0000010010101101",
19365 => "0000010010101101",
19366 => "0000010010101110",
19367 => "0000010010101110",
19368 => "0000010010101110",
19369 => "0000010010101110",
19370 => "0000010010101111",
19371 => "0000010010101111",
19372 => "0000010010101111",
19373 => "0000010010110000",
19374 => "0000010010110000",
19375 => "0000010010110000",
19376 => "0000010010110000",
19377 => "0000010010110001",
19378 => "0000010010110001",
19379 => "0000010010110001",
19380 => "0000010010110010",
19381 => "0000010010110010",
19382 => "0000010010110010",
19383 => "0000010010110010",
19384 => "0000010010110011",
19385 => "0000010010110011",
19386 => "0000010010110011",
19387 => "0000010010110100",
19388 => "0000010010110100",
19389 => "0000010010110100",
19390 => "0000010010110100",
19391 => "0000010010110101",
19392 => "0000010010110101",
19393 => "0000010010110101",
19394 => "0000010010110110",
19395 => "0000010010110110",
19396 => "0000010010110110",
19397 => "0000010010110110",
19398 => "0000010010110111",
19399 => "0000010010110111",
19400 => "0000010010110111",
19401 => "0000010010110111",
19402 => "0000010010111000",
19403 => "0000010010111000",
19404 => "0000010010111000",
19405 => "0000010010111001",
19406 => "0000010010111001",
19407 => "0000010010111001",
19408 => "0000010010111001",
19409 => "0000010010111010",
19410 => "0000010010111010",
19411 => "0000010010111010",
19412 => "0000010010111011",
19413 => "0000010010111011",
19414 => "0000010010111011",
19415 => "0000010010111011",
19416 => "0000010010111100",
19417 => "0000010010111100",
19418 => "0000010010111100",
19419 => "0000010010111101",
19420 => "0000010010111101",
19421 => "0000010010111101",
19422 => "0000010010111101",
19423 => "0000010010111110",
19424 => "0000010010111110",
19425 => "0000010010111110",
19426 => "0000010010111111",
19427 => "0000010010111111",
19428 => "0000010010111111",
19429 => "0000010010111111",
19430 => "0000010011000000",
19431 => "0000010011000000",
19432 => "0000010011000000",
19433 => "0000010011000001",
19434 => "0000010011000001",
19435 => "0000010011000001",
19436 => "0000010011000001",
19437 => "0000010011000010",
19438 => "0000010011000010",
19439 => "0000010011000010",
19440 => "0000010011000011",
19441 => "0000010011000011",
19442 => "0000010011000011",
19443 => "0000010011000011",
19444 => "0000010011000100",
19445 => "0000010011000100",
19446 => "0000010011000100",
19447 => "0000010011000101",
19448 => "0000010011000101",
19449 => "0000010011000101",
19450 => "0000010011000101",
19451 => "0000010011000110",
19452 => "0000010011000110",
19453 => "0000010011000110",
19454 => "0000010011000111",
19455 => "0000010011000111",
19456 => "0000010011000111",
19457 => "0000010011001000",
19458 => "0000010011001000",
19459 => "0000010011001000",
19460 => "0000010011001000",
19461 => "0000010011001001",
19462 => "0000010011001001",
19463 => "0000010011001001",
19464 => "0000010011001010",
19465 => "0000010011001010",
19466 => "0000010011001010",
19467 => "0000010011001010",
19468 => "0000010011001011",
19469 => "0000010011001011",
19470 => "0000010011001011",
19471 => "0000010011001100",
19472 => "0000010011001100",
19473 => "0000010011001100",
19474 => "0000010011001100",
19475 => "0000010011001101",
19476 => "0000010011001101",
19477 => "0000010011001101",
19478 => "0000010011001110",
19479 => "0000010011001110",
19480 => "0000010011001110",
19481 => "0000010011001110",
19482 => "0000010011001111",
19483 => "0000010011001111",
19484 => "0000010011001111",
19485 => "0000010011010000",
19486 => "0000010011010000",
19487 => "0000010011010000",
19488 => "0000010011010000",
19489 => "0000010011010001",
19490 => "0000010011010001",
19491 => "0000010011010001",
19492 => "0000010011010010",
19493 => "0000010011010010",
19494 => "0000010011010010",
19495 => "0000010011010010",
19496 => "0000010011010011",
19497 => "0000010011010011",
19498 => "0000010011010011",
19499 => "0000010011010100",
19500 => "0000010011010100",
19501 => "0000010011010100",
19502 => "0000010011010101",
19503 => "0000010011010101",
19504 => "0000010011010101",
19505 => "0000010011010101",
19506 => "0000010011010110",
19507 => "0000010011010110",
19508 => "0000010011010110",
19509 => "0000010011010111",
19510 => "0000010011010111",
19511 => "0000010011010111",
19512 => "0000010011010111",
19513 => "0000010011011000",
19514 => "0000010011011000",
19515 => "0000010011011000",
19516 => "0000010011011001",
19517 => "0000010011011001",
19518 => "0000010011011001",
19519 => "0000010011011001",
19520 => "0000010011011010",
19521 => "0000010011011010",
19522 => "0000010011011010",
19523 => "0000010011011011",
19524 => "0000010011011011",
19525 => "0000010011011011",
19526 => "0000010011011011",
19527 => "0000010011011100",
19528 => "0000010011011100",
19529 => "0000010011011100",
19530 => "0000010011011101",
19531 => "0000010011011101",
19532 => "0000010011011101",
19533 => "0000010011011110",
19534 => "0000010011011110",
19535 => "0000010011011110",
19536 => "0000010011011110",
19537 => "0000010011011111",
19538 => "0000010011011111",
19539 => "0000010011011111",
19540 => "0000010011100000",
19541 => "0000010011100000",
19542 => "0000010011100000",
19543 => "0000010011100000",
19544 => "0000010011100001",
19545 => "0000010011100001",
19546 => "0000010011100001",
19547 => "0000010011100010",
19548 => "0000010011100010",
19549 => "0000010011100010",
19550 => "0000010011100011",
19551 => "0000010011100011",
19552 => "0000010011100011",
19553 => "0000010011100011",
19554 => "0000010011100100",
19555 => "0000010011100100",
19556 => "0000010011100100",
19557 => "0000010011100101",
19558 => "0000010011100101",
19559 => "0000010011100101",
19560 => "0000010011100101",
19561 => "0000010011100110",
19562 => "0000010011100110",
19563 => "0000010011100110",
19564 => "0000010011100111",
19565 => "0000010011100111",
19566 => "0000010011100111",
19567 => "0000010011101000",
19568 => "0000010011101000",
19569 => "0000010011101000",
19570 => "0000010011101000",
19571 => "0000010011101001",
19572 => "0000010011101001",
19573 => "0000010011101001",
19574 => "0000010011101010",
19575 => "0000010011101010",
19576 => "0000010011101010",
19577 => "0000010011101010",
19578 => "0000010011101011",
19579 => "0000010011101011",
19580 => "0000010011101011",
19581 => "0000010011101100",
19582 => "0000010011101100",
19583 => "0000010011101100",
19584 => "0000010011101101",
19585 => "0000010011101101",
19586 => "0000010011101101",
19587 => "0000010011101101",
19588 => "0000010011101110",
19589 => "0000010011101110",
19590 => "0000010011101110",
19591 => "0000010011101111",
19592 => "0000010011101111",
19593 => "0000010011101111",
19594 => "0000010011110000",
19595 => "0000010011110000",
19596 => "0000010011110000",
19597 => "0000010011110000",
19598 => "0000010011110001",
19599 => "0000010011110001",
19600 => "0000010011110001",
19601 => "0000010011110010",
19602 => "0000010011110010",
19603 => "0000010011110010",
19604 => "0000010011110010",
19605 => "0000010011110011",
19606 => "0000010011110011",
19607 => "0000010011110011",
19608 => "0000010011110100",
19609 => "0000010011110100",
19610 => "0000010011110100",
19611 => "0000010011110101",
19612 => "0000010011110101",
19613 => "0000010011110101",
19614 => "0000010011110101",
19615 => "0000010011110110",
19616 => "0000010011110110",
19617 => "0000010011110110",
19618 => "0000010011110111",
19619 => "0000010011110111",
19620 => "0000010011110111",
19621 => "0000010011111000",
19622 => "0000010011111000",
19623 => "0000010011111000",
19624 => "0000010011111000",
19625 => "0000010011111001",
19626 => "0000010011111001",
19627 => "0000010011111001",
19628 => "0000010011111010",
19629 => "0000010011111010",
19630 => "0000010011111010",
19631 => "0000010011111011",
19632 => "0000010011111011",
19633 => "0000010011111011",
19634 => "0000010011111011",
19635 => "0000010011111100",
19636 => "0000010011111100",
19637 => "0000010011111100",
19638 => "0000010011111101",
19639 => "0000010011111101",
19640 => "0000010011111101",
19641 => "0000010011111110",
19642 => "0000010011111110",
19643 => "0000010011111110",
19644 => "0000010011111110",
19645 => "0000010011111111",
19646 => "0000010011111111",
19647 => "0000010011111111",
19648 => "0000010100000000",
19649 => "0000010100000000",
19650 => "0000010100000000",
19651 => "0000010100000001",
19652 => "0000010100000001",
19653 => "0000010100000001",
19654 => "0000010100000001",
19655 => "0000010100000010",
19656 => "0000010100000010",
19657 => "0000010100000010",
19658 => "0000010100000011",
19659 => "0000010100000011",
19660 => "0000010100000011",
19661 => "0000010100000100",
19662 => "0000010100000100",
19663 => "0000010100000100",
19664 => "0000010100000100",
19665 => "0000010100000101",
19666 => "0000010100000101",
19667 => "0000010100000101",
19668 => "0000010100000110",
19669 => "0000010100000110",
19670 => "0000010100000110",
19671 => "0000010100000111",
19672 => "0000010100000111",
19673 => "0000010100000111",
19674 => "0000010100000111",
19675 => "0000010100001000",
19676 => "0000010100001000",
19677 => "0000010100001000",
19678 => "0000010100001001",
19679 => "0000010100001001",
19680 => "0000010100001001",
19681 => "0000010100001010",
19682 => "0000010100001010",
19683 => "0000010100001010",
19684 => "0000010100001010",
19685 => "0000010100001011",
19686 => "0000010100001011",
19687 => "0000010100001011",
19688 => "0000010100001100",
19689 => "0000010100001100",
19690 => "0000010100001100",
19691 => "0000010100001101",
19692 => "0000010100001101",
19693 => "0000010100001101",
19694 => "0000010100001110",
19695 => "0000010100001110",
19696 => "0000010100001110",
19697 => "0000010100001110",
19698 => "0000010100001111",
19699 => "0000010100001111",
19700 => "0000010100001111",
19701 => "0000010100010000",
19702 => "0000010100010000",
19703 => "0000010100010000",
19704 => "0000010100010001",
19705 => "0000010100010001",
19706 => "0000010100010001",
19707 => "0000010100010001",
19708 => "0000010100010010",
19709 => "0000010100010010",
19710 => "0000010100010010",
19711 => "0000010100010011",
19712 => "0000010100010011",
19713 => "0000010100010011",
19714 => "0000010100010100",
19715 => "0000010100010100",
19716 => "0000010100010100",
19717 => "0000010100010101",
19718 => "0000010100010101",
19719 => "0000010100010101",
19720 => "0000010100010101",
19721 => "0000010100010110",
19722 => "0000010100010110",
19723 => "0000010100010110",
19724 => "0000010100010111",
19725 => "0000010100010111",
19726 => "0000010100010111",
19727 => "0000010100011000",
19728 => "0000010100011000",
19729 => "0000010100011000",
19730 => "0000010100011000",
19731 => "0000010100011001",
19732 => "0000010100011001",
19733 => "0000010100011001",
19734 => "0000010100011010",
19735 => "0000010100011010",
19736 => "0000010100011010",
19737 => "0000010100011011",
19738 => "0000010100011011",
19739 => "0000010100011011",
19740 => "0000010100011100",
19741 => "0000010100011100",
19742 => "0000010100011100",
19743 => "0000010100011100",
19744 => "0000010100011101",
19745 => "0000010100011101",
19746 => "0000010100011101",
19747 => "0000010100011110",
19748 => "0000010100011110",
19749 => "0000010100011110",
19750 => "0000010100011111",
19751 => "0000010100011111",
19752 => "0000010100011111",
19753 => "0000010100100000",
19754 => "0000010100100000",
19755 => "0000010100100000",
19756 => "0000010100100000",
19757 => "0000010100100001",
19758 => "0000010100100001",
19759 => "0000010100100001",
19760 => "0000010100100010",
19761 => "0000010100100010",
19762 => "0000010100100010",
19763 => "0000010100100011",
19764 => "0000010100100011",
19765 => "0000010100100011",
19766 => "0000010100100100",
19767 => "0000010100100100",
19768 => "0000010100100100",
19769 => "0000010100100100",
19770 => "0000010100100101",
19771 => "0000010100100101",
19772 => "0000010100100101",
19773 => "0000010100100110",
19774 => "0000010100100110",
19775 => "0000010100100110",
19776 => "0000010100100111",
19777 => "0000010100100111",
19778 => "0000010100100111",
19779 => "0000010100101000",
19780 => "0000010100101000",
19781 => "0000010100101000",
19782 => "0000010100101000",
19783 => "0000010100101001",
19784 => "0000010100101001",
19785 => "0000010100101001",
19786 => "0000010100101010",
19787 => "0000010100101010",
19788 => "0000010100101010",
19789 => "0000010100101011",
19790 => "0000010100101011",
19791 => "0000010100101011",
19792 => "0000010100101100",
19793 => "0000010100101100",
19794 => "0000010100101100",
19795 => "0000010100101100",
19796 => "0000010100101101",
19797 => "0000010100101101",
19798 => "0000010100101101",
19799 => "0000010100101110",
19800 => "0000010100101110",
19801 => "0000010100101110",
19802 => "0000010100101111",
19803 => "0000010100101111",
19804 => "0000010100101111",
19805 => "0000010100110000",
19806 => "0000010100110000",
19807 => "0000010100110000",
19808 => "0000010100110001",
19809 => "0000010100110001",
19810 => "0000010100110001",
19811 => "0000010100110001",
19812 => "0000010100110010",
19813 => "0000010100110010",
19814 => "0000010100110010",
19815 => "0000010100110011",
19816 => "0000010100110011",
19817 => "0000010100110011",
19818 => "0000010100110100",
19819 => "0000010100110100",
19820 => "0000010100110100",
19821 => "0000010100110101",
19822 => "0000010100110101",
19823 => "0000010100110101",
19824 => "0000010100110110",
19825 => "0000010100110110",
19826 => "0000010100110110",
19827 => "0000010100110110",
19828 => "0000010100110111",
19829 => "0000010100110111",
19830 => "0000010100110111",
19831 => "0000010100111000",
19832 => "0000010100111000",
19833 => "0000010100111000",
19834 => "0000010100111001",
19835 => "0000010100111001",
19836 => "0000010100111001",
19837 => "0000010100111010",
19838 => "0000010100111010",
19839 => "0000010100111010",
19840 => "0000010100111011",
19841 => "0000010100111011",
19842 => "0000010100111011",
19843 => "0000010100111011",
19844 => "0000010100111100",
19845 => "0000010100111100",
19846 => "0000010100111100",
19847 => "0000010100111101",
19848 => "0000010100111101",
19849 => "0000010100111101",
19850 => "0000010100111110",
19851 => "0000010100111110",
19852 => "0000010100111110",
19853 => "0000010100111111",
19854 => "0000010100111111",
19855 => "0000010100111111",
19856 => "0000010101000000",
19857 => "0000010101000000",
19858 => "0000010101000000",
19859 => "0000010101000000",
19860 => "0000010101000001",
19861 => "0000010101000001",
19862 => "0000010101000001",
19863 => "0000010101000010",
19864 => "0000010101000010",
19865 => "0000010101000010",
19866 => "0000010101000011",
19867 => "0000010101000011",
19868 => "0000010101000011",
19869 => "0000010101000100",
19870 => "0000010101000100",
19871 => "0000010101000100",
19872 => "0000010101000101",
19873 => "0000010101000101",
19874 => "0000010101000101",
19875 => "0000010101000110",
19876 => "0000010101000110",
19877 => "0000010101000110",
19878 => "0000010101000110",
19879 => "0000010101000111",
19880 => "0000010101000111",
19881 => "0000010101000111",
19882 => "0000010101001000",
19883 => "0000010101001000",
19884 => "0000010101001000",
19885 => "0000010101001001",
19886 => "0000010101001001",
19887 => "0000010101001001",
19888 => "0000010101001010",
19889 => "0000010101001010",
19890 => "0000010101001010",
19891 => "0000010101001011",
19892 => "0000010101001011",
19893 => "0000010101001011",
19894 => "0000010101001100",
19895 => "0000010101001100",
19896 => "0000010101001100",
19897 => "0000010101001101",
19898 => "0000010101001101",
19899 => "0000010101001101",
19900 => "0000010101001101",
19901 => "0000010101001110",
19902 => "0000010101001110",
19903 => "0000010101001110",
19904 => "0000010101001111",
19905 => "0000010101001111",
19906 => "0000010101001111",
19907 => "0000010101010000",
19908 => "0000010101010000",
19909 => "0000010101010000",
19910 => "0000010101010001",
19911 => "0000010101010001",
19912 => "0000010101010001",
19913 => "0000010101010010",
19914 => "0000010101010010",
19915 => "0000010101010010",
19916 => "0000010101010011",
19917 => "0000010101010011",
19918 => "0000010101010011",
19919 => "0000010101010100",
19920 => "0000010101010100",
19921 => "0000010101010100",
19922 => "0000010101010100",
19923 => "0000010101010101",
19924 => "0000010101010101",
19925 => "0000010101010101",
19926 => "0000010101010110",
19927 => "0000010101010110",
19928 => "0000010101010110",
19929 => "0000010101010111",
19930 => "0000010101010111",
19931 => "0000010101010111",
19932 => "0000010101011000",
19933 => "0000010101011000",
19934 => "0000010101011000",
19935 => "0000010101011001",
19936 => "0000010101011001",
19937 => "0000010101011001",
19938 => "0000010101011010",
19939 => "0000010101011010",
19940 => "0000010101011010",
19941 => "0000010101011011",
19942 => "0000010101011011",
19943 => "0000010101011011",
19944 => "0000010101011100",
19945 => "0000010101011100",
19946 => "0000010101011100",
19947 => "0000010101011100",
19948 => "0000010101011101",
19949 => "0000010101011101",
19950 => "0000010101011101",
19951 => "0000010101011110",
19952 => "0000010101011110",
19953 => "0000010101011110",
19954 => "0000010101011111",
19955 => "0000010101011111",
19956 => "0000010101011111",
19957 => "0000010101100000",
19958 => "0000010101100000",
19959 => "0000010101100000",
19960 => "0000010101100001",
19961 => "0000010101100001",
19962 => "0000010101100001",
19963 => "0000010101100010",
19964 => "0000010101100010",
19965 => "0000010101100010",
19966 => "0000010101100011",
19967 => "0000010101100011",
19968 => "0000010101100011",
19969 => "0000010101100100",
19970 => "0000010101100100",
19971 => "0000010101100100",
19972 => "0000010101100101",
19973 => "0000010101100101",
19974 => "0000010101100101",
19975 => "0000010101100101",
19976 => "0000010101100110",
19977 => "0000010101100110",
19978 => "0000010101100110",
19979 => "0000010101100111",
19980 => "0000010101100111",
19981 => "0000010101100111",
19982 => "0000010101101000",
19983 => "0000010101101000",
19984 => "0000010101101000",
19985 => "0000010101101001",
19986 => "0000010101101001",
19987 => "0000010101101001",
19988 => "0000010101101010",
19989 => "0000010101101010",
19990 => "0000010101101010",
19991 => "0000010101101011",
19992 => "0000010101101011",
19993 => "0000010101101011",
19994 => "0000010101101100",
19995 => "0000010101101100",
19996 => "0000010101101100",
19997 => "0000010101101101",
19998 => "0000010101101101",
19999 => "0000010101101101",
20000 => "0000010101101110",
20001 => "0000010101101110",
20002 => "0000010101101110",
20003 => "0000010101101111",
20004 => "0000010101101111",
20005 => "0000010101101111",
20006 => "0000010101110000",
20007 => "0000010101110000",
20008 => "0000010101110000",
20009 => "0000010101110001",
20010 => "0000010101110001",
20011 => "0000010101110001",
20012 => "0000010101110001",
20013 => "0000010101110010",
20014 => "0000010101110010",
20015 => "0000010101110010",
20016 => "0000010101110011",
20017 => "0000010101110011",
20018 => "0000010101110011",
20019 => "0000010101110100",
20020 => "0000010101110100",
20021 => "0000010101110100",
20022 => "0000010101110101",
20023 => "0000010101110101",
20024 => "0000010101110101",
20025 => "0000010101110110",
20026 => "0000010101110110",
20027 => "0000010101110110",
20028 => "0000010101110111",
20029 => "0000010101110111",
20030 => "0000010101110111",
20031 => "0000010101111000",
20032 => "0000010101111000",
20033 => "0000010101111000",
20034 => "0000010101111001",
20035 => "0000010101111001",
20036 => "0000010101111001",
20037 => "0000010101111010",
20038 => "0000010101111010",
20039 => "0000010101111010",
20040 => "0000010101111011",
20041 => "0000010101111011",
20042 => "0000010101111011",
20043 => "0000010101111100",
20044 => "0000010101111100",
20045 => "0000010101111100",
20046 => "0000010101111101",
20047 => "0000010101111101",
20048 => "0000010101111101",
20049 => "0000010101111110",
20050 => "0000010101111110",
20051 => "0000010101111110",
20052 => "0000010101111111",
20053 => "0000010101111111",
20054 => "0000010101111111",
20055 => "0000010110000000",
20056 => "0000010110000000",
20057 => "0000010110000000",
20058 => "0000010110000001",
20059 => "0000010110000001",
20060 => "0000010110000001",
20061 => "0000010110000010",
20062 => "0000010110000010",
20063 => "0000010110000010",
20064 => "0000010110000011",
20065 => "0000010110000011",
20066 => "0000010110000011",
20067 => "0000010110000100",
20068 => "0000010110000100",
20069 => "0000010110000100",
20070 => "0000010110000101",
20071 => "0000010110000101",
20072 => "0000010110000101",
20073 => "0000010110000101",
20074 => "0000010110000110",
20075 => "0000010110000110",
20076 => "0000010110000110",
20077 => "0000010110000111",
20078 => "0000010110000111",
20079 => "0000010110000111",
20080 => "0000010110001000",
20081 => "0000010110001000",
20082 => "0000010110001000",
20083 => "0000010110001001",
20084 => "0000010110001001",
20085 => "0000010110001001",
20086 => "0000010110001010",
20087 => "0000010110001010",
20088 => "0000010110001010",
20089 => "0000010110001011",
20090 => "0000010110001011",
20091 => "0000010110001011",
20092 => "0000010110001100",
20093 => "0000010110001100",
20094 => "0000010110001100",
20095 => "0000010110001101",
20096 => "0000010110001101",
20097 => "0000010110001101",
20098 => "0000010110001110",
20099 => "0000010110001110",
20100 => "0000010110001110",
20101 => "0000010110001111",
20102 => "0000010110001111",
20103 => "0000010110001111",
20104 => "0000010110010000",
20105 => "0000010110010000",
20106 => "0000010110010000",
20107 => "0000010110010001",
20108 => "0000010110010001",
20109 => "0000010110010001",
20110 => "0000010110010010",
20111 => "0000010110010010",
20112 => "0000010110010010",
20113 => "0000010110010011",
20114 => "0000010110010011",
20115 => "0000010110010011",
20116 => "0000010110010100",
20117 => "0000010110010100",
20118 => "0000010110010100",
20119 => "0000010110010101",
20120 => "0000010110010101",
20121 => "0000010110010101",
20122 => "0000010110010110",
20123 => "0000010110010110",
20124 => "0000010110010110",
20125 => "0000010110010111",
20126 => "0000010110010111",
20127 => "0000010110010111",
20128 => "0000010110011000",
20129 => "0000010110011000",
20130 => "0000010110011000",
20131 => "0000010110011001",
20132 => "0000010110011001",
20133 => "0000010110011001",
20134 => "0000010110011010",
20135 => "0000010110011010",
20136 => "0000010110011010",
20137 => "0000010110011011",
20138 => "0000010110011011",
20139 => "0000010110011011",
20140 => "0000010110011100",
20141 => "0000010110011100",
20142 => "0000010110011100",
20143 => "0000010110011101",
20144 => "0000010110011101",
20145 => "0000010110011101",
20146 => "0000010110011110",
20147 => "0000010110011110",
20148 => "0000010110011110",
20149 => "0000010110011111",
20150 => "0000010110011111",
20151 => "0000010110011111",
20152 => "0000010110100000",
20153 => "0000010110100000",
20154 => "0000010110100000",
20155 => "0000010110100001",
20156 => "0000010110100001",
20157 => "0000010110100001",
20158 => "0000010110100010",
20159 => "0000010110100010",
20160 => "0000010110100011",
20161 => "0000010110100011",
20162 => "0000010110100011",
20163 => "0000010110100100",
20164 => "0000010110100100",
20165 => "0000010110100100",
20166 => "0000010110100101",
20167 => "0000010110100101",
20168 => "0000010110100101",
20169 => "0000010110100110",
20170 => "0000010110100110",
20171 => "0000010110100110",
20172 => "0000010110100111",
20173 => "0000010110100111",
20174 => "0000010110100111",
20175 => "0000010110101000",
20176 => "0000010110101000",
20177 => "0000010110101000",
20178 => "0000010110101001",
20179 => "0000010110101001",
20180 => "0000010110101001",
20181 => "0000010110101010",
20182 => "0000010110101010",
20183 => "0000010110101010",
20184 => "0000010110101011",
20185 => "0000010110101011",
20186 => "0000010110101011",
20187 => "0000010110101100",
20188 => "0000010110101100",
20189 => "0000010110101100",
20190 => "0000010110101101",
20191 => "0000010110101101",
20192 => "0000010110101101",
20193 => "0000010110101110",
20194 => "0000010110101110",
20195 => "0000010110101110",
20196 => "0000010110101111",
20197 => "0000010110101111",
20198 => "0000010110101111",
20199 => "0000010110110000",
20200 => "0000010110110000",
20201 => "0000010110110000",
20202 => "0000010110110001",
20203 => "0000010110110001",
20204 => "0000010110110001",
20205 => "0000010110110010",
20206 => "0000010110110010",
20207 => "0000010110110010",
20208 => "0000010110110011",
20209 => "0000010110110011",
20210 => "0000010110110011",
20211 => "0000010110110100",
20212 => "0000010110110100",
20213 => "0000010110110100",
20214 => "0000010110110101",
20215 => "0000010110110101",
20216 => "0000010110110101",
20217 => "0000010110110110",
20218 => "0000010110110110",
20219 => "0000010110110111",
20220 => "0000010110110111",
20221 => "0000010110110111",
20222 => "0000010110111000",
20223 => "0000010110111000",
20224 => "0000010110111000",
20225 => "0000010110111001",
20226 => "0000010110111001",
20227 => "0000010110111001",
20228 => "0000010110111010",
20229 => "0000010110111010",
20230 => "0000010110111010",
20231 => "0000010110111011",
20232 => "0000010110111011",
20233 => "0000010110111011",
20234 => "0000010110111100",
20235 => "0000010110111100",
20236 => "0000010110111100",
20237 => "0000010110111101",
20238 => "0000010110111101",
20239 => "0000010110111101",
20240 => "0000010110111110",
20241 => "0000010110111110",
20242 => "0000010110111110",
20243 => "0000010110111111",
20244 => "0000010110111111",
20245 => "0000010110111111",
20246 => "0000010111000000",
20247 => "0000010111000000",
20248 => "0000010111000000",
20249 => "0000010111000001",
20250 => "0000010111000001",
20251 => "0000010111000001",
20252 => "0000010111000010",
20253 => "0000010111000010",
20254 => "0000010111000010",
20255 => "0000010111000011",
20256 => "0000010111000011",
20257 => "0000010111000100",
20258 => "0000010111000100",
20259 => "0000010111000100",
20260 => "0000010111000101",
20261 => "0000010111000101",
20262 => "0000010111000101",
20263 => "0000010111000110",
20264 => "0000010111000110",
20265 => "0000010111000110",
20266 => "0000010111000111",
20267 => "0000010111000111",
20268 => "0000010111000111",
20269 => "0000010111001000",
20270 => "0000010111001000",
20271 => "0000010111001000",
20272 => "0000010111001001",
20273 => "0000010111001001",
20274 => "0000010111001001",
20275 => "0000010111001010",
20276 => "0000010111001010",
20277 => "0000010111001010",
20278 => "0000010111001011",
20279 => "0000010111001011",
20280 => "0000010111001011",
20281 => "0000010111001100",
20282 => "0000010111001100",
20283 => "0000010111001100",
20284 => "0000010111001101",
20285 => "0000010111001101",
20286 => "0000010111001110",
20287 => "0000010111001110",
20288 => "0000010111001110",
20289 => "0000010111001111",
20290 => "0000010111001111",
20291 => "0000010111001111",
20292 => "0000010111010000",
20293 => "0000010111010000",
20294 => "0000010111010000",
20295 => "0000010111010001",
20296 => "0000010111010001",
20297 => "0000010111010001",
20298 => "0000010111010010",
20299 => "0000010111010010",
20300 => "0000010111010010",
20301 => "0000010111010011",
20302 => "0000010111010011",
20303 => "0000010111010011",
20304 => "0000010111010100",
20305 => "0000010111010100",
20306 => "0000010111010100",
20307 => "0000010111010101",
20308 => "0000010111010101",
20309 => "0000010111010110",
20310 => "0000010111010110",
20311 => "0000010111010110",
20312 => "0000010111010111",
20313 => "0000010111010111",
20314 => "0000010111010111",
20315 => "0000010111011000",
20316 => "0000010111011000",
20317 => "0000010111011000",
20318 => "0000010111011001",
20319 => "0000010111011001",
20320 => "0000010111011001",
20321 => "0000010111011010",
20322 => "0000010111011010",
20323 => "0000010111011010",
20324 => "0000010111011011",
20325 => "0000010111011011",
20326 => "0000010111011011",
20327 => "0000010111011100",
20328 => "0000010111011100",
20329 => "0000010111011100",
20330 => "0000010111011101",
20331 => "0000010111011101",
20332 => "0000010111011110",
20333 => "0000010111011110",
20334 => "0000010111011110",
20335 => "0000010111011111",
20336 => "0000010111011111",
20337 => "0000010111011111",
20338 => "0000010111100000",
20339 => "0000010111100000",
20340 => "0000010111100000",
20341 => "0000010111100001",
20342 => "0000010111100001",
20343 => "0000010111100001",
20344 => "0000010111100010",
20345 => "0000010111100010",
20346 => "0000010111100010",
20347 => "0000010111100011",
20348 => "0000010111100011",
20349 => "0000010111100011",
20350 => "0000010111100100",
20351 => "0000010111100100",
20352 => "0000010111100101",
20353 => "0000010111100101",
20354 => "0000010111100101",
20355 => "0000010111100110",
20356 => "0000010111100110",
20357 => "0000010111100110",
20358 => "0000010111100111",
20359 => "0000010111100111",
20360 => "0000010111100111",
20361 => "0000010111101000",
20362 => "0000010111101000",
20363 => "0000010111101000",
20364 => "0000010111101001",
20365 => "0000010111101001",
20366 => "0000010111101001",
20367 => "0000010111101010",
20368 => "0000010111101010",
20369 => "0000010111101011",
20370 => "0000010111101011",
20371 => "0000010111101011",
20372 => "0000010111101100",
20373 => "0000010111101100",
20374 => "0000010111101100",
20375 => "0000010111101101",
20376 => "0000010111101101",
20377 => "0000010111101101",
20378 => "0000010111101110",
20379 => "0000010111101110",
20380 => "0000010111101110",
20381 => "0000010111101111",
20382 => "0000010111101111",
20383 => "0000010111101111",
20384 => "0000010111110000",
20385 => "0000010111110000",
20386 => "0000010111110001",
20387 => "0000010111110001",
20388 => "0000010111110001",
20389 => "0000010111110010",
20390 => "0000010111110010",
20391 => "0000010111110010",
20392 => "0000010111110011",
20393 => "0000010111110011",
20394 => "0000010111110011",
20395 => "0000010111110100",
20396 => "0000010111110100",
20397 => "0000010111110100",
20398 => "0000010111110101",
20399 => "0000010111110101",
20400 => "0000010111110110",
20401 => "0000010111110110",
20402 => "0000010111110110",
20403 => "0000010111110111",
20404 => "0000010111110111",
20405 => "0000010111110111",
20406 => "0000010111111000",
20407 => "0000010111111000",
20408 => "0000010111111000",
20409 => "0000010111111001",
20410 => "0000010111111001",
20411 => "0000010111111001",
20412 => "0000010111111010",
20413 => "0000010111111010",
20414 => "0000010111111010",
20415 => "0000010111111011",
20416 => "0000010111111011",
20417 => "0000010111111100",
20418 => "0000010111111100",
20419 => "0000010111111100",
20420 => "0000010111111101",
20421 => "0000010111111101",
20422 => "0000010111111101",
20423 => "0000010111111110",
20424 => "0000010111111110",
20425 => "0000010111111110",
20426 => "0000010111111111",
20427 => "0000010111111111",
20428 => "0000010111111111",
20429 => "0000011000000000",
20430 => "0000011000000000",
20431 => "0000011000000001",
20432 => "0000011000000001",
20433 => "0000011000000001",
20434 => "0000011000000010",
20435 => "0000011000000010",
20436 => "0000011000000010",
20437 => "0000011000000011",
20438 => "0000011000000011",
20439 => "0000011000000011",
20440 => "0000011000000100",
20441 => "0000011000000100",
20442 => "0000011000000100",
20443 => "0000011000000101",
20444 => "0000011000000101",
20445 => "0000011000000110",
20446 => "0000011000000110",
20447 => "0000011000000110",
20448 => "0000011000000111",
20449 => "0000011000000111",
20450 => "0000011000000111",
20451 => "0000011000001000",
20452 => "0000011000001000",
20453 => "0000011000001000",
20454 => "0000011000001001",
20455 => "0000011000001001",
20456 => "0000011000001010",
20457 => "0000011000001010",
20458 => "0000011000001010",
20459 => "0000011000001011",
20460 => "0000011000001011",
20461 => "0000011000001011",
20462 => "0000011000001100",
20463 => "0000011000001100",
20464 => "0000011000001100",
20465 => "0000011000001101",
20466 => "0000011000001101",
20467 => "0000011000001101",
20468 => "0000011000001110",
20469 => "0000011000001110",
20470 => "0000011000001111",
20471 => "0000011000001111",
20472 => "0000011000001111",
20473 => "0000011000010000",
20474 => "0000011000010000",
20475 => "0000011000010000",
20476 => "0000011000010001",
20477 => "0000011000010001",
20478 => "0000011000010001",
20479 => "0000011000010010",
20480 => "0000011000010010",
20481 => "0000011000010011",
20482 => "0000011000010011",
20483 => "0000011000010011",
20484 => "0000011000010100",
20485 => "0000011000010100",
20486 => "0000011000010100",
20487 => "0000011000010101",
20488 => "0000011000010101",
20489 => "0000011000010101",
20490 => "0000011000010110",
20491 => "0000011000010110",
20492 => "0000011000010111",
20493 => "0000011000010111",
20494 => "0000011000010111",
20495 => "0000011000011000",
20496 => "0000011000011000",
20497 => "0000011000011000",
20498 => "0000011000011001",
20499 => "0000011000011001",
20500 => "0000011000011001",
20501 => "0000011000011010",
20502 => "0000011000011010",
20503 => "0000011000011010",
20504 => "0000011000011011",
20505 => "0000011000011011",
20506 => "0000011000011100",
20507 => "0000011000011100",
20508 => "0000011000011100",
20509 => "0000011000011101",
20510 => "0000011000011101",
20511 => "0000011000011101",
20512 => "0000011000011110",
20513 => "0000011000011110",
20514 => "0000011000011110",
20515 => "0000011000011111",
20516 => "0000011000011111",
20517 => "0000011000100000",
20518 => "0000011000100000",
20519 => "0000011000100000",
20520 => "0000011000100001",
20521 => "0000011000100001",
20522 => "0000011000100001",
20523 => "0000011000100010",
20524 => "0000011000100010",
20525 => "0000011000100011",
20526 => "0000011000100011",
20527 => "0000011000100011",
20528 => "0000011000100100",
20529 => "0000011000100100",
20530 => "0000011000100100",
20531 => "0000011000100101",
20532 => "0000011000100101",
20533 => "0000011000100101",
20534 => "0000011000100110",
20535 => "0000011000100110",
20536 => "0000011000100111",
20537 => "0000011000100111",
20538 => "0000011000100111",
20539 => "0000011000101000",
20540 => "0000011000101000",
20541 => "0000011000101000",
20542 => "0000011000101001",
20543 => "0000011000101001",
20544 => "0000011000101001",
20545 => "0000011000101010",
20546 => "0000011000101010",
20547 => "0000011000101011",
20548 => "0000011000101011",
20549 => "0000011000101011",
20550 => "0000011000101100",
20551 => "0000011000101100",
20552 => "0000011000101100",
20553 => "0000011000101101",
20554 => "0000011000101101",
20555 => "0000011000101101",
20556 => "0000011000101110",
20557 => "0000011000101110",
20558 => "0000011000101111",
20559 => "0000011000101111",
20560 => "0000011000101111",
20561 => "0000011000110000",
20562 => "0000011000110000",
20563 => "0000011000110000",
20564 => "0000011000110001",
20565 => "0000011000110001",
20566 => "0000011000110010",
20567 => "0000011000110010",
20568 => "0000011000110010",
20569 => "0000011000110011",
20570 => "0000011000110011",
20571 => "0000011000110011",
20572 => "0000011000110100",
20573 => "0000011000110100",
20574 => "0000011000110100",
20575 => "0000011000110101",
20576 => "0000011000110101",
20577 => "0000011000110110",
20578 => "0000011000110110",
20579 => "0000011000110110",
20580 => "0000011000110111",
20581 => "0000011000110111",
20582 => "0000011000110111",
20583 => "0000011000111000",
20584 => "0000011000111000",
20585 => "0000011000111001",
20586 => "0000011000111001",
20587 => "0000011000111001",
20588 => "0000011000111010",
20589 => "0000011000111010",
20590 => "0000011000111010",
20591 => "0000011000111011",
20592 => "0000011000111011",
20593 => "0000011000111100",
20594 => "0000011000111100",
20595 => "0000011000111100",
20596 => "0000011000111101",
20597 => "0000011000111101",
20598 => "0000011000111101",
20599 => "0000011000111110",
20600 => "0000011000111110",
20601 => "0000011000111110",
20602 => "0000011000111111",
20603 => "0000011000111111",
20604 => "0000011001000000",
20605 => "0000011001000000",
20606 => "0000011001000000",
20607 => "0000011001000001",
20608 => "0000011001000001",
20609 => "0000011001000001",
20610 => "0000011001000010",
20611 => "0000011001000010",
20612 => "0000011001000011",
20613 => "0000011001000011",
20614 => "0000011001000011",
20615 => "0000011001000100",
20616 => "0000011001000100",
20617 => "0000011001000100",
20618 => "0000011001000101",
20619 => "0000011001000101",
20620 => "0000011001000110",
20621 => "0000011001000110",
20622 => "0000011001000110",
20623 => "0000011001000111",
20624 => "0000011001000111",
20625 => "0000011001000111",
20626 => "0000011001001000",
20627 => "0000011001001000",
20628 => "0000011001001001",
20629 => "0000011001001001",
20630 => "0000011001001001",
20631 => "0000011001001010",
20632 => "0000011001001010",
20633 => "0000011001001010",
20634 => "0000011001001011",
20635 => "0000011001001011",
20636 => "0000011001001100",
20637 => "0000011001001100",
20638 => "0000011001001100",
20639 => "0000011001001101",
20640 => "0000011001001101",
20641 => "0000011001001101",
20642 => "0000011001001110",
20643 => "0000011001001110",
20644 => "0000011001001111",
20645 => "0000011001001111",
20646 => "0000011001001111",
20647 => "0000011001010000",
20648 => "0000011001010000",
20649 => "0000011001010000",
20650 => "0000011001010001",
20651 => "0000011001010001",
20652 => "0000011001010010",
20653 => "0000011001010010",
20654 => "0000011001010010",
20655 => "0000011001010011",
20656 => "0000011001010011",
20657 => "0000011001010011",
20658 => "0000011001010100",
20659 => "0000011001010100",
20660 => "0000011001010101",
20661 => "0000011001010101",
20662 => "0000011001010101",
20663 => "0000011001010110",
20664 => "0000011001010110",
20665 => "0000011001010110",
20666 => "0000011001010111",
20667 => "0000011001010111",
20668 => "0000011001011000",
20669 => "0000011001011000",
20670 => "0000011001011000",
20671 => "0000011001011001",
20672 => "0000011001011001",
20673 => "0000011001011001",
20674 => "0000011001011010",
20675 => "0000011001011010",
20676 => "0000011001011011",
20677 => "0000011001011011",
20678 => "0000011001011011",
20679 => "0000011001011100",
20680 => "0000011001011100",
20681 => "0000011001011100",
20682 => "0000011001011101",
20683 => "0000011001011101",
20684 => "0000011001011110",
20685 => "0000011001011110",
20686 => "0000011001011110",
20687 => "0000011001011111",
20688 => "0000011001011111",
20689 => "0000011001011111",
20690 => "0000011001100000",
20691 => "0000011001100000",
20692 => "0000011001100001",
20693 => "0000011001100001",
20694 => "0000011001100001",
20695 => "0000011001100010",
20696 => "0000011001100010",
20697 => "0000011001100011",
20698 => "0000011001100011",
20699 => "0000011001100011",
20700 => "0000011001100100",
20701 => "0000011001100100",
20702 => "0000011001100100",
20703 => "0000011001100101",
20704 => "0000011001100101",
20705 => "0000011001100110",
20706 => "0000011001100110",
20707 => "0000011001100110",
20708 => "0000011001100111",
20709 => "0000011001100111",
20710 => "0000011001100111",
20711 => "0000011001101000",
20712 => "0000011001101000",
20713 => "0000011001101001",
20714 => "0000011001101001",
20715 => "0000011001101001",
20716 => "0000011001101010",
20717 => "0000011001101010",
20718 => "0000011001101010",
20719 => "0000011001101011",
20720 => "0000011001101011",
20721 => "0000011001101100",
20722 => "0000011001101100",
20723 => "0000011001101100",
20724 => "0000011001101101",
20725 => "0000011001101101",
20726 => "0000011001101110",
20727 => "0000011001101110",
20728 => "0000011001101110",
20729 => "0000011001101111",
20730 => "0000011001101111",
20731 => "0000011001101111",
20732 => "0000011001110000",
20733 => "0000011001110000",
20734 => "0000011001110001",
20735 => "0000011001110001",
20736 => "0000011001110001",
20737 => "0000011001110010",
20738 => "0000011001110010",
20739 => "0000011001110011",
20740 => "0000011001110011",
20741 => "0000011001110011",
20742 => "0000011001110100",
20743 => "0000011001110100",
20744 => "0000011001110100",
20745 => "0000011001110101",
20746 => "0000011001110101",
20747 => "0000011001110110",
20748 => "0000011001110110",
20749 => "0000011001110110",
20750 => "0000011001110111",
20751 => "0000011001110111",
20752 => "0000011001110111",
20753 => "0000011001111000",
20754 => "0000011001111000",
20755 => "0000011001111001",
20756 => "0000011001111001",
20757 => "0000011001111001",
20758 => "0000011001111010",
20759 => "0000011001111010",
20760 => "0000011001111011",
20761 => "0000011001111011",
20762 => "0000011001111011",
20763 => "0000011001111100",
20764 => "0000011001111100",
20765 => "0000011001111100",
20766 => "0000011001111101",
20767 => "0000011001111101",
20768 => "0000011001111110",
20769 => "0000011001111110",
20770 => "0000011001111110",
20771 => "0000011001111111",
20772 => "0000011001111111",
20773 => "0000011010000000",
20774 => "0000011010000000",
20775 => "0000011010000000",
20776 => "0000011010000001",
20777 => "0000011010000001",
20778 => "0000011010000001",
20779 => "0000011010000010",
20780 => "0000011010000010",
20781 => "0000011010000011",
20782 => "0000011010000011",
20783 => "0000011010000011",
20784 => "0000011010000100",
20785 => "0000011010000100",
20786 => "0000011010000101",
20787 => "0000011010000101",
20788 => "0000011010000101",
20789 => "0000011010000110",
20790 => "0000011010000110",
20791 => "0000011010000111",
20792 => "0000011010000111",
20793 => "0000011010000111",
20794 => "0000011010001000",
20795 => "0000011010001000",
20796 => "0000011010001000",
20797 => "0000011010001001",
20798 => "0000011010001001",
20799 => "0000011010001010",
20800 => "0000011010001010",
20801 => "0000011010001010",
20802 => "0000011010001011",
20803 => "0000011010001011",
20804 => "0000011010001100",
20805 => "0000011010001100",
20806 => "0000011010001100",
20807 => "0000011010001101",
20808 => "0000011010001101",
20809 => "0000011010001101",
20810 => "0000011010001110",
20811 => "0000011010001110",
20812 => "0000011010001111",
20813 => "0000011010001111",
20814 => "0000011010001111",
20815 => "0000011010010000",
20816 => "0000011010010000",
20817 => "0000011010010001",
20818 => "0000011010010001",
20819 => "0000011010010001",
20820 => "0000011010010010",
20821 => "0000011010010010",
20822 => "0000011010010011",
20823 => "0000011010010011",
20824 => "0000011010010011",
20825 => "0000011010010100",
20826 => "0000011010010100",
20827 => "0000011010010101",
20828 => "0000011010010101",
20829 => "0000011010010101",
20830 => "0000011010010110",
20831 => "0000011010010110",
20832 => "0000011010010110",
20833 => "0000011010010111",
20834 => "0000011010010111",
20835 => "0000011010011000",
20836 => "0000011010011000",
20837 => "0000011010011000",
20838 => "0000011010011001",
20839 => "0000011010011001",
20840 => "0000011010011010",
20841 => "0000011010011010",
20842 => "0000011010011010",
20843 => "0000011010011011",
20844 => "0000011010011011",
20845 => "0000011010011100",
20846 => "0000011010011100",
20847 => "0000011010011100",
20848 => "0000011010011101",
20849 => "0000011010011101",
20850 => "0000011010011101",
20851 => "0000011010011110",
20852 => "0000011010011110",
20853 => "0000011010011111",
20854 => "0000011010011111",
20855 => "0000011010011111",
20856 => "0000011010100000",
20857 => "0000011010100000",
20858 => "0000011010100001",
20859 => "0000011010100001",
20860 => "0000011010100001",
20861 => "0000011010100010",
20862 => "0000011010100010",
20863 => "0000011010100011",
20864 => "0000011010100011",
20865 => "0000011010100011",
20866 => "0000011010100100",
20867 => "0000011010100100",
20868 => "0000011010100101",
20869 => "0000011010100101",
20870 => "0000011010100101",
20871 => "0000011010100110",
20872 => "0000011010100110",
20873 => "0000011010100111",
20874 => "0000011010100111",
20875 => "0000011010100111",
20876 => "0000011010101000",
20877 => "0000011010101000",
20878 => "0000011010101001",
20879 => "0000011010101001",
20880 => "0000011010101001",
20881 => "0000011010101010",
20882 => "0000011010101010",
20883 => "0000011010101010",
20884 => "0000011010101011",
20885 => "0000011010101011",
20886 => "0000011010101100",
20887 => "0000011010101100",
20888 => "0000011010101100",
20889 => "0000011010101101",
20890 => "0000011010101101",
20891 => "0000011010101110",
20892 => "0000011010101110",
20893 => "0000011010101110",
20894 => "0000011010101111",
20895 => "0000011010101111",
20896 => "0000011010110000",
20897 => "0000011010110000",
20898 => "0000011010110000",
20899 => "0000011010110001",
20900 => "0000011010110001",
20901 => "0000011010110010",
20902 => "0000011010110010",
20903 => "0000011010110010",
20904 => "0000011010110011",
20905 => "0000011010110011",
20906 => "0000011010110100",
20907 => "0000011010110100",
20908 => "0000011010110100",
20909 => "0000011010110101",
20910 => "0000011010110101",
20911 => "0000011010110110",
20912 => "0000011010110110",
20913 => "0000011010110110",
20914 => "0000011010110111",
20915 => "0000011010110111",
20916 => "0000011010111000",
20917 => "0000011010111000",
20918 => "0000011010111000",
20919 => "0000011010111001",
20920 => "0000011010111001",
20921 => "0000011010111010",
20922 => "0000011010111010",
20923 => "0000011010111010",
20924 => "0000011010111011",
20925 => "0000011010111011",
20926 => "0000011010111100",
20927 => "0000011010111100",
20928 => "0000011010111100",
20929 => "0000011010111101",
20930 => "0000011010111101",
20931 => "0000011010111110",
20932 => "0000011010111110",
20933 => "0000011010111110",
20934 => "0000011010111111",
20935 => "0000011010111111",
20936 => "0000011011000000",
20937 => "0000011011000000",
20938 => "0000011011000000",
20939 => "0000011011000001",
20940 => "0000011011000001",
20941 => "0000011011000010",
20942 => "0000011011000010",
20943 => "0000011011000010",
20944 => "0000011011000011",
20945 => "0000011011000011",
20946 => "0000011011000100",
20947 => "0000011011000100",
20948 => "0000011011000100",
20949 => "0000011011000101",
20950 => "0000011011000101",
20951 => "0000011011000110",
20952 => "0000011011000110",
20953 => "0000011011000110",
20954 => "0000011011000111",
20955 => "0000011011000111",
20956 => "0000011011001000",
20957 => "0000011011001000",
20958 => "0000011011001000",
20959 => "0000011011001001",
20960 => "0000011011001001",
20961 => "0000011011001010",
20962 => "0000011011001010",
20963 => "0000011011001010",
20964 => "0000011011001011",
20965 => "0000011011001011",
20966 => "0000011011001100",
20967 => "0000011011001100",
20968 => "0000011011001100",
20969 => "0000011011001101",
20970 => "0000011011001101",
20971 => "0000011011001110",
20972 => "0000011011001110",
20973 => "0000011011001110",
20974 => "0000011011001111",
20975 => "0000011011001111",
20976 => "0000011011010000",
20977 => "0000011011010000",
20978 => "0000011011010000",
20979 => "0000011011010001",
20980 => "0000011011010001",
20981 => "0000011011010010",
20982 => "0000011011010010",
20983 => "0000011011010010",
20984 => "0000011011010011",
20985 => "0000011011010011",
20986 => "0000011011010100",
20987 => "0000011011010100",
20988 => "0000011011010100",
20989 => "0000011011010101",
20990 => "0000011011010101",
20991 => "0000011011010110",
20992 => "0000011011010110",
20993 => "0000011011010110",
20994 => "0000011011010111",
20995 => "0000011011010111",
20996 => "0000011011011000",
20997 => "0000011011011000",
20998 => "0000011011011000",
20999 => "0000011011011001",
21000 => "0000011011011001",
21001 => "0000011011011010",
21002 => "0000011011011010",
21003 => "0000011011011011",
21004 => "0000011011011011",
21005 => "0000011011011011",
21006 => "0000011011011100",
21007 => "0000011011011100",
21008 => "0000011011011101",
21009 => "0000011011011101",
21010 => "0000011011011101",
21011 => "0000011011011110",
21012 => "0000011011011110",
21013 => "0000011011011111",
21014 => "0000011011011111",
21015 => "0000011011011111",
21016 => "0000011011100000",
21017 => "0000011011100000",
21018 => "0000011011100001",
21019 => "0000011011100001",
21020 => "0000011011100001",
21021 => "0000011011100010",
21022 => "0000011011100010",
21023 => "0000011011100011",
21024 => "0000011011100011",
21025 => "0000011011100011",
21026 => "0000011011100100",
21027 => "0000011011100100",
21028 => "0000011011100101",
21029 => "0000011011100101",
21030 => "0000011011100101",
21031 => "0000011011100110",
21032 => "0000011011100110",
21033 => "0000011011100111",
21034 => "0000011011100111",
21035 => "0000011011101000",
21036 => "0000011011101000",
21037 => "0000011011101000",
21038 => "0000011011101001",
21039 => "0000011011101001",
21040 => "0000011011101010",
21041 => "0000011011101010",
21042 => "0000011011101010",
21043 => "0000011011101011",
21044 => "0000011011101011",
21045 => "0000011011101100",
21046 => "0000011011101100",
21047 => "0000011011101100",
21048 => "0000011011101101",
21049 => "0000011011101101",
21050 => "0000011011101110",
21051 => "0000011011101110",
21052 => "0000011011101110",
21053 => "0000011011101111",
21054 => "0000011011101111",
21055 => "0000011011110000",
21056 => "0000011011110000",
21057 => "0000011011110001",
21058 => "0000011011110001",
21059 => "0000011011110001",
21060 => "0000011011110010",
21061 => "0000011011110010",
21062 => "0000011011110011",
21063 => "0000011011110011",
21064 => "0000011011110011",
21065 => "0000011011110100",
21066 => "0000011011110100",
21067 => "0000011011110101",
21068 => "0000011011110101",
21069 => "0000011011110101",
21070 => "0000011011110110",
21071 => "0000011011110110",
21072 => "0000011011110111",
21073 => "0000011011110111",
21074 => "0000011011111000",
21075 => "0000011011111000",
21076 => "0000011011111000",
21077 => "0000011011111001",
21078 => "0000011011111001",
21079 => "0000011011111010",
21080 => "0000011011111010",
21081 => "0000011011111010",
21082 => "0000011011111011",
21083 => "0000011011111011",
21084 => "0000011011111100",
21085 => "0000011011111100",
21086 => "0000011011111100",
21087 => "0000011011111101",
21088 => "0000011011111101",
21089 => "0000011011111110",
21090 => "0000011011111110",
21091 => "0000011011111111",
21092 => "0000011011111111",
21093 => "0000011011111111",
21094 => "0000011100000000",
21095 => "0000011100000000",
21096 => "0000011100000001",
21097 => "0000011100000001",
21098 => "0000011100000001",
21099 => "0000011100000010",
21100 => "0000011100000010",
21101 => "0000011100000011",
21102 => "0000011100000011",
21103 => "0000011100000011",
21104 => "0000011100000100",
21105 => "0000011100000100",
21106 => "0000011100000101",
21107 => "0000011100000101",
21108 => "0000011100000110",
21109 => "0000011100000110",
21110 => "0000011100000110",
21111 => "0000011100000111",
21112 => "0000011100000111",
21113 => "0000011100001000",
21114 => "0000011100001000",
21115 => "0000011100001000",
21116 => "0000011100001001",
21117 => "0000011100001001",
21118 => "0000011100001010",
21119 => "0000011100001010",
21120 => "0000011100001011",
21121 => "0000011100001011",
21122 => "0000011100001011",
21123 => "0000011100001100",
21124 => "0000011100001100",
21125 => "0000011100001101",
21126 => "0000011100001101",
21127 => "0000011100001101",
21128 => "0000011100001110",
21129 => "0000011100001110",
21130 => "0000011100001111",
21131 => "0000011100001111",
21132 => "0000011100010000",
21133 => "0000011100010000",
21134 => "0000011100010000",
21135 => "0000011100010001",
21136 => "0000011100010001",
21137 => "0000011100010010",
21138 => "0000011100010010",
21139 => "0000011100010010",
21140 => "0000011100010011",
21141 => "0000011100010011",
21142 => "0000011100010100",
21143 => "0000011100010100",
21144 => "0000011100010101",
21145 => "0000011100010101",
21146 => "0000011100010101",
21147 => "0000011100010110",
21148 => "0000011100010110",
21149 => "0000011100010111",
21150 => "0000011100010111",
21151 => "0000011100010111",
21152 => "0000011100011000",
21153 => "0000011100011000",
21154 => "0000011100011001",
21155 => "0000011100011001",
21156 => "0000011100011010",
21157 => "0000011100011010",
21158 => "0000011100011010",
21159 => "0000011100011011",
21160 => "0000011100011011",
21161 => "0000011100011100",
21162 => "0000011100011100",
21163 => "0000011100011101",
21164 => "0000011100011101",
21165 => "0000011100011101",
21166 => "0000011100011110",
21167 => "0000011100011110",
21168 => "0000011100011111",
21169 => "0000011100011111",
21170 => "0000011100011111",
21171 => "0000011100100000",
21172 => "0000011100100000",
21173 => "0000011100100001",
21174 => "0000011100100001",
21175 => "0000011100100010",
21176 => "0000011100100010",
21177 => "0000011100100010",
21178 => "0000011100100011",
21179 => "0000011100100011",
21180 => "0000011100100100",
21181 => "0000011100100100",
21182 => "0000011100100101",
21183 => "0000011100100101",
21184 => "0000011100100101",
21185 => "0000011100100110",
21186 => "0000011100100110",
21187 => "0000011100100111",
21188 => "0000011100100111",
21189 => "0000011100100111",
21190 => "0000011100101000",
21191 => "0000011100101000",
21192 => "0000011100101001",
21193 => "0000011100101001",
21194 => "0000011100101010",
21195 => "0000011100101010",
21196 => "0000011100101010",
21197 => "0000011100101011",
21198 => "0000011100101011",
21199 => "0000011100101100",
21200 => "0000011100101100",
21201 => "0000011100101101",
21202 => "0000011100101101",
21203 => "0000011100101101",
21204 => "0000011100101110",
21205 => "0000011100101110",
21206 => "0000011100101111",
21207 => "0000011100101111",
21208 => "0000011100101111",
21209 => "0000011100110000",
21210 => "0000011100110000",
21211 => "0000011100110001",
21212 => "0000011100110001",
21213 => "0000011100110010",
21214 => "0000011100110010",
21215 => "0000011100110010",
21216 => "0000011100110011",
21217 => "0000011100110011",
21218 => "0000011100110100",
21219 => "0000011100110100",
21220 => "0000011100110101",
21221 => "0000011100110101",
21222 => "0000011100110101",
21223 => "0000011100110110",
21224 => "0000011100110110",
21225 => "0000011100110111",
21226 => "0000011100110111",
21227 => "0000011100111000",
21228 => "0000011100111000",
21229 => "0000011100111000",
21230 => "0000011100111001",
21231 => "0000011100111001",
21232 => "0000011100111010",
21233 => "0000011100111010",
21234 => "0000011100111011",
21235 => "0000011100111011",
21236 => "0000011100111011",
21237 => "0000011100111100",
21238 => "0000011100111100",
21239 => "0000011100111101",
21240 => "0000011100111101",
21241 => "0000011100111110",
21242 => "0000011100111110",
21243 => "0000011100111110",
21244 => "0000011100111111",
21245 => "0000011100111111",
21246 => "0000011101000000",
21247 => "0000011101000000",
21248 => "0000011101000001",
21249 => "0000011101000001",
21250 => "0000011101000001",
21251 => "0000011101000010",
21252 => "0000011101000010",
21253 => "0000011101000011",
21254 => "0000011101000011",
21255 => "0000011101000100",
21256 => "0000011101000100",
21257 => "0000011101000100",
21258 => "0000011101000101",
21259 => "0000011101000101",
21260 => "0000011101000110",
21261 => "0000011101000110",
21262 => "0000011101000111",
21263 => "0000011101000111",
21264 => "0000011101000111",
21265 => "0000011101001000",
21266 => "0000011101001000",
21267 => "0000011101001001",
21268 => "0000011101001001",
21269 => "0000011101001010",
21270 => "0000011101001010",
21271 => "0000011101001010",
21272 => "0000011101001011",
21273 => "0000011101001011",
21274 => "0000011101001100",
21275 => "0000011101001100",
21276 => "0000011101001101",
21277 => "0000011101001101",
21278 => "0000011101001101",
21279 => "0000011101001110",
21280 => "0000011101001110",
21281 => "0000011101001111",
21282 => "0000011101001111",
21283 => "0000011101010000",
21284 => "0000011101010000",
21285 => "0000011101010000",
21286 => "0000011101010001",
21287 => "0000011101010001",
21288 => "0000011101010010",
21289 => "0000011101010010",
21290 => "0000011101010011",
21291 => "0000011101010011",
21292 => "0000011101010011",
21293 => "0000011101010100",
21294 => "0000011101010100",
21295 => "0000011101010101",
21296 => "0000011101010101",
21297 => "0000011101010110",
21298 => "0000011101010110",
21299 => "0000011101010110",
21300 => "0000011101010111",
21301 => "0000011101010111",
21302 => "0000011101011000",
21303 => "0000011101011000",
21304 => "0000011101011001",
21305 => "0000011101011001",
21306 => "0000011101011001",
21307 => "0000011101011010",
21308 => "0000011101011010",
21309 => "0000011101011011",
21310 => "0000011101011011",
21311 => "0000011101011100",
21312 => "0000011101011100",
21313 => "0000011101011101",
21314 => "0000011101011101",
21315 => "0000011101011101",
21316 => "0000011101011110",
21317 => "0000011101011110",
21318 => "0000011101011111",
21319 => "0000011101011111",
21320 => "0000011101100000",
21321 => "0000011101100000",
21322 => "0000011101100000",
21323 => "0000011101100001",
21324 => "0000011101100001",
21325 => "0000011101100010",
21326 => "0000011101100010",
21327 => "0000011101100011",
21328 => "0000011101100011",
21329 => "0000011101100011",
21330 => "0000011101100100",
21331 => "0000011101100100",
21332 => "0000011101100101",
21333 => "0000011101100101",
21334 => "0000011101100110",
21335 => "0000011101100110",
21336 => "0000011101100111",
21337 => "0000011101100111",
21338 => "0000011101100111",
21339 => "0000011101101000",
21340 => "0000011101101000",
21341 => "0000011101101001",
21342 => "0000011101101001",
21343 => "0000011101101010",
21344 => "0000011101101010",
21345 => "0000011101101010",
21346 => "0000011101101011",
21347 => "0000011101101011",
21348 => "0000011101101100",
21349 => "0000011101101100",
21350 => "0000011101101101",
21351 => "0000011101101101",
21352 => "0000011101101101",
21353 => "0000011101101110",
21354 => "0000011101101110",
21355 => "0000011101101111",
21356 => "0000011101101111",
21357 => "0000011101110000",
21358 => "0000011101110000",
21359 => "0000011101110001",
21360 => "0000011101110001",
21361 => "0000011101110001",
21362 => "0000011101110010",
21363 => "0000011101110010",
21364 => "0000011101110011",
21365 => "0000011101110011",
21366 => "0000011101110100",
21367 => "0000011101110100",
21368 => "0000011101110101",
21369 => "0000011101110101",
21370 => "0000011101110101",
21371 => "0000011101110110",
21372 => "0000011101110110",
21373 => "0000011101110111",
21374 => "0000011101110111",
21375 => "0000011101111000",
21376 => "0000011101111000",
21377 => "0000011101111000",
21378 => "0000011101111001",
21379 => "0000011101111001",
21380 => "0000011101111010",
21381 => "0000011101111010",
21382 => "0000011101111011",
21383 => "0000011101111011",
21384 => "0000011101111100",
21385 => "0000011101111100",
21386 => "0000011101111100",
21387 => "0000011101111101",
21388 => "0000011101111101",
21389 => "0000011101111110",
21390 => "0000011101111110",
21391 => "0000011101111111",
21392 => "0000011101111111",
21393 => "0000011110000000",
21394 => "0000011110000000",
21395 => "0000011110000000",
21396 => "0000011110000001",
21397 => "0000011110000001",
21398 => "0000011110000010",
21399 => "0000011110000010",
21400 => "0000011110000011",
21401 => "0000011110000011",
21402 => "0000011110000011",
21403 => "0000011110000100",
21404 => "0000011110000100",
21405 => "0000011110000101",
21406 => "0000011110000101",
21407 => "0000011110000110",
21408 => "0000011110000110",
21409 => "0000011110000111",
21410 => "0000011110000111",
21411 => "0000011110000111",
21412 => "0000011110001000",
21413 => "0000011110001000",
21414 => "0000011110001001",
21415 => "0000011110001001",
21416 => "0000011110001010",
21417 => "0000011110001010",
21418 => "0000011110001011",
21419 => "0000011110001011",
21420 => "0000011110001011",
21421 => "0000011110001100",
21422 => "0000011110001100",
21423 => "0000011110001101",
21424 => "0000011110001101",
21425 => "0000011110001110",
21426 => "0000011110001110",
21427 => "0000011110001111",
21428 => "0000011110001111",
21429 => "0000011110001111",
21430 => "0000011110010000",
21431 => "0000011110010000",
21432 => "0000011110010001",
21433 => "0000011110010001",
21434 => "0000011110010010",
21435 => "0000011110010010",
21436 => "0000011110010011",
21437 => "0000011110010011",
21438 => "0000011110010011",
21439 => "0000011110010100",
21440 => "0000011110010100",
21441 => "0000011110010101",
21442 => "0000011110010101",
21443 => "0000011110010110",
21444 => "0000011110010110",
21445 => "0000011110010111",
21446 => "0000011110010111",
21447 => "0000011110010111",
21448 => "0000011110011000",
21449 => "0000011110011000",
21450 => "0000011110011001",
21451 => "0000011110011001",
21452 => "0000011110011010",
21453 => "0000011110011010",
21454 => "0000011110011011",
21455 => "0000011110011011",
21456 => "0000011110011011",
21457 => "0000011110011100",
21458 => "0000011110011100",
21459 => "0000011110011101",
21460 => "0000011110011101",
21461 => "0000011110011110",
21462 => "0000011110011110",
21463 => "0000011110011111",
21464 => "0000011110011111",
21465 => "0000011110100000",
21466 => "0000011110100000",
21467 => "0000011110100000",
21468 => "0000011110100001",
21469 => "0000011110100001",
21470 => "0000011110100010",
21471 => "0000011110100010",
21472 => "0000011110100011",
21473 => "0000011110100011",
21474 => "0000011110100100",
21475 => "0000011110100100",
21476 => "0000011110100100",
21477 => "0000011110100101",
21478 => "0000011110100101",
21479 => "0000011110100110",
21480 => "0000011110100110",
21481 => "0000011110100111",
21482 => "0000011110100111",
21483 => "0000011110101000",
21484 => "0000011110101000",
21485 => "0000011110101000",
21486 => "0000011110101001",
21487 => "0000011110101001",
21488 => "0000011110101010",
21489 => "0000011110101010",
21490 => "0000011110101011",
21491 => "0000011110101011",
21492 => "0000011110101100",
21493 => "0000011110101100",
21494 => "0000011110101101",
21495 => "0000011110101101",
21496 => "0000011110101101",
21497 => "0000011110101110",
21498 => "0000011110101110",
21499 => "0000011110101111",
21500 => "0000011110101111",
21501 => "0000011110110000",
21502 => "0000011110110000",
21503 => "0000011110110001",
21504 => "0000011110110001",
21505 => "0000011110110010",
21506 => "0000011110110010",
21507 => "0000011110110010",
21508 => "0000011110110011",
21509 => "0000011110110011",
21510 => "0000011110110100",
21511 => "0000011110110100",
21512 => "0000011110110101",
21513 => "0000011110110101",
21514 => "0000011110110110",
21515 => "0000011110110110",
21516 => "0000011110110110",
21517 => "0000011110110111",
21518 => "0000011110110111",
21519 => "0000011110111000",
21520 => "0000011110111000",
21521 => "0000011110111001",
21522 => "0000011110111001",
21523 => "0000011110111010",
21524 => "0000011110111010",
21525 => "0000011110111011",
21526 => "0000011110111011",
21527 => "0000011110111011",
21528 => "0000011110111100",
21529 => "0000011110111100",
21530 => "0000011110111101",
21531 => "0000011110111101",
21532 => "0000011110111110",
21533 => "0000011110111110",
21534 => "0000011110111111",
21535 => "0000011110111111",
21536 => "0000011111000000",
21537 => "0000011111000000",
21538 => "0000011111000000",
21539 => "0000011111000001",
21540 => "0000011111000001",
21541 => "0000011111000010",
21542 => "0000011111000010",
21543 => "0000011111000011",
21544 => "0000011111000011",
21545 => "0000011111000100",
21546 => "0000011111000100",
21547 => "0000011111000101",
21548 => "0000011111000101",
21549 => "0000011111000101",
21550 => "0000011111000110",
21551 => "0000011111000110",
21552 => "0000011111000111",
21553 => "0000011111000111",
21554 => "0000011111001000",
21555 => "0000011111001000",
21556 => "0000011111001001",
21557 => "0000011111001001",
21558 => "0000011111001010",
21559 => "0000011111001010",
21560 => "0000011111001011",
21561 => "0000011111001011",
21562 => "0000011111001011",
21563 => "0000011111001100",
21564 => "0000011111001100",
21565 => "0000011111001101",
21566 => "0000011111001101",
21567 => "0000011111001110",
21568 => "0000011111001110",
21569 => "0000011111001111",
21570 => "0000011111001111",
21571 => "0000011111010000",
21572 => "0000011111010000",
21573 => "0000011111010000",
21574 => "0000011111010001",
21575 => "0000011111010001",
21576 => "0000011111010010",
21577 => "0000011111010010",
21578 => "0000011111010011",
21579 => "0000011111010011",
21580 => "0000011111010100",
21581 => "0000011111010100",
21582 => "0000011111010101",
21583 => "0000011111010101",
21584 => "0000011111010110",
21585 => "0000011111010110",
21586 => "0000011111010110",
21587 => "0000011111010111",
21588 => "0000011111010111",
21589 => "0000011111011000",
21590 => "0000011111011000",
21591 => "0000011111011001",
21592 => "0000011111011001",
21593 => "0000011111011010",
21594 => "0000011111011010",
21595 => "0000011111011011",
21596 => "0000011111011011",
21597 => "0000011111011100",
21598 => "0000011111011100",
21599 => "0000011111011100",
21600 => "0000011111011101",
21601 => "0000011111011101",
21602 => "0000011111011110",
21603 => "0000011111011110",
21604 => "0000011111011111",
21605 => "0000011111011111",
21606 => "0000011111100000",
21607 => "0000011111100000",
21608 => "0000011111100001",
21609 => "0000011111100001",
21610 => "0000011111100010",
21611 => "0000011111100010",
21612 => "0000011111100010",
21613 => "0000011111100011",
21614 => "0000011111100011",
21615 => "0000011111100100",
21616 => "0000011111100100",
21617 => "0000011111100101",
21618 => "0000011111100101",
21619 => "0000011111100110",
21620 => "0000011111100110",
21621 => "0000011111100111",
21622 => "0000011111100111",
21623 => "0000011111101000",
21624 => "0000011111101000",
21625 => "0000011111101000",
21626 => "0000011111101001",
21627 => "0000011111101001",
21628 => "0000011111101010",
21629 => "0000011111101010",
21630 => "0000011111101011",
21631 => "0000011111101011",
21632 => "0000011111101100",
21633 => "0000011111101100",
21634 => "0000011111101101",
21635 => "0000011111101101",
21636 => "0000011111101110",
21637 => "0000011111101110",
21638 => "0000011111101110",
21639 => "0000011111101111",
21640 => "0000011111101111",
21641 => "0000011111110000",
21642 => "0000011111110000",
21643 => "0000011111110001",
21644 => "0000011111110001",
21645 => "0000011111110010",
21646 => "0000011111110010",
21647 => "0000011111110011",
21648 => "0000011111110011",
21649 => "0000011111110100",
21650 => "0000011111110100",
21651 => "0000011111110101",
21652 => "0000011111110101",
21653 => "0000011111110101",
21654 => "0000011111110110",
21655 => "0000011111110110",
21656 => "0000011111110111",
21657 => "0000011111110111",
21658 => "0000011111111000",
21659 => "0000011111111000",
21660 => "0000011111111001",
21661 => "0000011111111001",
21662 => "0000011111111010",
21663 => "0000011111111010",
21664 => "0000011111111011",
21665 => "0000011111111011",
21666 => "0000011111111100",
21667 => "0000011111111100",
21668 => "0000011111111100",
21669 => "0000011111111101",
21670 => "0000011111111101",
21671 => "0000011111111110",
21672 => "0000011111111110",
21673 => "0000011111111111",
21674 => "0000011111111111",
21675 => "0000100000000000",
21676 => "0000100000000000",
21677 => "0000100000000000",
21678 => "0000100000000010",
21679 => "0000100000000010",
21680 => "0000100000000010",
21681 => "0000100000000010",
21682 => "0000100000000100",
21683 => "0000100000000100",
21684 => "0000100000000100",
21685 => "0000100000000100",
21686 => "0000100000000100",
21687 => "0000100000000110",
21688 => "0000100000000110",
21689 => "0000100000000110",
21690 => "0000100000000110",
21691 => "0000100000001000",
21692 => "0000100000001000",
21693 => "0000100000001000",
21694 => "0000100000001000",
21695 => "0000100000001010",
21696 => "0000100000001010",
21697 => "0000100000001010",
21698 => "0000100000001010",
21699 => "0000100000001100",
21700 => "0000100000001100",
21701 => "0000100000001100",
21702 => "0000100000001100",
21703 => "0000100000001100",
21704 => "0000100000001110",
21705 => "0000100000001110",
21706 => "0000100000001110",
21707 => "0000100000001110",
21708 => "0000100000010000",
21709 => "0000100000010000",
21710 => "0000100000010000",
21711 => "0000100000010000",
21712 => "0000100000010010",
21713 => "0000100000010010",
21714 => "0000100000010010",
21715 => "0000100000010010",
21716 => "0000100000010100",
21717 => "0000100000010100",
21718 => "0000100000010100",
21719 => "0000100000010100",
21720 => "0000100000010100",
21721 => "0000100000010110",
21722 => "0000100000010110",
21723 => "0000100000010110",
21724 => "0000100000010110",
21725 => "0000100000011000",
21726 => "0000100000011000",
21727 => "0000100000011000",
21728 => "0000100000011000",
21729 => "0000100000011010",
21730 => "0000100000011010",
21731 => "0000100000011010",
21732 => "0000100000011010",
21733 => "0000100000011100",
21734 => "0000100000011100",
21735 => "0000100000011100",
21736 => "0000100000011100",
21737 => "0000100000011110",
21738 => "0000100000011110",
21739 => "0000100000011110",
21740 => "0000100000011110",
21741 => "0000100000011110",
21742 => "0000100000100000",
21743 => "0000100000100000",
21744 => "0000100000100000",
21745 => "0000100000100000",
21746 => "0000100000100010",
21747 => "0000100000100010",
21748 => "0000100000100010",
21749 => "0000100000100010",
21750 => "0000100000100100",
21751 => "0000100000100100",
21752 => "0000100000100100",
21753 => "0000100000100100",
21754 => "0000100000100110",
21755 => "0000100000100110",
21756 => "0000100000100110",
21757 => "0000100000100110",
21758 => "0000100000101000",
21759 => "0000100000101000",
21760 => "0000100000101000",
21761 => "0000100000101000",
21762 => "0000100000101000",
21763 => "0000100000101010",
21764 => "0000100000101010",
21765 => "0000100000101010",
21766 => "0000100000101010",
21767 => "0000100000101100",
21768 => "0000100000101100",
21769 => "0000100000101100",
21770 => "0000100000101100",
21771 => "0000100000101110",
21772 => "0000100000101110",
21773 => "0000100000101110",
21774 => "0000100000101110",
21775 => "0000100000110000",
21776 => "0000100000110000",
21777 => "0000100000110000",
21778 => "0000100000110000",
21779 => "0000100000110010",
21780 => "0000100000110010",
21781 => "0000100000110010",
21782 => "0000100000110010",
21783 => "0000100000110010",
21784 => "0000100000110100",
21785 => "0000100000110100",
21786 => "0000100000110100",
21787 => "0000100000110100",
21788 => "0000100000110110",
21789 => "0000100000110110",
21790 => "0000100000110110",
21791 => "0000100000110110",
21792 => "0000100000111000",
21793 => "0000100000111000",
21794 => "0000100000111000",
21795 => "0000100000111000",
21796 => "0000100000111010",
21797 => "0000100000111010",
21798 => "0000100000111010",
21799 => "0000100000111010",
21800 => "0000100000111100",
21801 => "0000100000111100",
21802 => "0000100000111100",
21803 => "0000100000111100",
21804 => "0000100000111110",
21805 => "0000100000111110",
21806 => "0000100000111110",
21807 => "0000100000111110",
21808 => "0000100000111110",
21809 => "0000100001000000",
21810 => "0000100001000000",
21811 => "0000100001000000",
21812 => "0000100001000000",
21813 => "0000100001000010",
21814 => "0000100001000010",
21815 => "0000100001000010",
21816 => "0000100001000010",
21817 => "0000100001000100",
21818 => "0000100001000100",
21819 => "0000100001000100",
21820 => "0000100001000100",
21821 => "0000100001000110",
21822 => "0000100001000110",
21823 => "0000100001000110",
21824 => "0000100001000110",
21825 => "0000100001001000",
21826 => "0000100001001000",
21827 => "0000100001001000",
21828 => "0000100001001000",
21829 => "0000100001001010",
21830 => "0000100001001010",
21831 => "0000100001001010",
21832 => "0000100001001010",
21833 => "0000100001001100",
21834 => "0000100001001100",
21835 => "0000100001001100",
21836 => "0000100001001100",
21837 => "0000100001001110",
21838 => "0000100001001110",
21839 => "0000100001001110",
21840 => "0000100001001110",
21841 => "0000100001001110",
21842 => "0000100001010000",
21843 => "0000100001010000",
21844 => "0000100001010000",
21845 => "0000100001010000",
21846 => "0000100001010010",
21847 => "0000100001010010",
21848 => "0000100001010010",
21849 => "0000100001010010",
21850 => "0000100001010100",
21851 => "0000100001010100",
21852 => "0000100001010100",
21853 => "0000100001010100",
21854 => "0000100001010110",
21855 => "0000100001010110",
21856 => "0000100001010110",
21857 => "0000100001010110",
21858 => "0000100001011000",
21859 => "0000100001011000",
21860 => "0000100001011000",
21861 => "0000100001011000",
21862 => "0000100001011010",
21863 => "0000100001011010",
21864 => "0000100001011010",
21865 => "0000100001011010",
21866 => "0000100001011100",
21867 => "0000100001011100",
21868 => "0000100001011100",
21869 => "0000100001011100",
21870 => "0000100001011110",
21871 => "0000100001011110",
21872 => "0000100001011110",
21873 => "0000100001011110",
21874 => "0000100001100000",
21875 => "0000100001100000",
21876 => "0000100001100000",
21877 => "0000100001100000",
21878 => "0000100001100010",
21879 => "0000100001100010",
21880 => "0000100001100010",
21881 => "0000100001100010",
21882 => "0000100001100010",
21883 => "0000100001100100",
21884 => "0000100001100100",
21885 => "0000100001100100",
21886 => "0000100001100100",
21887 => "0000100001100110",
21888 => "0000100001100110",
21889 => "0000100001100110",
21890 => "0000100001100110",
21891 => "0000100001101000",
21892 => "0000100001101000",
21893 => "0000100001101000",
21894 => "0000100001101000",
21895 => "0000100001101010",
21896 => "0000100001101010",
21897 => "0000100001101010",
21898 => "0000100001101010",
21899 => "0000100001101100",
21900 => "0000100001101100",
21901 => "0000100001101100",
21902 => "0000100001101100",
21903 => "0000100001101110",
21904 => "0000100001101110",
21905 => "0000100001101110",
21906 => "0000100001101110",
21907 => "0000100001110000",
21908 => "0000100001110000",
21909 => "0000100001110000",
21910 => "0000100001110000",
21911 => "0000100001110010",
21912 => "0000100001110010",
21913 => "0000100001110010",
21914 => "0000100001110010",
21915 => "0000100001110100",
21916 => "0000100001110100",
21917 => "0000100001110100",
21918 => "0000100001110100",
21919 => "0000100001110110",
21920 => "0000100001110110",
21921 => "0000100001110110",
21922 => "0000100001110110",
21923 => "0000100001111000",
21924 => "0000100001111000",
21925 => "0000100001111000",
21926 => "0000100001111000",
21927 => "0000100001111010",
21928 => "0000100001111010",
21929 => "0000100001111010",
21930 => "0000100001111010",
21931 => "0000100001111100",
21932 => "0000100001111100",
21933 => "0000100001111100",
21934 => "0000100001111100",
21935 => "0000100001111110",
21936 => "0000100001111110",
21937 => "0000100001111110",
21938 => "0000100001111110",
21939 => "0000100010000000",
21940 => "0000100010000000",
21941 => "0000100010000000",
21942 => "0000100010000000",
21943 => "0000100010000010",
21944 => "0000100010000010",
21945 => "0000100010000010",
21946 => "0000100010000010",
21947 => "0000100010000100",
21948 => "0000100010000100",
21949 => "0000100010000100",
21950 => "0000100010000100",
21951 => "0000100010000110",
21952 => "0000100010000110",
21953 => "0000100010000110",
21954 => "0000100010000110",
21955 => "0000100010000110",
21956 => "0000100010001000",
21957 => "0000100010001000",
21958 => "0000100010001000",
21959 => "0000100010001000",
21960 => "0000100010001010",
21961 => "0000100010001010",
21962 => "0000100010001010",
21963 => "0000100010001010",
21964 => "0000100010001100",
21965 => "0000100010001100",
21966 => "0000100010001100",
21967 => "0000100010001100",
21968 => "0000100010001110",
21969 => "0000100010001110",
21970 => "0000100010001110",
21971 => "0000100010001110",
21972 => "0000100010010000",
21973 => "0000100010010000",
21974 => "0000100010010000",
21975 => "0000100010010000",
21976 => "0000100010010010",
21977 => "0000100010010010",
21978 => "0000100010010010",
21979 => "0000100010010010",
21980 => "0000100010010100",
21981 => "0000100010010100",
21982 => "0000100010010100",
21983 => "0000100010010100",
21984 => "0000100010010110",
21985 => "0000100010010110",
21986 => "0000100010010110",
21987 => "0000100010010110",
21988 => "0000100010011000",
21989 => "0000100010011000",
21990 => "0000100010011000",
21991 => "0000100010011000",
21992 => "0000100010011010",
21993 => "0000100010011010",
21994 => "0000100010011010",
21995 => "0000100010011010",
21996 => "0000100010011100",
21997 => "0000100010011100",
21998 => "0000100010011100",
21999 => "0000100010011100",
22000 => "0000100010011110",
22001 => "0000100010011110",
22002 => "0000100010011110",
22003 => "0000100010011110",
22004 => "0000100010100000",
22005 => "0000100010100000",
22006 => "0000100010100000",
22007 => "0000100010100010",
22008 => "0000100010100010",
22009 => "0000100010100010",
22010 => "0000100010100010",
22011 => "0000100010100100",
22012 => "0000100010100100",
22013 => "0000100010100100",
22014 => "0000100010100100",
22015 => "0000100010100110",
22016 => "0000100010100110",
22017 => "0000100010100110",
22018 => "0000100010100110",
22019 => "0000100010101000",
22020 => "0000100010101000",
22021 => "0000100010101000",
22022 => "0000100010101000",
22023 => "0000100010101010",
22024 => "0000100010101010",
22025 => "0000100010101010",
22026 => "0000100010101010",
22027 => "0000100010101100",
22028 => "0000100010101100",
22029 => "0000100010101100",
22030 => "0000100010101100",
22031 => "0000100010101110",
22032 => "0000100010101110",
22033 => "0000100010101110",
22034 => "0000100010101110",
22035 => "0000100010110000",
22036 => "0000100010110000",
22037 => "0000100010110000",
22038 => "0000100010110000",
22039 => "0000100010110010",
22040 => "0000100010110010",
22041 => "0000100010110010",
22042 => "0000100010110010",
22043 => "0000100010110100",
22044 => "0000100010110100",
22045 => "0000100010110100",
22046 => "0000100010110100",
22047 => "0000100010110110",
22048 => "0000100010110110",
22049 => "0000100010110110",
22050 => "0000100010110110",
22051 => "0000100010111000",
22052 => "0000100010111000",
22053 => "0000100010111000",
22054 => "0000100010111000",
22055 => "0000100010111010",
22056 => "0000100010111010",
22057 => "0000100010111010",
22058 => "0000100010111010",
22059 => "0000100010111100",
22060 => "0000100010111100",
22061 => "0000100010111100",
22062 => "0000100010111100",
22063 => "0000100010111110",
22064 => "0000100010111110",
22065 => "0000100010111110",
22066 => "0000100010111110",
22067 => "0000100011000000",
22068 => "0000100011000000",
22069 => "0000100011000000",
22070 => "0000100011000000",
22071 => "0000100011000010",
22072 => "0000100011000010",
22073 => "0000100011000010",
22074 => "0000100011000010",
22075 => "0000100011000100",
22076 => "0000100011000100",
22077 => "0000100011000100",
22078 => "0000100011000100",
22079 => "0000100011000110",
22080 => "0000100011000110",
22081 => "0000100011000110",
22082 => "0000100011001000",
22083 => "0000100011001000",
22084 => "0000100011001000",
22085 => "0000100011001000",
22086 => "0000100011001010",
22087 => "0000100011001010",
22088 => "0000100011001010",
22089 => "0000100011001010",
22090 => "0000100011001100",
22091 => "0000100011001100",
22092 => "0000100011001100",
22093 => "0000100011001100",
22094 => "0000100011001110",
22095 => "0000100011001110",
22096 => "0000100011001110",
22097 => "0000100011001110",
22098 => "0000100011010000",
22099 => "0000100011010000",
22100 => "0000100011010000",
22101 => "0000100011010000",
22102 => "0000100011010010",
22103 => "0000100011010010",
22104 => "0000100011010010",
22105 => "0000100011010010",
22106 => "0000100011010100",
22107 => "0000100011010100",
22108 => "0000100011010100",
22109 => "0000100011010100",
22110 => "0000100011010110",
22111 => "0000100011010110",
22112 => "0000100011010110",
22113 => "0000100011010110",
22114 => "0000100011011000",
22115 => "0000100011011000",
22116 => "0000100011011000",
22117 => "0000100011011000",
22118 => "0000100011011010",
22119 => "0000100011011010",
22120 => "0000100011011010",
22121 => "0000100011011100",
22122 => "0000100011011100",
22123 => "0000100011011100",
22124 => "0000100011011100",
22125 => "0000100011011110",
22126 => "0000100011011110",
22127 => "0000100011011110",
22128 => "0000100011011110",
22129 => "0000100011100000",
22130 => "0000100011100000",
22131 => "0000100011100000",
22132 => "0000100011100000",
22133 => "0000100011100010",
22134 => "0000100011100010",
22135 => "0000100011100010",
22136 => "0000100011100010",
22137 => "0000100011100100",
22138 => "0000100011100100",
22139 => "0000100011100100",
22140 => "0000100011100100",
22141 => "0000100011100110",
22142 => "0000100011100110",
22143 => "0000100011100110",
22144 => "0000100011100110",
22145 => "0000100011101000",
22146 => "0000100011101000",
22147 => "0000100011101000",
22148 => "0000100011101000",
22149 => "0000100011101010",
22150 => "0000100011101010",
22151 => "0000100011101010",
22152 => "0000100011101100",
22153 => "0000100011101100",
22154 => "0000100011101100",
22155 => "0000100011101100",
22156 => "0000100011101110",
22157 => "0000100011101110",
22158 => "0000100011101110",
22159 => "0000100011101110",
22160 => "0000100011110000",
22161 => "0000100011110000",
22162 => "0000100011110000",
22163 => "0000100011110000",
22164 => "0000100011110010",
22165 => "0000100011110010",
22166 => "0000100011110010",
22167 => "0000100011110010",
22168 => "0000100011110100",
22169 => "0000100011110100",
22170 => "0000100011110100",
22171 => "0000100011110100",
22172 => "0000100011110110",
22173 => "0000100011110110",
22174 => "0000100011110110",
22175 => "0000100011111000",
22176 => "0000100011111000",
22177 => "0000100011111000",
22178 => "0000100011111000",
22179 => "0000100011111010",
22180 => "0000100011111010",
22181 => "0000100011111010",
22182 => "0000100011111010",
22183 => "0000100011111100",
22184 => "0000100011111100",
22185 => "0000100011111100",
22186 => "0000100011111100",
22187 => "0000100011111110",
22188 => "0000100011111110",
22189 => "0000100011111110",
22190 => "0000100011111110",
22191 => "0000100100000000",
22192 => "0000100100000000",
22193 => "0000100100000000",
22194 => "0000100100000000",
22195 => "0000100100000010",
22196 => "0000100100000010",
22197 => "0000100100000010",
22198 => "0000100100000100",
22199 => "0000100100000100",
22200 => "0000100100000100",
22201 => "0000100100000100",
22202 => "0000100100000110",
22203 => "0000100100000110",
22204 => "0000100100000110",
22205 => "0000100100000110",
22206 => "0000100100001000",
22207 => "0000100100001000",
22208 => "0000100100001000",
22209 => "0000100100001000",
22210 => "0000100100001010",
22211 => "0000100100001010",
22212 => "0000100100001010",
22213 => "0000100100001010",
22214 => "0000100100001100",
22215 => "0000100100001100",
22216 => "0000100100001100",
22217 => "0000100100001110",
22218 => "0000100100001110",
22219 => "0000100100001110",
22220 => "0000100100001110",
22221 => "0000100100010000",
22222 => "0000100100010000",
22223 => "0000100100010000",
22224 => "0000100100010000",
22225 => "0000100100010010",
22226 => "0000100100010010",
22227 => "0000100100010010",
22228 => "0000100100010010",
22229 => "0000100100010100",
22230 => "0000100100010100",
22231 => "0000100100010100",
22232 => "0000100100010100",
22233 => "0000100100010110",
22234 => "0000100100010110",
22235 => "0000100100010110",
22236 => "0000100100011000",
22237 => "0000100100011000",
22238 => "0000100100011000",
22239 => "0000100100011000",
22240 => "0000100100011010",
22241 => "0000100100011010",
22242 => "0000100100011010",
22243 => "0000100100011010",
22244 => "0000100100011100",
22245 => "0000100100011100",
22246 => "0000100100011100",
22247 => "0000100100011100",
22248 => "0000100100011110",
22249 => "0000100100011110",
22250 => "0000100100011110",
22251 => "0000100100011110",
22252 => "0000100100100000",
22253 => "0000100100100000",
22254 => "0000100100100000",
22255 => "0000100100100010",
22256 => "0000100100100010",
22257 => "0000100100100010",
22258 => "0000100100100010",
22259 => "0000100100100100",
22260 => "0000100100100100",
22261 => "0000100100100100",
22262 => "0000100100100100",
22263 => "0000100100100110",
22264 => "0000100100100110",
22265 => "0000100100100110",
22266 => "0000100100100110",
22267 => "0000100100101000",
22268 => "0000100100101000",
22269 => "0000100100101000",
22270 => "0000100100101010",
22271 => "0000100100101010",
22272 => "0000100100101010",
22273 => "0000100100101010",
22274 => "0000100100101100",
22275 => "0000100100101100",
22276 => "0000100100101100",
22277 => "0000100100101100",
22278 => "0000100100101110",
22279 => "0000100100101110",
22280 => "0000100100101110",
22281 => "0000100100101110",
22282 => "0000100100110000",
22283 => "0000100100110000",
22284 => "0000100100110000",
22285 => "0000100100110010",
22286 => "0000100100110010",
22287 => "0000100100110010",
22288 => "0000100100110010",
22289 => "0000100100110100",
22290 => "0000100100110100",
22291 => "0000100100110100",
22292 => "0000100100110100",
22293 => "0000100100110110",
22294 => "0000100100110110",
22295 => "0000100100110110",
22296 => "0000100100110110",
22297 => "0000100100111000",
22298 => "0000100100111000",
22299 => "0000100100111000",
22300 => "0000100100111010",
22301 => "0000100100111010",
22302 => "0000100100111010",
22303 => "0000100100111010",
22304 => "0000100100111100",
22305 => "0000100100111100",
22306 => "0000100100111100",
22307 => "0000100100111100",
22308 => "0000100100111110",
22309 => "0000100100111110",
22310 => "0000100100111110",
22311 => "0000100100111110",
22312 => "0000100101000000",
22313 => "0000100101000000",
22314 => "0000100101000000",
22315 => "0000100101000010",
22316 => "0000100101000010",
22317 => "0000100101000010",
22318 => "0000100101000010",
22319 => "0000100101000100",
22320 => "0000100101000100",
22321 => "0000100101000100",
22322 => "0000100101000100",
22323 => "0000100101000110",
22324 => "0000100101000110",
22325 => "0000100101000110",
22326 => "0000100101000110",
22327 => "0000100101001000",
22328 => "0000100101001000",
22329 => "0000100101001000",
22330 => "0000100101001010",
22331 => "0000100101001010",
22332 => "0000100101001010",
22333 => "0000100101001010",
22334 => "0000100101001100",
22335 => "0000100101001100",
22336 => "0000100101001100",
22337 => "0000100101001100",
22338 => "0000100101001110",
22339 => "0000100101001110",
22340 => "0000100101001110",
22341 => "0000100101010000",
22342 => "0000100101010000",
22343 => "0000100101010000",
22344 => "0000100101010000",
22345 => "0000100101010010",
22346 => "0000100101010010",
22347 => "0000100101010010",
22348 => "0000100101010010",
22349 => "0000100101010100",
22350 => "0000100101010100",
22351 => "0000100101010100",
22352 => "0000100101010100",
22353 => "0000100101010110",
22354 => "0000100101010110",
22355 => "0000100101010110",
22356 => "0000100101011000",
22357 => "0000100101011000",
22358 => "0000100101011000",
22359 => "0000100101011000",
22360 => "0000100101011010",
22361 => "0000100101011010",
22362 => "0000100101011010",
22363 => "0000100101011010",
22364 => "0000100101011100",
22365 => "0000100101011100",
22366 => "0000100101011100",
22367 => "0000100101011110",
22368 => "0000100101011110",
22369 => "0000100101011110",
22370 => "0000100101011110",
22371 => "0000100101100000",
22372 => "0000100101100000",
22373 => "0000100101100000",
22374 => "0000100101100000",
22375 => "0000100101100010",
22376 => "0000100101100010",
22377 => "0000100101100010",
22378 => "0000100101100100",
22379 => "0000100101100100",
22380 => "0000100101100100",
22381 => "0000100101100100",
22382 => "0000100101100110",
22383 => "0000100101100110",
22384 => "0000100101100110",
22385 => "0000100101100110",
22386 => "0000100101101000",
22387 => "0000100101101000",
22388 => "0000100101101000",
22389 => "0000100101101010",
22390 => "0000100101101010",
22391 => "0000100101101010",
22392 => "0000100101101010",
22393 => "0000100101101100",
22394 => "0000100101101100",
22395 => "0000100101101100",
22396 => "0000100101101100",
22397 => "0000100101101110",
22398 => "0000100101101110",
22399 => "0000100101101110",
22400 => "0000100101110000",
22401 => "0000100101110000",
22402 => "0000100101110000",
22403 => "0000100101110000",
22404 => "0000100101110010",
22405 => "0000100101110010",
22406 => "0000100101110010",
22407 => "0000100101110010",
22408 => "0000100101110100",
22409 => "0000100101110100",
22410 => "0000100101110100",
22411 => "0000100101110110",
22412 => "0000100101110110",
22413 => "0000100101110110",
22414 => "0000100101110110",
22415 => "0000100101111000",
22416 => "0000100101111000",
22417 => "0000100101111000",
22418 => "0000100101111000",
22419 => "0000100101111010",
22420 => "0000100101111010",
22421 => "0000100101111010",
22422 => "0000100101111100",
22423 => "0000100101111100",
22424 => "0000100101111100",
22425 => "0000100101111100",
22426 => "0000100101111110",
22427 => "0000100101111110",
22428 => "0000100101111110",
22429 => "0000100101111110",
22430 => "0000100110000000",
22431 => "0000100110000000",
22432 => "0000100110000000",
22433 => "0000100110000010",
22434 => "0000100110000010",
22435 => "0000100110000010",
22436 => "0000100110000010",
22437 => "0000100110000100",
22438 => "0000100110000100",
22439 => "0000100110000100",
22440 => "0000100110000110",
22441 => "0000100110000110",
22442 => "0000100110000110",
22443 => "0000100110000110",
22444 => "0000100110001000",
22445 => "0000100110001000",
22446 => "0000100110001000",
22447 => "0000100110001000",
22448 => "0000100110001010",
22449 => "0000100110001010",
22450 => "0000100110001010",
22451 => "0000100110001100",
22452 => "0000100110001100",
22453 => "0000100110001100",
22454 => "0000100110001100",
22455 => "0000100110001110",
22456 => "0000100110001110",
22457 => "0000100110001110",
22458 => "0000100110001110",
22459 => "0000100110010000",
22460 => "0000100110010000",
22461 => "0000100110010000",
22462 => "0000100110010010",
22463 => "0000100110010010",
22464 => "0000100110010010",
22465 => "0000100110010010",
22466 => "0000100110010100",
22467 => "0000100110010100",
22468 => "0000100110010100",
22469 => "0000100110010110",
22470 => "0000100110010110",
22471 => "0000100110010110",
22472 => "0000100110010110",
22473 => "0000100110011000",
22474 => "0000100110011000",
22475 => "0000100110011000",
22476 => "0000100110011000",
22477 => "0000100110011010",
22478 => "0000100110011010",
22479 => "0000100110011010",
22480 => "0000100110011100",
22481 => "0000100110011100",
22482 => "0000100110011100",
22483 => "0000100110011100",
22484 => "0000100110011110",
22485 => "0000100110011110",
22486 => "0000100110011110",
22487 => "0000100110100000",
22488 => "0000100110100000",
22489 => "0000100110100000",
22490 => "0000100110100000",
22491 => "0000100110100010",
22492 => "0000100110100010",
22493 => "0000100110100010",
22494 => "0000100110100010",
22495 => "0000100110100100",
22496 => "0000100110100100",
22497 => "0000100110100100",
22498 => "0000100110100110",
22499 => "0000100110100110",
22500 => "0000100110100110",
22501 => "0000100110100110",
22502 => "0000100110101000",
22503 => "0000100110101000",
22504 => "0000100110101000",
22505 => "0000100110101010",
22506 => "0000100110101010",
22507 => "0000100110101010",
22508 => "0000100110101010",
22509 => "0000100110101100",
22510 => "0000100110101100",
22511 => "0000100110101100",
22512 => "0000100110101100",
22513 => "0000100110101110",
22514 => "0000100110101110",
22515 => "0000100110101110",
22516 => "0000100110110000",
22517 => "0000100110110000",
22518 => "0000100110110000",
22519 => "0000100110110000",
22520 => "0000100110110010",
22521 => "0000100110110010",
22522 => "0000100110110010",
22523 => "0000100110110100",
22524 => "0000100110110100",
22525 => "0000100110110100",
22526 => "0000100110110100",
22527 => "0000100110110110",
22528 => "0000100110110110",
22529 => "0000100110110110",
22530 => "0000100110111000",
22531 => "0000100110111000",
22532 => "0000100110111000",
22533 => "0000100110111000",
22534 => "0000100110111010",
22535 => "0000100110111010",
22536 => "0000100110111010",
22537 => "0000100110111010",
22538 => "0000100110111100",
22539 => "0000100110111100",
22540 => "0000100110111100",
22541 => "0000100110111110",
22542 => "0000100110111110",
22543 => "0000100110111110",
22544 => "0000100110111110",
22545 => "0000100111000000",
22546 => "0000100111000000",
22547 => "0000100111000000",
22548 => "0000100111000010",
22549 => "0000100111000010",
22550 => "0000100111000010",
22551 => "0000100111000010",
22552 => "0000100111000100",
22553 => "0000100111000100",
22554 => "0000100111000100",
22555 => "0000100111000110",
22556 => "0000100111000110",
22557 => "0000100111000110",
22558 => "0000100111000110",
22559 => "0000100111001000",
22560 => "0000100111001000",
22561 => "0000100111001000",
22562 => "0000100111001010",
22563 => "0000100111001010",
22564 => "0000100111001010",
22565 => "0000100111001010",
22566 => "0000100111001100",
22567 => "0000100111001100",
22568 => "0000100111001100",
22569 => "0000100111001110",
22570 => "0000100111001110",
22571 => "0000100111001110",
22572 => "0000100111001110",
22573 => "0000100111010000",
22574 => "0000100111010000",
22575 => "0000100111010000",
22576 => "0000100111010000",
22577 => "0000100111010010",
22578 => "0000100111010010",
22579 => "0000100111010010",
22580 => "0000100111010100",
22581 => "0000100111010100",
22582 => "0000100111010100",
22583 => "0000100111010100",
22584 => "0000100111010110",
22585 => "0000100111010110",
22586 => "0000100111010110",
22587 => "0000100111011000",
22588 => "0000100111011000",
22589 => "0000100111011000",
22590 => "0000100111011000",
22591 => "0000100111011010",
22592 => "0000100111011010",
22593 => "0000100111011010",
22594 => "0000100111011100",
22595 => "0000100111011100",
22596 => "0000100111011100",
22597 => "0000100111011100",
22598 => "0000100111011110",
22599 => "0000100111011110",
22600 => "0000100111011110",
22601 => "0000100111100000",
22602 => "0000100111100000",
22603 => "0000100111100000",
22604 => "0000100111100000",
22605 => "0000100111100010",
22606 => "0000100111100010",
22607 => "0000100111100010",
22608 => "0000100111100100",
22609 => "0000100111100100",
22610 => "0000100111100100",
22611 => "0000100111100100",
22612 => "0000100111100110",
22613 => "0000100111100110",
22614 => "0000100111100110",
22615 => "0000100111101000",
22616 => "0000100111101000",
22617 => "0000100111101000",
22618 => "0000100111101000",
22619 => "0000100111101010",
22620 => "0000100111101010",
22621 => "0000100111101010",
22622 => "0000100111101100",
22623 => "0000100111101100",
22624 => "0000100111101100",
22625 => "0000100111101100",
22626 => "0000100111101110",
22627 => "0000100111101110",
22628 => "0000100111101110",
22629 => "0000100111110000",
22630 => "0000100111110000",
22631 => "0000100111110000",
22632 => "0000100111110000",
22633 => "0000100111110010",
22634 => "0000100111110010",
22635 => "0000100111110010",
22636 => "0000100111110100",
22637 => "0000100111110100",
22638 => "0000100111110100",
22639 => "0000100111110100",
22640 => "0000100111110110",
22641 => "0000100111110110",
22642 => "0000100111110110",
22643 => "0000100111111000",
22644 => "0000100111111000",
22645 => "0000100111111000",
22646 => "0000100111111000",
22647 => "0000100111111010",
22648 => "0000100111111010",
22649 => "0000100111111010",
22650 => "0000100111111100",
22651 => "0000100111111100",
22652 => "0000100111111100",
22653 => "0000100111111100",
22654 => "0000100111111110",
22655 => "0000100111111110",
22656 => "0000100111111110",
22657 => "0000101000000000",
22658 => "0000101000000000",
22659 => "0000101000000000",
22660 => "0000101000000000",
22661 => "0000101000000010",
22662 => "0000101000000010",
22663 => "0000101000000010",
22664 => "0000101000000100",
22665 => "0000101000000100",
22666 => "0000101000000100",
22667 => "0000101000000110",
22668 => "0000101000000110",
22669 => "0000101000000110",
22670 => "0000101000000110",
22671 => "0000101000001000",
22672 => "0000101000001000",
22673 => "0000101000001000",
22674 => "0000101000001010",
22675 => "0000101000001010",
22676 => "0000101000001010",
22677 => "0000101000001010",
22678 => "0000101000001100",
22679 => "0000101000001100",
22680 => "0000101000001100",
22681 => "0000101000001110",
22682 => "0000101000001110",
22683 => "0000101000001110",
22684 => "0000101000001110",
22685 => "0000101000010000",
22686 => "0000101000010000",
22687 => "0000101000010000",
22688 => "0000101000010010",
22689 => "0000101000010010",
22690 => "0000101000010010",
22691 => "0000101000010010",
22692 => "0000101000010100",
22693 => "0000101000010100",
22694 => "0000101000010100",
22695 => "0000101000010110",
22696 => "0000101000010110",
22697 => "0000101000010110",
22698 => "0000101000010110",
22699 => "0000101000011000",
22700 => "0000101000011000",
22701 => "0000101000011000",
22702 => "0000101000011010",
22703 => "0000101000011010",
22704 => "0000101000011010",
22705 => "0000101000011100",
22706 => "0000101000011100",
22707 => "0000101000011100",
22708 => "0000101000011100",
22709 => "0000101000011110",
22710 => "0000101000011110",
22711 => "0000101000011110",
22712 => "0000101000100000",
22713 => "0000101000100000",
22714 => "0000101000100000",
22715 => "0000101000100000",
22716 => "0000101000100010",
22717 => "0000101000100010",
22718 => "0000101000100010",
22719 => "0000101000100100",
22720 => "0000101000100100",
22721 => "0000101000100100",
22722 => "0000101000100100",
22723 => "0000101000100110",
22724 => "0000101000100110",
22725 => "0000101000100110",
22726 => "0000101000101000",
22727 => "0000101000101000",
22728 => "0000101000101000",
22729 => "0000101000101010",
22730 => "0000101000101010",
22731 => "0000101000101010",
22732 => "0000101000101010",
22733 => "0000101000101100",
22734 => "0000101000101100",
22735 => "0000101000101100",
22736 => "0000101000101110",
22737 => "0000101000101110",
22738 => "0000101000101110",
22739 => "0000101000101110",
22740 => "0000101000110000",
22741 => "0000101000110000",
22742 => "0000101000110000",
22743 => "0000101000110010",
22744 => "0000101000110010",
22745 => "0000101000110010",
22746 => "0000101000110010",
22747 => "0000101000110100",
22748 => "0000101000110100",
22749 => "0000101000110100",
22750 => "0000101000110110",
22751 => "0000101000110110",
22752 => "0000101000110110",
22753 => "0000101000111000",
22754 => "0000101000111000",
22755 => "0000101000111000",
22756 => "0000101000111000",
22757 => "0000101000111010",
22758 => "0000101000111010",
22759 => "0000101000111010",
22760 => "0000101000111100",
22761 => "0000101000111100",
22762 => "0000101000111100",
22763 => "0000101000111100",
22764 => "0000101000111110",
22765 => "0000101000111110",
22766 => "0000101000111110",
22767 => "0000101001000000",
22768 => "0000101001000000",
22769 => "0000101001000000",
22770 => "0000101001000010",
22771 => "0000101001000010",
22772 => "0000101001000010",
22773 => "0000101001000010",
22774 => "0000101001000100",
22775 => "0000101001000100",
22776 => "0000101001000100",
22777 => "0000101001000110",
22778 => "0000101001000110",
22779 => "0000101001000110",
22780 => "0000101001000110",
22781 => "0000101001001000",
22782 => "0000101001001000",
22783 => "0000101001001000",
22784 => "0000101001001010",
22785 => "0000101001001010",
22786 => "0000101001001010",
22787 => "0000101001001100",
22788 => "0000101001001100",
22789 => "0000101001001100",
22790 => "0000101001001100",
22791 => "0000101001001110",
22792 => "0000101001001110",
22793 => "0000101001001110",
22794 => "0000101001010000",
22795 => "0000101001010000",
22796 => "0000101001010000",
22797 => "0000101001010010",
22798 => "0000101001010010",
22799 => "0000101001010010",
22800 => "0000101001010010",
22801 => "0000101001010100",
22802 => "0000101001010100",
22803 => "0000101001010100",
22804 => "0000101001010110",
22805 => "0000101001010110",
22806 => "0000101001010110",
22807 => "0000101001010110",
22808 => "0000101001011000",
22809 => "0000101001011000",
22810 => "0000101001011000",
22811 => "0000101001011010",
22812 => "0000101001011010",
22813 => "0000101001011010",
22814 => "0000101001011100",
22815 => "0000101001011100",
22816 => "0000101001011100",
22817 => "0000101001011100",
22818 => "0000101001011110",
22819 => "0000101001011110",
22820 => "0000101001011110",
22821 => "0000101001100000",
22822 => "0000101001100000",
22823 => "0000101001100000",
22824 => "0000101001100010",
22825 => "0000101001100010",
22826 => "0000101001100010",
22827 => "0000101001100010",
22828 => "0000101001100100",
22829 => "0000101001100100",
22830 => "0000101001100100",
22831 => "0000101001100110",
22832 => "0000101001100110",
22833 => "0000101001100110",
22834 => "0000101001101000",
22835 => "0000101001101000",
22836 => "0000101001101000",
22837 => "0000101001101000",
22838 => "0000101001101010",
22839 => "0000101001101010",
22840 => "0000101001101010",
22841 => "0000101001101100",
22842 => "0000101001101100",
22843 => "0000101001101100",
22844 => "0000101001101110",
22845 => "0000101001101110",
22846 => "0000101001101110",
22847 => "0000101001101110",
22848 => "0000101001110000",
22849 => "0000101001110000",
22850 => "0000101001110000",
22851 => "0000101001110010",
22852 => "0000101001110010",
22853 => "0000101001110010",
22854 => "0000101001110100",
22855 => "0000101001110100",
22856 => "0000101001110100",
22857 => "0000101001110100",
22858 => "0000101001110110",
22859 => "0000101001110110",
22860 => "0000101001110110",
22861 => "0000101001111000",
22862 => "0000101001111000",
22863 => "0000101001111000",
22864 => "0000101001111010",
22865 => "0000101001111010",
22866 => "0000101001111010",
22867 => "0000101001111010",
22868 => "0000101001111100",
22869 => "0000101001111100",
22870 => "0000101001111100",
22871 => "0000101001111110",
22872 => "0000101001111110",
22873 => "0000101001111110",
22874 => "0000101010000000",
22875 => "0000101010000000",
22876 => "0000101010000000",
22877 => "0000101010000000",
22878 => "0000101010000010",
22879 => "0000101010000010",
22880 => "0000101010000010",
22881 => "0000101010000100",
22882 => "0000101010000100",
22883 => "0000101010000100",
22884 => "0000101010000110",
22885 => "0000101010000110",
22886 => "0000101010000110",
22887 => "0000101010000110",
22888 => "0000101010001000",
22889 => "0000101010001000",
22890 => "0000101010001000",
22891 => "0000101010001010",
22892 => "0000101010001010",
22893 => "0000101010001010",
22894 => "0000101010001100",
22895 => "0000101010001100",
22896 => "0000101010001100",
22897 => "0000101010001100",
22898 => "0000101010001110",
22899 => "0000101010001110",
22900 => "0000101010001110",
22901 => "0000101010010000",
22902 => "0000101010010000",
22903 => "0000101010010000",
22904 => "0000101010010010",
22905 => "0000101010010010",
22906 => "0000101010010010",
22907 => "0000101010010100",
22908 => "0000101010010100",
22909 => "0000101010010100",
22910 => "0000101010010100",
22911 => "0000101010010110",
22912 => "0000101010010110",
22913 => "0000101010010110",
22914 => "0000101010011000",
22915 => "0000101010011000",
22916 => "0000101010011000",
22917 => "0000101010011010",
22918 => "0000101010011010",
22919 => "0000101010011010",
22920 => "0000101010011010",
22921 => "0000101010011100",
22922 => "0000101010011100",
22923 => "0000101010011100",
22924 => "0000101010011110",
22925 => "0000101010011110",
22926 => "0000101010011110",
22927 => "0000101010100000",
22928 => "0000101010100000",
22929 => "0000101010100000",
22930 => "0000101010100000",
22931 => "0000101010100010",
22932 => "0000101010100010",
22933 => "0000101010100010",
22934 => "0000101010100100",
22935 => "0000101010100100",
22936 => "0000101010100100",
22937 => "0000101010100110",
22938 => "0000101010100110",
22939 => "0000101010100110",
22940 => "0000101010101000",
22941 => "0000101010101000",
22942 => "0000101010101000",
22943 => "0000101010101000",
22944 => "0000101010101010",
22945 => "0000101010101010",
22946 => "0000101010101010",
22947 => "0000101010101100",
22948 => "0000101010101100",
22949 => "0000101010101100",
22950 => "0000101010101110",
22951 => "0000101010101110",
22952 => "0000101010101110",
22953 => "0000101010110000",
22954 => "0000101010110000",
22955 => "0000101010110000",
22956 => "0000101010110000",
22957 => "0000101010110010",
22958 => "0000101010110010",
22959 => "0000101010110010",
22960 => "0000101010110100",
22961 => "0000101010110100",
22962 => "0000101010110100",
22963 => "0000101010110110",
22964 => "0000101010110110",
22965 => "0000101010110110",
22966 => "0000101010110110",
22967 => "0000101010111000",
22968 => "0000101010111000",
22969 => "0000101010111000",
22970 => "0000101010111010",
22971 => "0000101010111010",
22972 => "0000101010111010",
22973 => "0000101010111100",
22974 => "0000101010111100",
22975 => "0000101010111100",
22976 => "0000101010111110",
22977 => "0000101010111110",
22978 => "0000101010111110",
22979 => "0000101010111110",
22980 => "0000101011000000",
22981 => "0000101011000000",
22982 => "0000101011000000",
22983 => "0000101011000010",
22984 => "0000101011000010",
22985 => "0000101011000010",
22986 => "0000101011000100",
22987 => "0000101011000100",
22988 => "0000101011000100",
22989 => "0000101011000110",
22990 => "0000101011000110",
22991 => "0000101011000110",
22992 => "0000101011000110",
22993 => "0000101011001000",
22994 => "0000101011001000",
22995 => "0000101011001000",
22996 => "0000101011001010",
22997 => "0000101011001010",
22998 => "0000101011001010",
22999 => "0000101011001100",
23000 => "0000101011001100",
23001 => "0000101011001100",
23002 => "0000101011001110",
23003 => "0000101011001110",
23004 => "0000101011001110",
23005 => "0000101011010000",
23006 => "0000101011010000",
23007 => "0000101011010000",
23008 => "0000101011010000",
23009 => "0000101011010010",
23010 => "0000101011010010",
23011 => "0000101011010010",
23012 => "0000101011010100",
23013 => "0000101011010100",
23014 => "0000101011010100",
23015 => "0000101011010110",
23016 => "0000101011010110",
23017 => "0000101011010110",
23018 => "0000101011011000",
23019 => "0000101011011000",
23020 => "0000101011011000",
23021 => "0000101011011000",
23022 => "0000101011011010",
23023 => "0000101011011010",
23024 => "0000101011011010",
23025 => "0000101011011100",
23026 => "0000101011011100",
23027 => "0000101011011100",
23028 => "0000101011011110",
23029 => "0000101011011110",
23030 => "0000101011011110",
23031 => "0000101011100000",
23032 => "0000101011100000",
23033 => "0000101011100000",
23034 => "0000101011100010",
23035 => "0000101011100010",
23036 => "0000101011100010",
23037 => "0000101011100010",
23038 => "0000101011100100",
23039 => "0000101011100100",
23040 => "0000101011100100",
23041 => "0000101011100110",
23042 => "0000101011100110",
23043 => "0000101011100110",
23044 => "0000101011101000",
23045 => "0000101011101000",
23046 => "0000101011101000",
23047 => "0000101011101010",
23048 => "0000101011101010",
23049 => "0000101011101010",
23050 => "0000101011101010",
23051 => "0000101011101100",
23052 => "0000101011101100",
23053 => "0000101011101100",
23054 => "0000101011101110",
23055 => "0000101011101110",
23056 => "0000101011101110",
23057 => "0000101011110000",
23058 => "0000101011110000",
23059 => "0000101011110000",
23060 => "0000101011110010",
23061 => "0000101011110010",
23062 => "0000101011110010",
23063 => "0000101011110100",
23064 => "0000101011110100",
23065 => "0000101011110100",
23066 => "0000101011110100",
23067 => "0000101011110110",
23068 => "0000101011110110",
23069 => "0000101011110110",
23070 => "0000101011111000",
23071 => "0000101011111000",
23072 => "0000101011111000",
23073 => "0000101011111010",
23074 => "0000101011111010",
23075 => "0000101011111010",
23076 => "0000101011111100",
23077 => "0000101011111100",
23078 => "0000101011111100",
23079 => "0000101011111110",
23080 => "0000101011111110",
23081 => "0000101011111110",
23082 => "0000101100000000",
23083 => "0000101100000000",
23084 => "0000101100000000",
23085 => "0000101100000000",
23086 => "0000101100000010",
23087 => "0000101100000010",
23088 => "0000101100000010",
23089 => "0000101100000100",
23090 => "0000101100000100",
23091 => "0000101100000100",
23092 => "0000101100000110",
23093 => "0000101100000110",
23094 => "0000101100000110",
23095 => "0000101100001000",
23096 => "0000101100001000",
23097 => "0000101100001000",
23098 => "0000101100001010",
23099 => "0000101100001010",
23100 => "0000101100001010",
23101 => "0000101100001010",
23102 => "0000101100001100",
23103 => "0000101100001100",
23104 => "0000101100001100",
23105 => "0000101100001110",
23106 => "0000101100001110",
23107 => "0000101100001110",
23108 => "0000101100010000",
23109 => "0000101100010000",
23110 => "0000101100010000",
23111 => "0000101100010010",
23112 => "0000101100010010",
23113 => "0000101100010010",
23114 => "0000101100010100",
23115 => "0000101100010100",
23116 => "0000101100010100",
23117 => "0000101100010110",
23118 => "0000101100010110",
23119 => "0000101100010110",
23120 => "0000101100010110",
23121 => "0000101100011000",
23122 => "0000101100011000",
23123 => "0000101100011000",
23124 => "0000101100011010",
23125 => "0000101100011010",
23126 => "0000101100011010",
23127 => "0000101100011100",
23128 => "0000101100011100",
23129 => "0000101100011100",
23130 => "0000101100011110",
23131 => "0000101100011110",
23132 => "0000101100011110",
23133 => "0000101100100000",
23134 => "0000101100100000",
23135 => "0000101100100000",
23136 => "0000101100100010",
23137 => "0000101100100010",
23138 => "0000101100100010",
23139 => "0000101100100100",
23140 => "0000101100100100",
23141 => "0000101100100100",
23142 => "0000101100100100",
23143 => "0000101100100110",
23144 => "0000101100100110",
23145 => "0000101100100110",
23146 => "0000101100101000",
23147 => "0000101100101000",
23148 => "0000101100101000",
23149 => "0000101100101010",
23150 => "0000101100101010",
23151 => "0000101100101010",
23152 => "0000101100101100",
23153 => "0000101100101100",
23154 => "0000101100101100",
23155 => "0000101100101110",
23156 => "0000101100101110",
23157 => "0000101100101110",
23158 => "0000101100110000",
23159 => "0000101100110000",
23160 => "0000101100110000",
23161 => "0000101100110010",
23162 => "0000101100110010",
23163 => "0000101100110010",
23164 => "0000101100110010",
23165 => "0000101100110100",
23166 => "0000101100110100",
23167 => "0000101100110100",
23168 => "0000101100110110",
23169 => "0000101100110110",
23170 => "0000101100110110",
23171 => "0000101100111000",
23172 => "0000101100111000",
23173 => "0000101100111000",
23174 => "0000101100111010",
23175 => "0000101100111010",
23176 => "0000101100111010",
23177 => "0000101100111100",
23178 => "0000101100111100",
23179 => "0000101100111100",
23180 => "0000101100111110",
23181 => "0000101100111110",
23182 => "0000101100111110",
23183 => "0000101101000000",
23184 => "0000101101000000",
23185 => "0000101101000000",
23186 => "0000101101000010",
23187 => "0000101101000010",
23188 => "0000101101000010",
23189 => "0000101101000010",
23190 => "0000101101000100",
23191 => "0000101101000100",
23192 => "0000101101000100",
23193 => "0000101101000110",
23194 => "0000101101000110",
23195 => "0000101101000110",
23196 => "0000101101001000",
23197 => "0000101101001000",
23198 => "0000101101001000",
23199 => "0000101101001010",
23200 => "0000101101001010",
23201 => "0000101101001010",
23202 => "0000101101001100",
23203 => "0000101101001100",
23204 => "0000101101001100",
23205 => "0000101101001110",
23206 => "0000101101001110",
23207 => "0000101101001110",
23208 => "0000101101010000",
23209 => "0000101101010000",
23210 => "0000101101010000",
23211 => "0000101101010010",
23212 => "0000101101010010",
23213 => "0000101101010010",
23214 => "0000101101010100",
23215 => "0000101101010100",
23216 => "0000101101010100",
23217 => "0000101101010100",
23218 => "0000101101010110",
23219 => "0000101101010110",
23220 => "0000101101010110",
23221 => "0000101101011000",
23222 => "0000101101011000",
23223 => "0000101101011000",
23224 => "0000101101011010",
23225 => "0000101101011010",
23226 => "0000101101011010",
23227 => "0000101101011100",
23228 => "0000101101011100",
23229 => "0000101101011100",
23230 => "0000101101011110",
23231 => "0000101101011110",
23232 => "0000101101011110",
23233 => "0000101101100000",
23234 => "0000101101100000",
23235 => "0000101101100000",
23236 => "0000101101100010",
23237 => "0000101101100010",
23238 => "0000101101100010",
23239 => "0000101101100100",
23240 => "0000101101100100",
23241 => "0000101101100100",
23242 => "0000101101100110",
23243 => "0000101101100110",
23244 => "0000101101100110",
23245 => "0000101101101000",
23246 => "0000101101101000",
23247 => "0000101101101000",
23248 => "0000101101101010",
23249 => "0000101101101010",
23250 => "0000101101101010",
23251 => "0000101101101100",
23252 => "0000101101101100",
23253 => "0000101101101100",
23254 => "0000101101101100",
23255 => "0000101101101110",
23256 => "0000101101101110",
23257 => "0000101101101110",
23258 => "0000101101110000",
23259 => "0000101101110000",
23260 => "0000101101110000",
23261 => "0000101101110010",
23262 => "0000101101110010",
23263 => "0000101101110010",
23264 => "0000101101110100",
23265 => "0000101101110100",
23266 => "0000101101110100",
23267 => "0000101101110110",
23268 => "0000101101110110",
23269 => "0000101101110110",
23270 => "0000101101111000",
23271 => "0000101101111000",
23272 => "0000101101111000",
23273 => "0000101101111010",
23274 => "0000101101111010",
23275 => "0000101101111010",
23276 => "0000101101111100",
23277 => "0000101101111100",
23278 => "0000101101111100",
23279 => "0000101101111110",
23280 => "0000101101111110",
23281 => "0000101101111110",
23282 => "0000101110000000",
23283 => "0000101110000000",
23284 => "0000101110000000",
23285 => "0000101110000010",
23286 => "0000101110000010",
23287 => "0000101110000010",
23288 => "0000101110000100",
23289 => "0000101110000100",
23290 => "0000101110000100",
23291 => "0000101110000110",
23292 => "0000101110000110",
23293 => "0000101110000110",
23294 => "0000101110001000",
23295 => "0000101110001000",
23296 => "0000101110001000",
23297 => "0000101110001010",
23298 => "0000101110001010",
23299 => "0000101110001010",
23300 => "0000101110001100",
23301 => "0000101110001100",
23302 => "0000101110001100",
23303 => "0000101110001100",
23304 => "0000101110001110",
23305 => "0000101110001110",
23306 => "0000101110001110",
23307 => "0000101110010000",
23308 => "0000101110010000",
23309 => "0000101110010000",
23310 => "0000101110010010",
23311 => "0000101110010010",
23312 => "0000101110010010",
23313 => "0000101110010100",
23314 => "0000101110010100",
23315 => "0000101110010100",
23316 => "0000101110010110",
23317 => "0000101110010110",
23318 => "0000101110010110",
23319 => "0000101110011000",
23320 => "0000101110011000",
23321 => "0000101110011000",
23322 => "0000101110011010",
23323 => "0000101110011010",
23324 => "0000101110011010",
23325 => "0000101110011100",
23326 => "0000101110011100",
23327 => "0000101110011100",
23328 => "0000101110011110",
23329 => "0000101110011110",
23330 => "0000101110011110",
23331 => "0000101110100000",
23332 => "0000101110100000",
23333 => "0000101110100000",
23334 => "0000101110100010",
23335 => "0000101110100010",
23336 => "0000101110100010",
23337 => "0000101110100100",
23338 => "0000101110100100",
23339 => "0000101110100100",
23340 => "0000101110100110",
23341 => "0000101110100110",
23342 => "0000101110100110",
23343 => "0000101110101000",
23344 => "0000101110101000",
23345 => "0000101110101000",
23346 => "0000101110101010",
23347 => "0000101110101010",
23348 => "0000101110101010",
23349 => "0000101110101100",
23350 => "0000101110101100",
23351 => "0000101110101100",
23352 => "0000101110101110",
23353 => "0000101110101110",
23354 => "0000101110101110",
23355 => "0000101110110000",
23356 => "0000101110110000",
23357 => "0000101110110000",
23358 => "0000101110110010",
23359 => "0000101110110010",
23360 => "0000101110110010",
23361 => "0000101110110100",
23362 => "0000101110110100",
23363 => "0000101110110100",
23364 => "0000101110110110",
23365 => "0000101110110110",
23366 => "0000101110110110",
23367 => "0000101110111000",
23368 => "0000101110111000",
23369 => "0000101110111000",
23370 => "0000101110111010",
23371 => "0000101110111010",
23372 => "0000101110111010",
23373 => "0000101110111100",
23374 => "0000101110111100",
23375 => "0000101110111100",
23376 => "0000101110111110",
23377 => "0000101110111110",
23378 => "0000101110111110",
23379 => "0000101111000000",
23380 => "0000101111000000",
23381 => "0000101111000000",
23382 => "0000101111000010",
23383 => "0000101111000010",
23384 => "0000101111000010",
23385 => "0000101111000100",
23386 => "0000101111000100",
23387 => "0000101111000100",
23388 => "0000101111000110",
23389 => "0000101111000110",
23390 => "0000101111000110",
23391 => "0000101111001000",
23392 => "0000101111001000",
23393 => "0000101111001000",
23394 => "0000101111001010",
23395 => "0000101111001010",
23396 => "0000101111001010",
23397 => "0000101111001100",
23398 => "0000101111001100",
23399 => "0000101111001100",
23400 => "0000101111001110",
23401 => "0000101111001110",
23402 => "0000101111001110",
23403 => "0000101111010000",
23404 => "0000101111010000",
23405 => "0000101111010000",
23406 => "0000101111010010",
23407 => "0000101111010010",
23408 => "0000101111010010",
23409 => "0000101111010100",
23410 => "0000101111010100",
23411 => "0000101111010100",
23412 => "0000101111010110",
23413 => "0000101111010110",
23414 => "0000101111010110",
23415 => "0000101111011000",
23416 => "0000101111011000",
23417 => "0000101111011000",
23418 => "0000101111011010",
23419 => "0000101111011010",
23420 => "0000101111011010",
23421 => "0000101111011100",
23422 => "0000101111011100",
23423 => "0000101111011100",
23424 => "0000101111011110",
23425 => "0000101111011110",
23426 => "0000101111011110",
23427 => "0000101111100000",
23428 => "0000101111100000",
23429 => "0000101111100000",
23430 => "0000101111100010",
23431 => "0000101111100010",
23432 => "0000101111100010",
23433 => "0000101111100100",
23434 => "0000101111100100",
23435 => "0000101111100100",
23436 => "0000101111100110",
23437 => "0000101111100110",
23438 => "0000101111100110",
23439 => "0000101111101000",
23440 => "0000101111101000",
23441 => "0000101111101000",
23442 => "0000101111101010",
23443 => "0000101111101010",
23444 => "0000101111101010",
23445 => "0000101111101100",
23446 => "0000101111101100",
23447 => "0000101111101100",
23448 => "0000101111101110",
23449 => "0000101111101110",
23450 => "0000101111101110",
23451 => "0000101111110000",
23452 => "0000101111110000",
23453 => "0000101111110010",
23454 => "0000101111110010",
23455 => "0000101111110010",
23456 => "0000101111110100",
23457 => "0000101111110100",
23458 => "0000101111110100",
23459 => "0000101111110110",
23460 => "0000101111110110",
23461 => "0000101111110110",
23462 => "0000101111111000",
23463 => "0000101111111000",
23464 => "0000101111111000",
23465 => "0000101111111010",
23466 => "0000101111111010",
23467 => "0000101111111010",
23468 => "0000101111111100",
23469 => "0000101111111100",
23470 => "0000101111111100",
23471 => "0000101111111110",
23472 => "0000101111111110",
23473 => "0000101111111110",
23474 => "0000110000000000",
23475 => "0000110000000000",
23476 => "0000110000000000",
23477 => "0000110000000010",
23478 => "0000110000000010",
23479 => "0000110000000010",
23480 => "0000110000000100",
23481 => "0000110000000100",
23482 => "0000110000000100",
23483 => "0000110000000110",
23484 => "0000110000000110",
23485 => "0000110000000110",
23486 => "0000110000001000",
23487 => "0000110000001000",
23488 => "0000110000001000",
23489 => "0000110000001010",
23490 => "0000110000001010",
23491 => "0000110000001010",
23492 => "0000110000001100",
23493 => "0000110000001100",
23494 => "0000110000001100",
23495 => "0000110000001110",
23496 => "0000110000001110",
23497 => "0000110000001110",
23498 => "0000110000010000",
23499 => "0000110000010000",
23500 => "0000110000010000",
23501 => "0000110000010010",
23502 => "0000110000010010",
23503 => "0000110000010100",
23504 => "0000110000010100",
23505 => "0000110000010100",
23506 => "0000110000010110",
23507 => "0000110000010110",
23508 => "0000110000010110",
23509 => "0000110000011000",
23510 => "0000110000011000",
23511 => "0000110000011000",
23512 => "0000110000011010",
23513 => "0000110000011010",
23514 => "0000110000011010",
23515 => "0000110000011100",
23516 => "0000110000011100",
23517 => "0000110000011100",
23518 => "0000110000011110",
23519 => "0000110000011110",
23520 => "0000110000011110",
23521 => "0000110000100000",
23522 => "0000110000100000",
23523 => "0000110000100000",
23524 => "0000110000100010",
23525 => "0000110000100010",
23526 => "0000110000100010",
23527 => "0000110000100100",
23528 => "0000110000100100",
23529 => "0000110000100100",
23530 => "0000110000100110",
23531 => "0000110000100110",
23532 => "0000110000100110",
23533 => "0000110000101000",
23534 => "0000110000101000",
23535 => "0000110000101000",
23536 => "0000110000101010",
23537 => "0000110000101010",
23538 => "0000110000101100",
23539 => "0000110000101100",
23540 => "0000110000101100",
23541 => "0000110000101110",
23542 => "0000110000101110",
23543 => "0000110000101110",
23544 => "0000110000110000",
23545 => "0000110000110000",
23546 => "0000110000110000",
23547 => "0000110000110010",
23548 => "0000110000110010",
23549 => "0000110000110010",
23550 => "0000110000110100",
23551 => "0000110000110100",
23552 => "0000110000110100",
23553 => "0000110000110110",
23554 => "0000110000110110",
23555 => "0000110000110110",
23556 => "0000110000111000",
23557 => "0000110000111000",
23558 => "0000110000111000",
23559 => "0000110000111010",
23560 => "0000110000111010",
23561 => "0000110000111010",
23562 => "0000110000111100",
23563 => "0000110000111100",
23564 => "0000110000111100",
23565 => "0000110000111110",
23566 => "0000110000111110",
23567 => "0000110001000000",
23568 => "0000110001000000",
23569 => "0000110001000000",
23570 => "0000110001000010",
23571 => "0000110001000010",
23572 => "0000110001000010",
23573 => "0000110001000100",
23574 => "0000110001000100",
23575 => "0000110001000100",
23576 => "0000110001000110",
23577 => "0000110001000110",
23578 => "0000110001000110",
23579 => "0000110001001000",
23580 => "0000110001001000",
23581 => "0000110001001000",
23582 => "0000110001001010",
23583 => "0000110001001010",
23584 => "0000110001001010",
23585 => "0000110001001100",
23586 => "0000110001001100",
23587 => "0000110001001100",
23588 => "0000110001001110",
23589 => "0000110001001110",
23590 => "0000110001001110",
23591 => "0000110001010000",
23592 => "0000110001010000",
23593 => "0000110001010010",
23594 => "0000110001010010",
23595 => "0000110001010010",
23596 => "0000110001010100",
23597 => "0000110001010100",
23598 => "0000110001010100",
23599 => "0000110001010110",
23600 => "0000110001010110",
23601 => "0000110001010110",
23602 => "0000110001011000",
23603 => "0000110001011000",
23604 => "0000110001011000",
23605 => "0000110001011010",
23606 => "0000110001011010",
23607 => "0000110001011010",
23608 => "0000110001011100",
23609 => "0000110001011100",
23610 => "0000110001011100",
23611 => "0000110001011110",
23612 => "0000110001011110",
23613 => "0000110001100000",
23614 => "0000110001100000",
23615 => "0000110001100000",
23616 => "0000110001100010",
23617 => "0000110001100010",
23618 => "0000110001100010",
23619 => "0000110001100100",
23620 => "0000110001100100",
23621 => "0000110001100100",
23622 => "0000110001100110",
23623 => "0000110001100110",
23624 => "0000110001100110",
23625 => "0000110001101000",
23626 => "0000110001101000",
23627 => "0000110001101000",
23628 => "0000110001101010",
23629 => "0000110001101010",
23630 => "0000110001101010",
23631 => "0000110001101100",
23632 => "0000110001101100",
23633 => "0000110001101110",
23634 => "0000110001101110",
23635 => "0000110001101110",
23636 => "0000110001110000",
23637 => "0000110001110000",
23638 => "0000110001110000",
23639 => "0000110001110010",
23640 => "0000110001110010",
23641 => "0000110001110010",
23642 => "0000110001110100",
23643 => "0000110001110100",
23644 => "0000110001110100",
23645 => "0000110001110110",
23646 => "0000110001110110",
23647 => "0000110001110110",
23648 => "0000110001111000",
23649 => "0000110001111000",
23650 => "0000110001111000",
23651 => "0000110001111010",
23652 => "0000110001111010",
23653 => "0000110001111100",
23654 => "0000110001111100",
23655 => "0000110001111100",
23656 => "0000110001111110",
23657 => "0000110001111110",
23658 => "0000110001111110",
23659 => "0000110010000000",
23660 => "0000110010000000",
23661 => "0000110010000000",
23662 => "0000110010000010",
23663 => "0000110010000010",
23664 => "0000110010000010",
23665 => "0000110010000100",
23666 => "0000110010000100",
23667 => "0000110010000100",
23668 => "0000110010000110",
23669 => "0000110010000110",
23670 => "0000110010001000",
23671 => "0000110010001000",
23672 => "0000110010001000",
23673 => "0000110010001010",
23674 => "0000110010001010",
23675 => "0000110010001010",
23676 => "0000110010001100",
23677 => "0000110010001100",
23678 => "0000110010001100",
23679 => "0000110010001110",
23680 => "0000110010001110",
23681 => "0000110010001110",
23682 => "0000110010010000",
23683 => "0000110010010000",
23684 => "0000110010010000",
23685 => "0000110010010010",
23686 => "0000110010010010",
23687 => "0000110010010100",
23688 => "0000110010010100",
23689 => "0000110010010100",
23690 => "0000110010010110",
23691 => "0000110010010110",
23692 => "0000110010010110",
23693 => "0000110010011000",
23694 => "0000110010011000",
23695 => "0000110010011000",
23696 => "0000110010011010",
23697 => "0000110010011010",
23698 => "0000110010011010",
23699 => "0000110010011100",
23700 => "0000110010011100",
23701 => "0000110010011110",
23702 => "0000110010011110",
23703 => "0000110010011110",
23704 => "0000110010100000",
23705 => "0000110010100000",
23706 => "0000110010100000",
23707 => "0000110010100010",
23708 => "0000110010100010",
23709 => "0000110010100010",
23710 => "0000110010100100",
23711 => "0000110010100100",
23712 => "0000110010100100",
23713 => "0000110010100110",
23714 => "0000110010100110",
23715 => "0000110010100110",
23716 => "0000110010101000",
23717 => "0000110010101000",
23718 => "0000110010101010",
23719 => "0000110010101010",
23720 => "0000110010101010",
23721 => "0000110010101100",
23722 => "0000110010101100",
23723 => "0000110010101100",
23724 => "0000110010101110",
23725 => "0000110010101110",
23726 => "0000110010101110",
23727 => "0000110010110000",
23728 => "0000110010110000",
23729 => "0000110010110000",
23730 => "0000110010110010",
23731 => "0000110010110010",
23732 => "0000110010110100",
23733 => "0000110010110100",
23734 => "0000110010110100",
23735 => "0000110010110110",
23736 => "0000110010110110",
23737 => "0000110010110110",
23738 => "0000110010111000",
23739 => "0000110010111000",
23740 => "0000110010111000",
23741 => "0000110010111010",
23742 => "0000110010111010",
23743 => "0000110010111010",
23744 => "0000110010111100",
23745 => "0000110010111100",
23746 => "0000110010111110",
23747 => "0000110010111110",
23748 => "0000110010111110",
23749 => "0000110011000000",
23750 => "0000110011000000",
23751 => "0000110011000000",
23752 => "0000110011000010",
23753 => "0000110011000010",
23754 => "0000110011000010",
23755 => "0000110011000100",
23756 => "0000110011000100",
23757 => "0000110011000110",
23758 => "0000110011000110",
23759 => "0000110011000110",
23760 => "0000110011001000",
23761 => "0000110011001000",
23762 => "0000110011001000",
23763 => "0000110011001010",
23764 => "0000110011001010",
23765 => "0000110011001010",
23766 => "0000110011001100",
23767 => "0000110011001100",
23768 => "0000110011001100",
23769 => "0000110011001110",
23770 => "0000110011001110",
23771 => "0000110011010000",
23772 => "0000110011010000",
23773 => "0000110011010000",
23774 => "0000110011010010",
23775 => "0000110011010010",
23776 => "0000110011010010",
23777 => "0000110011010100",
23778 => "0000110011010100",
23779 => "0000110011010100",
23780 => "0000110011010110",
23781 => "0000110011010110",
23782 => "0000110011011000",
23783 => "0000110011011000",
23784 => "0000110011011000",
23785 => "0000110011011010",
23786 => "0000110011011010",
23787 => "0000110011011010",
23788 => "0000110011011100",
23789 => "0000110011011100",
23790 => "0000110011011100",
23791 => "0000110011011110",
23792 => "0000110011011110",
23793 => "0000110011011110",
23794 => "0000110011100000",
23795 => "0000110011100000",
23796 => "0000110011100010",
23797 => "0000110011100010",
23798 => "0000110011100010",
23799 => "0000110011100100",
23800 => "0000110011100100",
23801 => "0000110011100100",
23802 => "0000110011100110",
23803 => "0000110011100110",
23804 => "0000110011100110",
23805 => "0000110011101000",
23806 => "0000110011101000",
23807 => "0000110011101010",
23808 => "0000110011101010",
23809 => "0000110011101010",
23810 => "0000110011101100",
23811 => "0000110011101100",
23812 => "0000110011101100",
23813 => "0000110011101110",
23814 => "0000110011101110",
23815 => "0000110011101110",
23816 => "0000110011110000",
23817 => "0000110011110000",
23818 => "0000110011110010",
23819 => "0000110011110010",
23820 => "0000110011110010",
23821 => "0000110011110100",
23822 => "0000110011110100",
23823 => "0000110011110100",
23824 => "0000110011110110",
23825 => "0000110011110110",
23826 => "0000110011110110",
23827 => "0000110011111000",
23828 => "0000110011111000",
23829 => "0000110011111010",
23830 => "0000110011111010",
23831 => "0000110011111010",
23832 => "0000110011111100",
23833 => "0000110011111100",
23834 => "0000110011111100",
23835 => "0000110011111110",
23836 => "0000110011111110",
23837 => "0000110011111110",
23838 => "0000110100000000",
23839 => "0000110100000000",
23840 => "0000110100000010",
23841 => "0000110100000010",
23842 => "0000110100000010",
23843 => "0000110100000100",
23844 => "0000110100000100",
23845 => "0000110100000100",
23846 => "0000110100000110",
23847 => "0000110100000110",
23848 => "0000110100000110",
23849 => "0000110100001000",
23850 => "0000110100001000",
23851 => "0000110100001010",
23852 => "0000110100001010",
23853 => "0000110100001010",
23854 => "0000110100001100",
23855 => "0000110100001100",
23856 => "0000110100001100",
23857 => "0000110100001110",
23858 => "0000110100001110",
23859 => "0000110100010000",
23860 => "0000110100010000",
23861 => "0000110100010000",
23862 => "0000110100010010",
23863 => "0000110100010010",
23864 => "0000110100010010",
23865 => "0000110100010100",
23866 => "0000110100010100",
23867 => "0000110100010100",
23868 => "0000110100010110",
23869 => "0000110100010110",
23870 => "0000110100011000",
23871 => "0000110100011000",
23872 => "0000110100011000",
23873 => "0000110100011010",
23874 => "0000110100011010",
23875 => "0000110100011010",
23876 => "0000110100011100",
23877 => "0000110100011100",
23878 => "0000110100011100",
23879 => "0000110100011110",
23880 => "0000110100011110",
23881 => "0000110100100000",
23882 => "0000110100100000",
23883 => "0000110100100000",
23884 => "0000110100100010",
23885 => "0000110100100010",
23886 => "0000110100100010",
23887 => "0000110100100100",
23888 => "0000110100100100",
23889 => "0000110100100110",
23890 => "0000110100100110",
23891 => "0000110100100110",
23892 => "0000110100101000",
23893 => "0000110100101000",
23894 => "0000110100101000",
23895 => "0000110100101010",
23896 => "0000110100101010",
23897 => "0000110100101100",
23898 => "0000110100101100",
23899 => "0000110100101100",
23900 => "0000110100101110",
23901 => "0000110100101110",
23902 => "0000110100101110",
23903 => "0000110100110000",
23904 => "0000110100110000",
23905 => "0000110100110000",
23906 => "0000110100110010",
23907 => "0000110100110010",
23908 => "0000110100110100",
23909 => "0000110100110100",
23910 => "0000110100110100",
23911 => "0000110100110110",
23912 => "0000110100110110",
23913 => "0000110100110110",
23914 => "0000110100111000",
23915 => "0000110100111000",
23916 => "0000110100111010",
23917 => "0000110100111010",
23918 => "0000110100111010",
23919 => "0000110100111100",
23920 => "0000110100111100",
23921 => "0000110100111100",
23922 => "0000110100111110",
23923 => "0000110100111110",
23924 => "0000110100111110",
23925 => "0000110101000000",
23926 => "0000110101000000",
23927 => "0000110101000010",
23928 => "0000110101000010",
23929 => "0000110101000010",
23930 => "0000110101000100",
23931 => "0000110101000100",
23932 => "0000110101000100",
23933 => "0000110101000110",
23934 => "0000110101000110",
23935 => "0000110101001000",
23936 => "0000110101001000",
23937 => "0000110101001000",
23938 => "0000110101001010",
23939 => "0000110101001010",
23940 => "0000110101001010",
23941 => "0000110101001100",
23942 => "0000110101001100",
23943 => "0000110101001110",
23944 => "0000110101001110",
23945 => "0000110101001110",
23946 => "0000110101010000",
23947 => "0000110101010000",
23948 => "0000110101010000",
23949 => "0000110101010010",
23950 => "0000110101010010",
23951 => "0000110101010100",
23952 => "0000110101010100",
23953 => "0000110101010100",
23954 => "0000110101010110",
23955 => "0000110101010110",
23956 => "0000110101010110",
23957 => "0000110101011000",
23958 => "0000110101011000",
23959 => "0000110101011010",
23960 => "0000110101011010",
23961 => "0000110101011010",
23962 => "0000110101011100",
23963 => "0000110101011100",
23964 => "0000110101011100",
23965 => "0000110101011110",
23966 => "0000110101011110",
23967 => "0000110101100000",
23968 => "0000110101100000",
23969 => "0000110101100000",
23970 => "0000110101100010",
23971 => "0000110101100010",
23972 => "0000110101100010",
23973 => "0000110101100100",
23974 => "0000110101100100",
23975 => "0000110101100110",
23976 => "0000110101100110",
23977 => "0000110101100110",
23978 => "0000110101101000",
23979 => "0000110101101000",
23980 => "0000110101101000",
23981 => "0000110101101010",
23982 => "0000110101101010",
23983 => "0000110101101100",
23984 => "0000110101101100",
23985 => "0000110101101100",
23986 => "0000110101101110",
23987 => "0000110101101110",
23988 => "0000110101101110",
23989 => "0000110101110000",
23990 => "0000110101110000",
23991 => "0000110101110010",
23992 => "0000110101110010",
23993 => "0000110101110010",
23994 => "0000110101110100",
23995 => "0000110101110100",
23996 => "0000110101110100",
23997 => "0000110101110110",
23998 => "0000110101110110",
23999 => "0000110101111000",
24000 => "0000110101111000",
24001 => "0000110101111000",
24002 => "0000110101111010",
24003 => "0000110101111010",
24004 => "0000110101111010",
24005 => "0000110101111100",
24006 => "0000110101111100",
24007 => "0000110101111110",
24008 => "0000110101111110",
24009 => "0000110101111110",
24010 => "0000110110000000",
24011 => "0000110110000000",
24012 => "0000110110000000",
24013 => "0000110110000010",
24014 => "0000110110000010",
24015 => "0000110110000100",
24016 => "0000110110000100",
24017 => "0000110110000100",
24018 => "0000110110000110",
24019 => "0000110110000110",
24020 => "0000110110000110",
24021 => "0000110110001000",
24022 => "0000110110001000",
24023 => "0000110110001010",
24024 => "0000110110001010",
24025 => "0000110110001010",
24026 => "0000110110001100",
24027 => "0000110110001100",
24028 => "0000110110001100",
24029 => "0000110110001110",
24030 => "0000110110001110",
24031 => "0000110110010000",
24032 => "0000110110010000",
24033 => "0000110110010000",
24034 => "0000110110010010",
24035 => "0000110110010010",
24036 => "0000110110010100",
24037 => "0000110110010100",
24038 => "0000110110010100",
24039 => "0000110110010110",
24040 => "0000110110010110",
24041 => "0000110110010110",
24042 => "0000110110011000",
24043 => "0000110110011000",
24044 => "0000110110011010",
24045 => "0000110110011010",
24046 => "0000110110011010",
24047 => "0000110110011100",
24048 => "0000110110011100",
24049 => "0000110110011100",
24050 => "0000110110011110",
24051 => "0000110110011110",
24052 => "0000110110100000",
24053 => "0000110110100000",
24054 => "0000110110100000",
24055 => "0000110110100010",
24056 => "0000110110100010",
24057 => "0000110110100010",
24058 => "0000110110100100",
24059 => "0000110110100100",
24060 => "0000110110100110",
24061 => "0000110110100110",
24062 => "0000110110100110",
24063 => "0000110110101000",
24064 => "0000110110101000",
24065 => "0000110110101010",
24066 => "0000110110101010",
24067 => "0000110110101010",
24068 => "0000110110101100",
24069 => "0000110110101100",
24070 => "0000110110101100",
24071 => "0000110110101110",
24072 => "0000110110101110",
24073 => "0000110110110000",
24074 => "0000110110110000",
24075 => "0000110110110000",
24076 => "0000110110110010",
24077 => "0000110110110010",
24078 => "0000110110110100",
24079 => "0000110110110100",
24080 => "0000110110110100",
24081 => "0000110110110110",
24082 => "0000110110110110",
24083 => "0000110110110110",
24084 => "0000110110111000",
24085 => "0000110110111000",
24086 => "0000110110111010",
24087 => "0000110110111010",
24088 => "0000110110111010",
24089 => "0000110110111100",
24090 => "0000110110111100",
24091 => "0000110110111100",
24092 => "0000110110111110",
24093 => "0000110110111110",
24094 => "0000110111000000",
24095 => "0000110111000000",
24096 => "0000110111000000",
24097 => "0000110111000010",
24098 => "0000110111000010",
24099 => "0000110111000100",
24100 => "0000110111000100",
24101 => "0000110111000100",
24102 => "0000110111000110",
24103 => "0000110111000110",
24104 => "0000110111000110",
24105 => "0000110111001000",
24106 => "0000110111001000",
24107 => "0000110111001010",
24108 => "0000110111001010",
24109 => "0000110111001010",
24110 => "0000110111001100",
24111 => "0000110111001100",
24112 => "0000110111001110",
24113 => "0000110111001110",
24114 => "0000110111001110",
24115 => "0000110111010000",
24116 => "0000110111010000",
24117 => "0000110111010000",
24118 => "0000110111010010",
24119 => "0000110111010010",
24120 => "0000110111010100",
24121 => "0000110111010100",
24122 => "0000110111010100",
24123 => "0000110111010110",
24124 => "0000110111010110",
24125 => "0000110111011000",
24126 => "0000110111011000",
24127 => "0000110111011000",
24128 => "0000110111011010",
24129 => "0000110111011010",
24130 => "0000110111011010",
24131 => "0000110111011100",
24132 => "0000110111011100",
24133 => "0000110111011110",
24134 => "0000110111011110",
24135 => "0000110111011110",
24136 => "0000110111100000",
24137 => "0000110111100000",
24138 => "0000110111100010",
24139 => "0000110111100010",
24140 => "0000110111100010",
24141 => "0000110111100100",
24142 => "0000110111100100",
24143 => "0000110111100110",
24144 => "0000110111100110",
24145 => "0000110111100110",
24146 => "0000110111101000",
24147 => "0000110111101000",
24148 => "0000110111101000",
24149 => "0000110111101010",
24150 => "0000110111101010",
24151 => "0000110111101100",
24152 => "0000110111101100",
24153 => "0000110111101100",
24154 => "0000110111101110",
24155 => "0000110111101110",
24156 => "0000110111110000",
24157 => "0000110111110000",
24158 => "0000110111110000",
24159 => "0000110111110010",
24160 => "0000110111110010",
24161 => "0000110111110010",
24162 => "0000110111110100",
24163 => "0000110111110100",
24164 => "0000110111110110",
24165 => "0000110111110110",
24166 => "0000110111110110",
24167 => "0000110111111000",
24168 => "0000110111111000",
24169 => "0000110111111010",
24170 => "0000110111111010",
24171 => "0000110111111010",
24172 => "0000110111111100",
24173 => "0000110111111100",
24174 => "0000110111111110",
24175 => "0000110111111110",
24176 => "0000110111111110",
24177 => "0000111000000000",
24178 => "0000111000000000",
24179 => "0000111000000000",
24180 => "0000111000000010",
24181 => "0000111000000010",
24182 => "0000111000000100",
24183 => "0000111000000100",
24184 => "0000111000000100",
24185 => "0000111000000110",
24186 => "0000111000000110",
24187 => "0000111000001000",
24188 => "0000111000001000",
24189 => "0000111000001000",
24190 => "0000111000001010",
24191 => "0000111000001010",
24192 => "0000111000001100",
24193 => "0000111000001100",
24194 => "0000111000001100",
24195 => "0000111000001110",
24196 => "0000111000001110",
24197 => "0000111000010000",
24198 => "0000111000010000",
24199 => "0000111000010000",
24200 => "0000111000010010",
24201 => "0000111000010010",
24202 => "0000111000010010",
24203 => "0000111000010100",
24204 => "0000111000010100",
24205 => "0000111000010110",
24206 => "0000111000010110",
24207 => "0000111000010110",
24208 => "0000111000011000",
24209 => "0000111000011000",
24210 => "0000111000011010",
24211 => "0000111000011010",
24212 => "0000111000011010",
24213 => "0000111000011100",
24214 => "0000111000011100",
24215 => "0000111000011110",
24216 => "0000111000011110",
24217 => "0000111000011110",
24218 => "0000111000100000",
24219 => "0000111000100000",
24220 => "0000111000100010",
24221 => "0000111000100010",
24222 => "0000111000100010",
24223 => "0000111000100100",
24224 => "0000111000100100",
24225 => "0000111000100100",
24226 => "0000111000100110",
24227 => "0000111000100110",
24228 => "0000111000101000",
24229 => "0000111000101000",
24230 => "0000111000101000",
24231 => "0000111000101010",
24232 => "0000111000101010",
24233 => "0000111000101100",
24234 => "0000111000101100",
24235 => "0000111000101100",
24236 => "0000111000101110",
24237 => "0000111000101110",
24238 => "0000111000110000",
24239 => "0000111000110000",
24240 => "0000111000110000",
24241 => "0000111000110010",
24242 => "0000111000110010",
24243 => "0000111000110100",
24244 => "0000111000110100",
24245 => "0000111000110100",
24246 => "0000111000110110",
24247 => "0000111000110110",
24248 => "0000111000111000",
24249 => "0000111000111000",
24250 => "0000111000111000",
24251 => "0000111000111010",
24252 => "0000111000111010",
24253 => "0000111000111100",
24254 => "0000111000111100",
24255 => "0000111000111100",
24256 => "0000111000111110",
24257 => "0000111000111110",
24258 => "0000111001000000",
24259 => "0000111001000000",
24260 => "0000111001000000",
24261 => "0000111001000010",
24262 => "0000111001000010",
24263 => "0000111001000010",
24264 => "0000111001000100",
24265 => "0000111001000100",
24266 => "0000111001000110",
24267 => "0000111001000110",
24268 => "0000111001000110",
24269 => "0000111001001000",
24270 => "0000111001001000",
24271 => "0000111001001010",
24272 => "0000111001001010",
24273 => "0000111001001010",
24274 => "0000111001001100",
24275 => "0000111001001100",
24276 => "0000111001001110",
24277 => "0000111001001110",
24278 => "0000111001001110",
24279 => "0000111001010000",
24280 => "0000111001010000",
24281 => "0000111001010010",
24282 => "0000111001010010",
24283 => "0000111001010010",
24284 => "0000111001010100",
24285 => "0000111001010100",
24286 => "0000111001010110",
24287 => "0000111001010110",
24288 => "0000111001010110",
24289 => "0000111001011000",
24290 => "0000111001011000",
24291 => "0000111001011010",
24292 => "0000111001011010",
24293 => "0000111001011010",
24294 => "0000111001011100",
24295 => "0000111001011100",
24296 => "0000111001011110",
24297 => "0000111001011110",
24298 => "0000111001011110",
24299 => "0000111001100000",
24300 => "0000111001100000",
24301 => "0000111001100010",
24302 => "0000111001100010",
24303 => "0000111001100010",
24304 => "0000111001100100",
24305 => "0000111001100100",
24306 => "0000111001100110",
24307 => "0000111001100110",
24308 => "0000111001100110",
24309 => "0000111001101000",
24310 => "0000111001101000",
24311 => "0000111001101010",
24312 => "0000111001101010",
24313 => "0000111001101010",
24314 => "0000111001101100",
24315 => "0000111001101100",
24316 => "0000111001101110",
24317 => "0000111001101110",
24318 => "0000111001101110",
24319 => "0000111001110000",
24320 => "0000111001110000",
24321 => "0000111001110010",
24322 => "0000111001110010",
24323 => "0000111001110010",
24324 => "0000111001110100",
24325 => "0000111001110100",
24326 => "0000111001110110",
24327 => "0000111001110110",
24328 => "0000111001110110",
24329 => "0000111001111000",
24330 => "0000111001111000",
24331 => "0000111001111010",
24332 => "0000111001111010",
24333 => "0000111001111010",
24334 => "0000111001111100",
24335 => "0000111001111100",
24336 => "0000111001111110",
24337 => "0000111001111110",
24338 => "0000111001111110",
24339 => "0000111010000000",
24340 => "0000111010000000",
24341 => "0000111010000010",
24342 => "0000111010000010",
24343 => "0000111010000010",
24344 => "0000111010000100",
24345 => "0000111010000100",
24346 => "0000111010000110",
24347 => "0000111010000110",
24348 => "0000111010000110",
24349 => "0000111010001000",
24350 => "0000111010001000",
24351 => "0000111010001010",
24352 => "0000111010001010",
24353 => "0000111010001010",
24354 => "0000111010001100",
24355 => "0000111010001100",
24356 => "0000111010001110",
24357 => "0000111010001110",
24358 => "0000111010001110",
24359 => "0000111010010000",
24360 => "0000111010010000",
24361 => "0000111010010010",
24362 => "0000111010010010",
24363 => "0000111010010010",
24364 => "0000111010010100",
24365 => "0000111010010100",
24366 => "0000111010010110",
24367 => "0000111010010110",
24368 => "0000111010010110",
24369 => "0000111010011000",
24370 => "0000111010011000",
24371 => "0000111010011010",
24372 => "0000111010011010",
24373 => "0000111010011100",
24374 => "0000111010011100",
24375 => "0000111010011100",
24376 => "0000111010011110",
24377 => "0000111010011110",
24378 => "0000111010100000",
24379 => "0000111010100000",
24380 => "0000111010100000",
24381 => "0000111010100010",
24382 => "0000111010100010",
24383 => "0000111010100100",
24384 => "0000111010100100",
24385 => "0000111010100100",
24386 => "0000111010100110",
24387 => "0000111010100110",
24388 => "0000111010101000",
24389 => "0000111010101000",
24390 => "0000111010101000",
24391 => "0000111010101010",
24392 => "0000111010101010",
24393 => "0000111010101100",
24394 => "0000111010101100",
24395 => "0000111010101100",
24396 => "0000111010101110",
24397 => "0000111010101110",
24398 => "0000111010110000",
24399 => "0000111010110000",
24400 => "0000111010110000",
24401 => "0000111010110010",
24402 => "0000111010110010",
24403 => "0000111010110100",
24404 => "0000111010110100",
24405 => "0000111010110100",
24406 => "0000111010110110",
24407 => "0000111010110110",
24408 => "0000111010111000",
24409 => "0000111010111000",
24410 => "0000111010111010",
24411 => "0000111010111010",
24412 => "0000111010111010",
24413 => "0000111010111100",
24414 => "0000111010111100",
24415 => "0000111010111110",
24416 => "0000111010111110",
24417 => "0000111010111110",
24418 => "0000111011000000",
24419 => "0000111011000000",
24420 => "0000111011000010",
24421 => "0000111011000010",
24422 => "0000111011000010",
24423 => "0000111011000100",
24424 => "0000111011000100",
24425 => "0000111011000110",
24426 => "0000111011000110",
24427 => "0000111011000110",
24428 => "0000111011001000",
24429 => "0000111011001000",
24430 => "0000111011001010",
24431 => "0000111011001010",
24432 => "0000111011001100",
24433 => "0000111011001100",
24434 => "0000111011001100",
24435 => "0000111011001110",
24436 => "0000111011001110",
24437 => "0000111011010000",
24438 => "0000111011010000",
24439 => "0000111011010000",
24440 => "0000111011010010",
24441 => "0000111011010010",
24442 => "0000111011010100",
24443 => "0000111011010100",
24444 => "0000111011010100",
24445 => "0000111011010110",
24446 => "0000111011010110",
24447 => "0000111011011000",
24448 => "0000111011011000",
24449 => "0000111011011000",
24450 => "0000111011011010",
24451 => "0000111011011010",
24452 => "0000111011011100",
24453 => "0000111011011100",
24454 => "0000111011011110",
24455 => "0000111011011110",
24456 => "0000111011011110",
24457 => "0000111011100000",
24458 => "0000111011100000",
24459 => "0000111011100010",
24460 => "0000111011100010",
24461 => "0000111011100010",
24462 => "0000111011100100",
24463 => "0000111011100100",
24464 => "0000111011100110",
24465 => "0000111011100110",
24466 => "0000111011100110",
24467 => "0000111011101000",
24468 => "0000111011101000",
24469 => "0000111011101010",
24470 => "0000111011101010",
24471 => "0000111011101100",
24472 => "0000111011101100",
24473 => "0000111011101100",
24474 => "0000111011101110",
24475 => "0000111011101110",
24476 => "0000111011110000",
24477 => "0000111011110000",
24478 => "0000111011110000",
24479 => "0000111011110010",
24480 => "0000111011110010",
24481 => "0000111011110100",
24482 => "0000111011110100",
24483 => "0000111011110100",
24484 => "0000111011110110",
24485 => "0000111011110110",
24486 => "0000111011111000",
24487 => "0000111011111000",
24488 => "0000111011111010",
24489 => "0000111011111010",
24490 => "0000111011111010",
24491 => "0000111011111100",
24492 => "0000111011111100",
24493 => "0000111011111110",
24494 => "0000111011111110",
24495 => "0000111011111110",
24496 => "0000111100000000",
24497 => "0000111100000000",
24498 => "0000111100000010",
24499 => "0000111100000010",
24500 => "0000111100000010",
24501 => "0000111100000100",
24502 => "0000111100000100",
24503 => "0000111100000110",
24504 => "0000111100000110",
24505 => "0000111100001000",
24506 => "0000111100001000",
24507 => "0000111100001000",
24508 => "0000111100001010",
24509 => "0000111100001010",
24510 => "0000111100001100",
24511 => "0000111100001100",
24512 => "0000111100001100",
24513 => "0000111100001110",
24514 => "0000111100001110",
24515 => "0000111100010000",
24516 => "0000111100010000",
24517 => "0000111100010010",
24518 => "0000111100010010",
24519 => "0000111100010010",
24520 => "0000111100010100",
24521 => "0000111100010100",
24522 => "0000111100010110",
24523 => "0000111100010110",
24524 => "0000111100010110",
24525 => "0000111100011000",
24526 => "0000111100011000",
24527 => "0000111100011010",
24528 => "0000111100011010",
24529 => "0000111100011100",
24530 => "0000111100011100",
24531 => "0000111100011100",
24532 => "0000111100011110",
24533 => "0000111100011110",
24534 => "0000111100100000",
24535 => "0000111100100000",
24536 => "0000111100100000",
24537 => "0000111100100010",
24538 => "0000111100100010",
24539 => "0000111100100100",
24540 => "0000111100100100",
24541 => "0000111100100110",
24542 => "0000111100100110",
24543 => "0000111100100110",
24544 => "0000111100101000",
24545 => "0000111100101000",
24546 => "0000111100101010",
24547 => "0000111100101010",
24548 => "0000111100101010",
24549 => "0000111100101100",
24550 => "0000111100101100",
24551 => "0000111100101110",
24552 => "0000111100101110",
24553 => "0000111100110000",
24554 => "0000111100110000",
24555 => "0000111100110000",
24556 => "0000111100110010",
24557 => "0000111100110010",
24558 => "0000111100110100",
24559 => "0000111100110100",
24560 => "0000111100110100",
24561 => "0000111100110110",
24562 => "0000111100110110",
24563 => "0000111100111000",
24564 => "0000111100111000",
24565 => "0000111100111010",
24566 => "0000111100111010",
24567 => "0000111100111010",
24568 => "0000111100111100",
24569 => "0000111100111100",
24570 => "0000111100111110",
24571 => "0000111100111110",
24572 => "0000111100111110",
24573 => "0000111101000000",
24574 => "0000111101000000",
24575 => "0000111101000010",
24576 => "0000111101000010",
24577 => "0000111101000100",
24578 => "0000111101000100",
24579 => "0000111101000100",
24580 => "0000111101000110",
24581 => "0000111101000110",
24582 => "0000111101001000",
24583 => "0000111101001000",
24584 => "0000111101001010",
24585 => "0000111101001010",
24586 => "0000111101001010",
24587 => "0000111101001100",
24588 => "0000111101001100",
24589 => "0000111101001110",
24590 => "0000111101001110",
24591 => "0000111101001110",
24592 => "0000111101010000",
24593 => "0000111101010000",
24594 => "0000111101010010",
24595 => "0000111101010010",
24596 => "0000111101010100",
24597 => "0000111101010100",
24598 => "0000111101010100",
24599 => "0000111101010110",
24600 => "0000111101010110",
24601 => "0000111101011000",
24602 => "0000111101011000",
24603 => "0000111101011010",
24604 => "0000111101011010",
24605 => "0000111101011010",
24606 => "0000111101011100",
24607 => "0000111101011100",
24608 => "0000111101011110",
24609 => "0000111101011110",
24610 => "0000111101100000",
24611 => "0000111101100000",
24612 => "0000111101100000",
24613 => "0000111101100010",
24614 => "0000111101100010",
24615 => "0000111101100100",
24616 => "0000111101100100",
24617 => "0000111101100100",
24618 => "0000111101100110",
24619 => "0000111101100110",
24620 => "0000111101101000",
24621 => "0000111101101000",
24622 => "0000111101101010",
24623 => "0000111101101010",
24624 => "0000111101101010",
24625 => "0000111101101100",
24626 => "0000111101101100",
24627 => "0000111101101110",
24628 => "0000111101101110",
24629 => "0000111101110000",
24630 => "0000111101110000",
24631 => "0000111101110000",
24632 => "0000111101110010",
24633 => "0000111101110010",
24634 => "0000111101110100",
24635 => "0000111101110100",
24636 => "0000111101110110",
24637 => "0000111101110110",
24638 => "0000111101110110",
24639 => "0000111101111000",
24640 => "0000111101111000",
24641 => "0000111101111010",
24642 => "0000111101111010",
24643 => "0000111101111010",
24644 => "0000111101111100",
24645 => "0000111101111100",
24646 => "0000111101111110",
24647 => "0000111101111110",
24648 => "0000111110000000",
24649 => "0000111110000000",
24650 => "0000111110000000",
24651 => "0000111110000010",
24652 => "0000111110000010",
24653 => "0000111110000100",
24654 => "0000111110000100",
24655 => "0000111110000110",
24656 => "0000111110000110",
24657 => "0000111110000110",
24658 => "0000111110001000",
24659 => "0000111110001000",
24660 => "0000111110001010",
24661 => "0000111110001010",
24662 => "0000111110001100",
24663 => "0000111110001100",
24664 => "0000111110001100",
24665 => "0000111110001110",
24666 => "0000111110001110",
24667 => "0000111110010000",
24668 => "0000111110010000",
24669 => "0000111110010010",
24670 => "0000111110010010",
24671 => "0000111110010010",
24672 => "0000111110010100",
24673 => "0000111110010100",
24674 => "0000111110010110",
24675 => "0000111110010110",
24676 => "0000111110011000",
24677 => "0000111110011000",
24678 => "0000111110011000",
24679 => "0000111110011010",
24680 => "0000111110011010",
24681 => "0000111110011100",
24682 => "0000111110011100",
24683 => "0000111110011110",
24684 => "0000111110011110",
24685 => "0000111110011110",
24686 => "0000111110100000",
24687 => "0000111110100000",
24688 => "0000111110100010",
24689 => "0000111110100010",
24690 => "0000111110100100",
24691 => "0000111110100100",
24692 => "0000111110100100",
24693 => "0000111110100110",
24694 => "0000111110100110",
24695 => "0000111110101000",
24696 => "0000111110101000",
24697 => "0000111110101010",
24698 => "0000111110101010",
24699 => "0000111110101010",
24700 => "0000111110101100",
24701 => "0000111110101100",
24702 => "0000111110101110",
24703 => "0000111110101110",
24704 => "0000111110110000",
24705 => "0000111110110000",
24706 => "0000111110110000",
24707 => "0000111110110010",
24708 => "0000111110110010",
24709 => "0000111110110100",
24710 => "0000111110110100",
24711 => "0000111110110110",
24712 => "0000111110110110",
24713 => "0000111110110110",
24714 => "0000111110111000",
24715 => "0000111110111000",
24716 => "0000111110111010",
24717 => "0000111110111010",
24718 => "0000111110111100",
24719 => "0000111110111100",
24720 => "0000111110111100",
24721 => "0000111110111110",
24722 => "0000111110111110",
24723 => "0000111111000000",
24724 => "0000111111000000",
24725 => "0000111111000010",
24726 => "0000111111000010",
24727 => "0000111111000010",
24728 => "0000111111000100",
24729 => "0000111111000100",
24730 => "0000111111000110",
24731 => "0000111111000110",
24732 => "0000111111001000",
24733 => "0000111111001000",
24734 => "0000111111001010",
24735 => "0000111111001010",
24736 => "0000111111001010",
24737 => "0000111111001100",
24738 => "0000111111001100",
24739 => "0000111111001110",
24740 => "0000111111001110",
24741 => "0000111111010000",
24742 => "0000111111010000",
24743 => "0000111111010000",
24744 => "0000111111010010",
24745 => "0000111111010010",
24746 => "0000111111010100",
24747 => "0000111111010100",
24748 => "0000111111010110",
24749 => "0000111111010110",
24750 => "0000111111010110",
24751 => "0000111111011000",
24752 => "0000111111011000",
24753 => "0000111111011010",
24754 => "0000111111011010",
24755 => "0000111111011100",
24756 => "0000111111011100",
24757 => "0000111111011100",
24758 => "0000111111011110",
24759 => "0000111111011110",
24760 => "0000111111100000",
24761 => "0000111111100000",
24762 => "0000111111100010",
24763 => "0000111111100010",
24764 => "0000111111100100",
24765 => "0000111111100100",
24766 => "0000111111100100",
24767 => "0000111111100110",
24768 => "0000111111100110",
24769 => "0000111111101000",
24770 => "0000111111101000",
24771 => "0000111111101010",
24772 => "0000111111101010",
24773 => "0000111111101010",
24774 => "0000111111101100",
24775 => "0000111111101100",
24776 => "0000111111101110",
24777 => "0000111111101110",
24778 => "0000111111110000",
24779 => "0000111111110000",
24780 => "0000111111110000",
24781 => "0000111111110010",
24782 => "0000111111110010",
24783 => "0000111111110100",
24784 => "0000111111110100",
24785 => "0000111111110110",
24786 => "0000111111110110",
24787 => "0000111111111000",
24788 => "0000111111111000",
24789 => "0000111111111000",
24790 => "0000111111111010",
24791 => "0000111111111010",
24792 => "0000111111111100",
24793 => "0000111111111100",
24794 => "0000111111111110",
24795 => "0000111111111110",
24796 => "0000111111111110",
24797 => "0001000000000000",
24798 => "0001000000000000",
24799 => "0001000000000000",
24800 => "0001000000000100",
24801 => "0001000000000100",
24802 => "0001000000000100",
24803 => "0001000000000100",
24804 => "0001000000000100",
24805 => "0001000000001000",
24806 => "0001000000001000",
24807 => "0001000000001000",
24808 => "0001000000001000",
24809 => "0001000000001100",
24810 => "0001000000001100",
24811 => "0001000000001100",
24812 => "0001000000001100",
24813 => "0001000000001100",
24814 => "0001000000010000",
24815 => "0001000000010000",
24816 => "0001000000010000",
24817 => "0001000000010000",
24818 => "0001000000010100",
24819 => "0001000000010100",
24820 => "0001000000010100",
24821 => "0001000000010100",
24822 => "0001000000010100",
24823 => "0001000000011000",
24824 => "0001000000011000",
24825 => "0001000000011000",
24826 => "0001000000011000",
24827 => "0001000000011100",
24828 => "0001000000011100",
24829 => "0001000000011100",
24830 => "0001000000011100",
24831 => "0001000000011100",
24832 => "0001000000100000",
24833 => "0001000000100000",
24834 => "0001000000100000",
24835 => "0001000000100000",
24836 => "0001000000100100",
24837 => "0001000000100100",
24838 => "0001000000100100",
24839 => "0001000000100100",
24840 => "0001000000100100",
24841 => "0001000000101000",
24842 => "0001000000101000",
24843 => "0001000000101000",
24844 => "0001000000101000",
24845 => "0001000000101100",
24846 => "0001000000101100",
24847 => "0001000000101100",
24848 => "0001000000101100",
24849 => "0001000000101100",
24850 => "0001000000110000",
24851 => "0001000000110000",
24852 => "0001000000110000",
24853 => "0001000000110000",
24854 => "0001000000110000",
24855 => "0001000000110100",
24856 => "0001000000110100",
24857 => "0001000000110100",
24858 => "0001000000110100",
24859 => "0001000000111000",
24860 => "0001000000111000",
24861 => "0001000000111000",
24862 => "0001000000111000",
24863 => "0001000000111000",
24864 => "0001000000111100",
24865 => "0001000000111100",
24866 => "0001000000111100",
24867 => "0001000000111100",
24868 => "0001000001000000",
24869 => "0001000001000000",
24870 => "0001000001000000",
24871 => "0001000001000000",
24872 => "0001000001000000",
24873 => "0001000001000100",
24874 => "0001000001000100",
24875 => "0001000001000100",
24876 => "0001000001000100",
24877 => "0001000001001000",
24878 => "0001000001001000",
24879 => "0001000001001000",
24880 => "0001000001001000",
24881 => "0001000001001000",
24882 => "0001000001001100",
24883 => "0001000001001100",
24884 => "0001000001001100",
24885 => "0001000001001100",
24886 => "0001000001010000",
24887 => "0001000001010000",
24888 => "0001000001010000",
24889 => "0001000001010000",
24890 => "0001000001010000",
24891 => "0001000001010100",
24892 => "0001000001010100",
24893 => "0001000001010100",
24894 => "0001000001010100",
24895 => "0001000001011000",
24896 => "0001000001011000",
24897 => "0001000001011000",
24898 => "0001000001011000",
24899 => "0001000001011000",
24900 => "0001000001011100",
24901 => "0001000001011100",
24902 => "0001000001011100",
24903 => "0001000001011100",
24904 => "0001000001100000",
24905 => "0001000001100000",
24906 => "0001000001100000",
24907 => "0001000001100000",
24908 => "0001000001100000",
24909 => "0001000001100100",
24910 => "0001000001100100",
24911 => "0001000001100100",
24912 => "0001000001100100",
24913 => "0001000001101000",
24914 => "0001000001101000",
24915 => "0001000001101000",
24916 => "0001000001101000",
24917 => "0001000001101100",
24918 => "0001000001101100",
24919 => "0001000001101100",
24920 => "0001000001101100",
24921 => "0001000001101100",
24922 => "0001000001110000",
24923 => "0001000001110000",
24924 => "0001000001110000",
24925 => "0001000001110000",
24926 => "0001000001110100",
24927 => "0001000001110100",
24928 => "0001000001110100",
24929 => "0001000001110100",
24930 => "0001000001110100",
24931 => "0001000001111000",
24932 => "0001000001111000",
24933 => "0001000001111000",
24934 => "0001000001111000",
24935 => "0001000001111100",
24936 => "0001000001111100",
24937 => "0001000001111100",
24938 => "0001000001111100",
24939 => "0001000001111100",
24940 => "0001000010000000",
24941 => "0001000010000000",
24942 => "0001000010000000",
24943 => "0001000010000000",
24944 => "0001000010000100",
24945 => "0001000010000100",
24946 => "0001000010000100",
24947 => "0001000010000100",
24948 => "0001000010000100",
24949 => "0001000010001000",
24950 => "0001000010001000",
24951 => "0001000010001000",
24952 => "0001000010001000",
24953 => "0001000010001100",
24954 => "0001000010001100",
24955 => "0001000010001100",
24956 => "0001000010001100",
24957 => "0001000010001100",
24958 => "0001000010010000",
24959 => "0001000010010000",
24960 => "0001000010010000",
24961 => "0001000010010000",
24962 => "0001000010010100",
24963 => "0001000010010100",
24964 => "0001000010010100",
24965 => "0001000010010100",
24966 => "0001000010011000",
24967 => "0001000010011000",
24968 => "0001000010011000",
24969 => "0001000010011000",
24970 => "0001000010011000",
24971 => "0001000010011100",
24972 => "0001000010011100",
24973 => "0001000010011100",
24974 => "0001000010011100",
24975 => "0001000010100000",
24976 => "0001000010100000",
24977 => "0001000010100000",
24978 => "0001000010100000",
24979 => "0001000010100000",
24980 => "0001000010100100",
24981 => "0001000010100100",
24982 => "0001000010100100",
24983 => "0001000010100100",
24984 => "0001000010101000",
24985 => "0001000010101000",
24986 => "0001000010101000",
24987 => "0001000010101000",
24988 => "0001000010101000",
24989 => "0001000010101100",
24990 => "0001000010101100",
24991 => "0001000010101100",
24992 => "0001000010101100",
24993 => "0001000010110000",
24994 => "0001000010110000",
24995 => "0001000010110000",
24996 => "0001000010110000",
24997 => "0001000010110100",
24998 => "0001000010110100",
24999 => "0001000010110100",
25000 => "0001000010110100",
25001 => "0001000010110100",
25002 => "0001000010111000",
25003 => "0001000010111000",
25004 => "0001000010111000",
25005 => "0001000010111000",
25006 => "0001000010111100",
25007 => "0001000010111100",
25008 => "0001000010111100",
25009 => "0001000010111100",
25010 => "0001000010111100",
25011 => "0001000011000000",
25012 => "0001000011000000",
25013 => "0001000011000000",
25014 => "0001000011000000",
25015 => "0001000011000100",
25016 => "0001000011000100",
25017 => "0001000011000100",
25018 => "0001000011000100",
25019 => "0001000011001000",
25020 => "0001000011001000",
25021 => "0001000011001000",
25022 => "0001000011001000",
25023 => "0001000011001000",
25024 => "0001000011001100",
25025 => "0001000011001100",
25026 => "0001000011001100",
25027 => "0001000011001100",
25028 => "0001000011010000",
25029 => "0001000011010000",
25030 => "0001000011010000",
25031 => "0001000011010000",
25032 => "0001000011010000",
25033 => "0001000011010100",
25034 => "0001000011010100",
25035 => "0001000011010100",
25036 => "0001000011010100",
25037 => "0001000011011000",
25038 => "0001000011011000",
25039 => "0001000011011000",
25040 => "0001000011011000",
25041 => "0001000011011100",
25042 => "0001000011011100",
25043 => "0001000011011100",
25044 => "0001000011011100",
25045 => "0001000011011100",
25046 => "0001000011100000",
25047 => "0001000011100000",
25048 => "0001000011100000",
25049 => "0001000011100000",
25050 => "0001000011100100",
25051 => "0001000011100100",
25052 => "0001000011100100",
25053 => "0001000011100100",
25054 => "0001000011101000",
25055 => "0001000011101000",
25056 => "0001000011101000",
25057 => "0001000011101000",
25058 => "0001000011101000",
25059 => "0001000011101100",
25060 => "0001000011101100",
25061 => "0001000011101100",
25062 => "0001000011101100",
25063 => "0001000011110000",
25064 => "0001000011110000",
25065 => "0001000011110000",
25066 => "0001000011110000",
25067 => "0001000011110000",
25068 => "0001000011110100",
25069 => "0001000011110100",
25070 => "0001000011110100",
25071 => "0001000011110100",
25072 => "0001000011111000",
25073 => "0001000011111000",
25074 => "0001000011111000",
25075 => "0001000011111000",
25076 => "0001000011111100",
25077 => "0001000011111100",
25078 => "0001000011111100",
25079 => "0001000011111100",
25080 => "0001000011111100",
25081 => "0001000100000000",
25082 => "0001000100000000",
25083 => "0001000100000000",
25084 => "0001000100000000",
25085 => "0001000100000100",
25086 => "0001000100000100",
25087 => "0001000100000100",
25088 => "0001000100000100",
25089 => "0001000100001000",
25090 => "0001000100001000",
25091 => "0001000100001000",
25092 => "0001000100001000",
25093 => "0001000100001000",
25094 => "0001000100001100",
25095 => "0001000100001100",
25096 => "0001000100001100",
25097 => "0001000100001100",
25098 => "0001000100010000",
25099 => "0001000100010000",
25100 => "0001000100010000",
25101 => "0001000100010000",
25102 => "0001000100010100",
25103 => "0001000100010100",
25104 => "0001000100010100",
25105 => "0001000100010100",
25106 => "0001000100010100",
25107 => "0001000100011000",
25108 => "0001000100011000",
25109 => "0001000100011000",
25110 => "0001000100011000",
25111 => "0001000100011100",
25112 => "0001000100011100",
25113 => "0001000100011100",
25114 => "0001000100011100",
25115 => "0001000100100000",
25116 => "0001000100100000",
25117 => "0001000100100000",
25118 => "0001000100100000",
25119 => "0001000100100000",
25120 => "0001000100100100",
25121 => "0001000100100100",
25122 => "0001000100100100",
25123 => "0001000100100100",
25124 => "0001000100101000",
25125 => "0001000100101000",
25126 => "0001000100101000",
25127 => "0001000100101000",
25128 => "0001000100101100",
25129 => "0001000100101100",
25130 => "0001000100101100",
25131 => "0001000100101100",
25132 => "0001000100110000",
25133 => "0001000100110000",
25134 => "0001000100110000",
25135 => "0001000100110000",
25136 => "0001000100110000",
25137 => "0001000100110100",
25138 => "0001000100110100",
25139 => "0001000100110100",
25140 => "0001000100110100",
25141 => "0001000100111000",
25142 => "0001000100111000",
25143 => "0001000100111000",
25144 => "0001000100111000",
25145 => "0001000100111100",
25146 => "0001000100111100",
25147 => "0001000100111100",
25148 => "0001000100111100",
25149 => "0001000100111100",
25150 => "0001000101000000",
25151 => "0001000101000000",
25152 => "0001000101000000",
25153 => "0001000101000000",
25154 => "0001000101000100",
25155 => "0001000101000100",
25156 => "0001000101000100",
25157 => "0001000101000100",
25158 => "0001000101001000",
25159 => "0001000101001000",
25160 => "0001000101001000",
25161 => "0001000101001000",
25162 => "0001000101001100",
25163 => "0001000101001100",
25164 => "0001000101001100",
25165 => "0001000101001100",
25166 => "0001000101001100",
25167 => "0001000101010000",
25168 => "0001000101010000",
25169 => "0001000101010000",
25170 => "0001000101010000",
25171 => "0001000101010100",
25172 => "0001000101010100",
25173 => "0001000101010100",
25174 => "0001000101010100",
25175 => "0001000101011000",
25176 => "0001000101011000",
25177 => "0001000101011000",
25178 => "0001000101011000",
25179 => "0001000101011000",
25180 => "0001000101011100",
25181 => "0001000101011100",
25182 => "0001000101011100",
25183 => "0001000101011100",
25184 => "0001000101100000",
25185 => "0001000101100000",
25186 => "0001000101100000",
25187 => "0001000101100000",
25188 => "0001000101100100",
25189 => "0001000101100100",
25190 => "0001000101100100",
25191 => "0001000101100100",
25192 => "0001000101101000",
25193 => "0001000101101000",
25194 => "0001000101101000",
25195 => "0001000101101000",
25196 => "0001000101101000",
25197 => "0001000101101100",
25198 => "0001000101101100",
25199 => "0001000101101100",
25200 => "0001000101101100",
25201 => "0001000101110000",
25202 => "0001000101110000",
25203 => "0001000101110000",
25204 => "0001000101110000",
25205 => "0001000101110100",
25206 => "0001000101110100",
25207 => "0001000101110100",
25208 => "0001000101110100",
25209 => "0001000101111000",
25210 => "0001000101111000",
25211 => "0001000101111000",
25212 => "0001000101111000",
25213 => "0001000101111000",
25214 => "0001000101111100",
25215 => "0001000101111100",
25216 => "0001000101111100",
25217 => "0001000101111100",
25218 => "0001000110000000",
25219 => "0001000110000000",
25220 => "0001000110000000",
25221 => "0001000110000000",
25222 => "0001000110000100",
25223 => "0001000110000100",
25224 => "0001000110000100",
25225 => "0001000110000100",
25226 => "0001000110001000",
25227 => "0001000110001000",
25228 => "0001000110001000",
25229 => "0001000110001000",
25230 => "0001000110001000",
25231 => "0001000110001100",
25232 => "0001000110001100",
25233 => "0001000110001100",
25234 => "0001000110001100",
25235 => "0001000110010000",
25236 => "0001000110010000",
25237 => "0001000110010000",
25238 => "0001000110010000",
25239 => "0001000110010100",
25240 => "0001000110010100",
25241 => "0001000110010100",
25242 => "0001000110010100",
25243 => "0001000110011000",
25244 => "0001000110011000",
25245 => "0001000110011000",
25246 => "0001000110011000",
25247 => "0001000110011100",
25248 => "0001000110011100",
25249 => "0001000110011100",
25250 => "0001000110011100",
25251 => "0001000110011100",
25252 => "0001000110100000",
25253 => "0001000110100000",
25254 => "0001000110100000",
25255 => "0001000110100000",
25256 => "0001000110100100",
25257 => "0001000110100100",
25258 => "0001000110100100",
25259 => "0001000110100100",
25260 => "0001000110101000",
25261 => "0001000110101000",
25262 => "0001000110101000",
25263 => "0001000110101000",
25264 => "0001000110101100",
25265 => "0001000110101100",
25266 => "0001000110101100",
25267 => "0001000110101100",
25268 => "0001000110110000",
25269 => "0001000110110000",
25270 => "0001000110110000",
25271 => "0001000110110000",
25272 => "0001000110110000",
25273 => "0001000110110100",
25274 => "0001000110110100",
25275 => "0001000110110100",
25276 => "0001000110110100",
25277 => "0001000110111000",
25278 => "0001000110111000",
25279 => "0001000110111000",
25280 => "0001000110111000",
25281 => "0001000110111100",
25282 => "0001000110111100",
25283 => "0001000110111100",
25284 => "0001000110111100",
25285 => "0001000111000000",
25286 => "0001000111000000",
25287 => "0001000111000000",
25288 => "0001000111000000",
25289 => "0001000111000100",
25290 => "0001000111000100",
25291 => "0001000111000100",
25292 => "0001000111000100",
25293 => "0001000111000100",
25294 => "0001000111001000",
25295 => "0001000111001000",
25296 => "0001000111001000",
25297 => "0001000111001000",
25298 => "0001000111001100",
25299 => "0001000111001100",
25300 => "0001000111001100",
25301 => "0001000111001100",
25302 => "0001000111010000",
25303 => "0001000111010000",
25304 => "0001000111010000",
25305 => "0001000111010000",
25306 => "0001000111010100",
25307 => "0001000111010100",
25308 => "0001000111010100",
25309 => "0001000111010100",
25310 => "0001000111011000",
25311 => "0001000111011000",
25312 => "0001000111011000",
25313 => "0001000111011000",
25314 => "0001000111011100",
25315 => "0001000111011100",
25316 => "0001000111011100",
25317 => "0001000111011100",
25318 => "0001000111011100",
25319 => "0001000111100000",
25320 => "0001000111100000",
25321 => "0001000111100000",
25322 => "0001000111100000",
25323 => "0001000111100100",
25324 => "0001000111100100",
25325 => "0001000111100100",
25326 => "0001000111100100",
25327 => "0001000111101000",
25328 => "0001000111101000",
25329 => "0001000111101000",
25330 => "0001000111101000",
25331 => "0001000111101100",
25332 => "0001000111101100",
25333 => "0001000111101100",
25334 => "0001000111101100",
25335 => "0001000111110000",
25336 => "0001000111110000",
25337 => "0001000111110000",
25338 => "0001000111110000",
25339 => "0001000111110100",
25340 => "0001000111110100",
25341 => "0001000111110100",
25342 => "0001000111110100",
25343 => "0001000111110100",
25344 => "0001000111111000",
25345 => "0001000111111000",
25346 => "0001000111111000",
25347 => "0001000111111000",
25348 => "0001000111111100",
25349 => "0001000111111100",
25350 => "0001000111111100",
25351 => "0001000111111100",
25352 => "0001001000000000",
25353 => "0001001000000000",
25354 => "0001001000000000",
25355 => "0001001000000000",
25356 => "0001001000000100",
25357 => "0001001000000100",
25358 => "0001001000000100",
25359 => "0001001000000100",
25360 => "0001001000001000",
25361 => "0001001000001000",
25362 => "0001001000001000",
25363 => "0001001000001000",
25364 => "0001001000001100",
25365 => "0001001000001100",
25366 => "0001001000001100",
25367 => "0001001000001100",
25368 => "0001001000010000",
25369 => "0001001000010000",
25370 => "0001001000010000",
25371 => "0001001000010000",
25372 => "0001001000010100",
25373 => "0001001000010100",
25374 => "0001001000010100",
25375 => "0001001000010100",
25376 => "0001001000010100",
25377 => "0001001000011000",
25378 => "0001001000011000",
25379 => "0001001000011000",
25380 => "0001001000011000",
25381 => "0001001000011100",
25382 => "0001001000011100",
25383 => "0001001000011100",
25384 => "0001001000011100",
25385 => "0001001000100000",
25386 => "0001001000100000",
25387 => "0001001000100000",
25388 => "0001001000100000",
25389 => "0001001000100100",
25390 => "0001001000100100",
25391 => "0001001000100100",
25392 => "0001001000100100",
25393 => "0001001000101000",
25394 => "0001001000101000",
25395 => "0001001000101000",
25396 => "0001001000101000",
25397 => "0001001000101100",
25398 => "0001001000101100",
25399 => "0001001000101100",
25400 => "0001001000101100",
25401 => "0001001000110000",
25402 => "0001001000110000",
25403 => "0001001000110000",
25404 => "0001001000110000",
25405 => "0001001000110100",
25406 => "0001001000110100",
25407 => "0001001000110100",
25408 => "0001001000110100",
25409 => "0001001000111000",
25410 => "0001001000111000",
25411 => "0001001000111000",
25412 => "0001001000111000",
25413 => "0001001000111000",
25414 => "0001001000111100",
25415 => "0001001000111100",
25416 => "0001001000111100",
25417 => "0001001000111100",
25418 => "0001001001000000",
25419 => "0001001001000000",
25420 => "0001001001000000",
25421 => "0001001001000000",
25422 => "0001001001000100",
25423 => "0001001001000100",
25424 => "0001001001000100",
25425 => "0001001001000100",
25426 => "0001001001001000",
25427 => "0001001001001000",
25428 => "0001001001001000",
25429 => "0001001001001000",
25430 => "0001001001001100",
25431 => "0001001001001100",
25432 => "0001001001001100",
25433 => "0001001001001100",
25434 => "0001001001010000",
25435 => "0001001001010000",
25436 => "0001001001010000",
25437 => "0001001001010000",
25438 => "0001001001010100",
25439 => "0001001001010100",
25440 => "0001001001010100",
25441 => "0001001001010100",
25442 => "0001001001011000",
25443 => "0001001001011000",
25444 => "0001001001011000",
25445 => "0001001001011000",
25446 => "0001001001011100",
25447 => "0001001001011100",
25448 => "0001001001011100",
25449 => "0001001001011100",
25450 => "0001001001100000",
25451 => "0001001001100000",
25452 => "0001001001100000",
25453 => "0001001001100000",
25454 => "0001001001100100",
25455 => "0001001001100100",
25456 => "0001001001100100",
25457 => "0001001001100100",
25458 => "0001001001101000",
25459 => "0001001001101000",
25460 => "0001001001101000",
25461 => "0001001001101000",
25462 => "0001001001101000",
25463 => "0001001001101100",
25464 => "0001001001101100",
25465 => "0001001001101100",
25466 => "0001001001101100",
25467 => "0001001001110000",
25468 => "0001001001110000",
25469 => "0001001001110000",
25470 => "0001001001110000",
25471 => "0001001001110100",
25472 => "0001001001110100",
25473 => "0001001001110100",
25474 => "0001001001110100",
25475 => "0001001001111000",
25476 => "0001001001111000",
25477 => "0001001001111000",
25478 => "0001001001111000",
25479 => "0001001001111100",
25480 => "0001001001111100",
25481 => "0001001001111100",
25482 => "0001001001111100",
25483 => "0001001010000000",
25484 => "0001001010000000",
25485 => "0001001010000000",
25486 => "0001001010000000",
25487 => "0001001010000100",
25488 => "0001001010000100",
25489 => "0001001010000100",
25490 => "0001001010000100",
25491 => "0001001010001000",
25492 => "0001001010001000",
25493 => "0001001010001000",
25494 => "0001001010001000",
25495 => "0001001010001100",
25496 => "0001001010001100",
25497 => "0001001010001100",
25498 => "0001001010001100",
25499 => "0001001010010000",
25500 => "0001001010010000",
25501 => "0001001010010000",
25502 => "0001001010010000",
25503 => "0001001010010100",
25504 => "0001001010010100",
25505 => "0001001010010100",
25506 => "0001001010010100",
25507 => "0001001010011000",
25508 => "0001001010011000",
25509 => "0001001010011000",
25510 => "0001001010011000",
25511 => "0001001010011100",
25512 => "0001001010011100",
25513 => "0001001010011100",
25514 => "0001001010011100",
25515 => "0001001010100000",
25516 => "0001001010100000",
25517 => "0001001010100000",
25518 => "0001001010100000",
25519 => "0001001010100100",
25520 => "0001001010100100",
25521 => "0001001010100100",
25522 => "0001001010100100",
25523 => "0001001010101000",
25524 => "0001001010101000",
25525 => "0001001010101000",
25526 => "0001001010101000",
25527 => "0001001010101100",
25528 => "0001001010101100",
25529 => "0001001010101100",
25530 => "0001001010101100",
25531 => "0001001010110000",
25532 => "0001001010110000",
25533 => "0001001010110000",
25534 => "0001001010110000",
25535 => "0001001010110100",
25536 => "0001001010110100",
25537 => "0001001010110100",
25538 => "0001001010110100",
25539 => "0001001010111000",
25540 => "0001001010111000",
25541 => "0001001010111000",
25542 => "0001001010111000",
25543 => "0001001010111100",
25544 => "0001001010111100",
25545 => "0001001010111100",
25546 => "0001001010111100",
25547 => "0001001011000000",
25548 => "0001001011000000",
25549 => "0001001011000000",
25550 => "0001001011000000",
25551 => "0001001011000100",
25552 => "0001001011000100",
25553 => "0001001011000100",
25554 => "0001001011000100",
25555 => "0001001011001000",
25556 => "0001001011001000",
25557 => "0001001011001000",
25558 => "0001001011001000",
25559 => "0001001011001100",
25560 => "0001001011001100",
25561 => "0001001011001100",
25562 => "0001001011001100",
25563 => "0001001011010000",
25564 => "0001001011010000",
25565 => "0001001011010000",
25566 => "0001001011010000",
25567 => "0001001011010100",
25568 => "0001001011010100",
25569 => "0001001011010100",
25570 => "0001001011010100",
25571 => "0001001011011000",
25572 => "0001001011011000",
25573 => "0001001011011000",
25574 => "0001001011011000",
25575 => "0001001011011100",
25576 => "0001001011011100",
25577 => "0001001011011100",
25578 => "0001001011011100",
25579 => "0001001011100000",
25580 => "0001001011100000",
25581 => "0001001011100000",
25582 => "0001001011100000",
25583 => "0001001011100100",
25584 => "0001001011100100",
25585 => "0001001011100100",
25586 => "0001001011100100",
25587 => "0001001011101000",
25588 => "0001001011101000",
25589 => "0001001011101000",
25590 => "0001001011101000",
25591 => "0001001011101100",
25592 => "0001001011101100",
25593 => "0001001011101100",
25594 => "0001001011101100",
25595 => "0001001011110000",
25596 => "0001001011110000",
25597 => "0001001011110000",
25598 => "0001001011110000",
25599 => "0001001011110100",
25600 => "0001001011110100",
25601 => "0001001011110100",
25602 => "0001001011110100",
25603 => "0001001011111000",
25604 => "0001001011111000",
25605 => "0001001011111000",
25606 => "0001001011111000",
25607 => "0001001011111100",
25608 => "0001001011111100",
25609 => "0001001011111100",
25610 => "0001001011111100",
25611 => "0001001100000000",
25612 => "0001001100000000",
25613 => "0001001100000000",
25614 => "0001001100000000",
25615 => "0001001100000100",
25616 => "0001001100000100",
25617 => "0001001100000100",
25618 => "0001001100000100",
25619 => "0001001100001000",
25620 => "0001001100001000",
25621 => "0001001100001000",
25622 => "0001001100001000",
25623 => "0001001100001100",
25624 => "0001001100001100",
25625 => "0001001100001100",
25626 => "0001001100001100",
25627 => "0001001100010000",
25628 => "0001001100010000",
25629 => "0001001100010000",
25630 => "0001001100010000",
25631 => "0001001100010100",
25632 => "0001001100010100",
25633 => "0001001100010100",
25634 => "0001001100011000",
25635 => "0001001100011000",
25636 => "0001001100011000",
25637 => "0001001100011000",
25638 => "0001001100011100",
25639 => "0001001100011100",
25640 => "0001001100011100",
25641 => "0001001100011100",
25642 => "0001001100100000",
25643 => "0001001100100000",
25644 => "0001001100100000",
25645 => "0001001100100000",
25646 => "0001001100100100",
25647 => "0001001100100100",
25648 => "0001001100100100",
25649 => "0001001100100100",
25650 => "0001001100101000",
25651 => "0001001100101000",
25652 => "0001001100101000",
25653 => "0001001100101000",
25654 => "0001001100101100",
25655 => "0001001100101100",
25656 => "0001001100101100",
25657 => "0001001100101100",
25658 => "0001001100110000",
25659 => "0001001100110000",
25660 => "0001001100110000",
25661 => "0001001100110000",
25662 => "0001001100110100",
25663 => "0001001100110100",
25664 => "0001001100110100",
25665 => "0001001100110100",
25666 => "0001001100111000",
25667 => "0001001100111000",
25668 => "0001001100111000",
25669 => "0001001100111000",
25670 => "0001001100111100",
25671 => "0001001100111100",
25672 => "0001001100111100",
25673 => "0001001100111100",
25674 => "0001001101000000",
25675 => "0001001101000000",
25676 => "0001001101000000",
25677 => "0001001101000000",
25678 => "0001001101000100",
25679 => "0001001101000100",
25680 => "0001001101000100",
25681 => "0001001101000100",
25682 => "0001001101001000",
25683 => "0001001101001000",
25684 => "0001001101001000",
25685 => "0001001101001100",
25686 => "0001001101001100",
25687 => "0001001101001100",
25688 => "0001001101001100",
25689 => "0001001101010000",
25690 => "0001001101010000",
25691 => "0001001101010000",
25692 => "0001001101010000",
25693 => "0001001101010100",
25694 => "0001001101010100",
25695 => "0001001101010100",
25696 => "0001001101010100",
25697 => "0001001101011000",
25698 => "0001001101011000",
25699 => "0001001101011000",
25700 => "0001001101011000",
25701 => "0001001101011100",
25702 => "0001001101011100",
25703 => "0001001101011100",
25704 => "0001001101011100",
25705 => "0001001101100000",
25706 => "0001001101100000",
25707 => "0001001101100000",
25708 => "0001001101100000",
25709 => "0001001101100100",
25710 => "0001001101100100",
25711 => "0001001101100100",
25712 => "0001001101100100",
25713 => "0001001101101000",
25714 => "0001001101101000",
25715 => "0001001101101000",
25716 => "0001001101101000",
25717 => "0001001101101100",
25718 => "0001001101101100",
25719 => "0001001101101100",
25720 => "0001001101101100",
25721 => "0001001101110000",
25722 => "0001001101110000",
25723 => "0001001101110000",
25724 => "0001001101110100",
25725 => "0001001101110100",
25726 => "0001001101110100",
25727 => "0001001101110100",
25728 => "0001001101111000",
25729 => "0001001101111000",
25730 => "0001001101111000",
25731 => "0001001101111000",
25732 => "0001001101111100",
25733 => "0001001101111100",
25734 => "0001001101111100",
25735 => "0001001101111100",
25736 => "0001001110000000",
25737 => "0001001110000000",
25738 => "0001001110000000",
25739 => "0001001110000000",
25740 => "0001001110000100",
25741 => "0001001110000100",
25742 => "0001001110000100",
25743 => "0001001110000100",
25744 => "0001001110001000",
25745 => "0001001110001000",
25746 => "0001001110001000",
25747 => "0001001110001000",
25748 => "0001001110001100",
25749 => "0001001110001100",
25750 => "0001001110001100",
25751 => "0001001110001100",
25752 => "0001001110010000",
25753 => "0001001110010000",
25754 => "0001001110010000",
25755 => "0001001110010100",
25756 => "0001001110010100",
25757 => "0001001110010100",
25758 => "0001001110010100",
25759 => "0001001110011000",
25760 => "0001001110011000",
25761 => "0001001110011000",
25762 => "0001001110011000",
25763 => "0001001110011100",
25764 => "0001001110011100",
25765 => "0001001110011100",
25766 => "0001001110011100",
25767 => "0001001110100000",
25768 => "0001001110100000",
25769 => "0001001110100000",
25770 => "0001001110100000",
25771 => "0001001110100100",
25772 => "0001001110100100",
25773 => "0001001110100100",
25774 => "0001001110100100",
25775 => "0001001110101000",
25776 => "0001001110101000",
25777 => "0001001110101000",
25778 => "0001001110101000",
25779 => "0001001110101100",
25780 => "0001001110101100",
25781 => "0001001110101100",
25782 => "0001001110110000",
25783 => "0001001110110000",
25784 => "0001001110110000",
25785 => "0001001110110000",
25786 => "0001001110110100",
25787 => "0001001110110100",
25788 => "0001001110110100",
25789 => "0001001110110100",
25790 => "0001001110111000",
25791 => "0001001110111000",
25792 => "0001001110111000",
25793 => "0001001110111000",
25794 => "0001001110111100",
25795 => "0001001110111100",
25796 => "0001001110111100",
25797 => "0001001110111100",
25798 => "0001001111000000",
25799 => "0001001111000000",
25800 => "0001001111000000",
25801 => "0001001111000000",
25802 => "0001001111000100",
25803 => "0001001111000100",
25804 => "0001001111000100",
25805 => "0001001111001000",
25806 => "0001001111001000",
25807 => "0001001111001000",
25808 => "0001001111001000",
25809 => "0001001111001100",
25810 => "0001001111001100",
25811 => "0001001111001100",
25812 => "0001001111001100",
25813 => "0001001111010000",
25814 => "0001001111010000",
25815 => "0001001111010000",
25816 => "0001001111010000",
25817 => "0001001111010100",
25818 => "0001001111010100",
25819 => "0001001111010100",
25820 => "0001001111010100",
25821 => "0001001111011000",
25822 => "0001001111011000",
25823 => "0001001111011000",
25824 => "0001001111011100",
25825 => "0001001111011100",
25826 => "0001001111011100",
25827 => "0001001111011100",
25828 => "0001001111100000",
25829 => "0001001111100000",
25830 => "0001001111100000",
25831 => "0001001111100000",
25832 => "0001001111100100",
25833 => "0001001111100100",
25834 => "0001001111100100",
25835 => "0001001111100100",
25836 => "0001001111101000",
25837 => "0001001111101000",
25838 => "0001001111101000",
25839 => "0001001111101000",
25840 => "0001001111101100",
25841 => "0001001111101100",
25842 => "0001001111101100",
25843 => "0001001111101100",
25844 => "0001001111110000",
25845 => "0001001111110000",
25846 => "0001001111110000",
25847 => "0001001111110100",
25848 => "0001001111110100",
25849 => "0001001111110100",
25850 => "0001001111110100",
25851 => "0001001111111000",
25852 => "0001001111111000",
25853 => "0001001111111000",
25854 => "0001001111111000",
25855 => "0001001111111100",
25856 => "0001001111111100",
25857 => "0001001111111100",
25858 => "0001001111111100",
25859 => "0001010000000000",
25860 => "0001010000000000",
25861 => "0001010000000000",
25862 => "0001010000000000",
25863 => "0001010000000100",
25864 => "0001010000000100",
25865 => "0001010000000100",
25866 => "0001010000001000",
25867 => "0001010000001000",
25868 => "0001010000001000",
25869 => "0001010000001000",
25870 => "0001010000001100",
25871 => "0001010000001100",
25872 => "0001010000001100",
25873 => "0001010000001100",
25874 => "0001010000010000",
25875 => "0001010000010000",
25876 => "0001010000010000",
25877 => "0001010000010000",
25878 => "0001010000010100",
25879 => "0001010000010100",
25880 => "0001010000010100",
25881 => "0001010000011000",
25882 => "0001010000011000",
25883 => "0001010000011000",
25884 => "0001010000011000",
25885 => "0001010000011100",
25886 => "0001010000011100",
25887 => "0001010000011100",
25888 => "0001010000011100",
25889 => "0001010000100000",
25890 => "0001010000100000",
25891 => "0001010000100000",
25892 => "0001010000100000",
25893 => "0001010000100100",
25894 => "0001010000100100",
25895 => "0001010000100100",
25896 => "0001010000100100",
25897 => "0001010000101000",
25898 => "0001010000101000",
25899 => "0001010000101000",
25900 => "0001010000101100",
25901 => "0001010000101100",
25902 => "0001010000101100",
25903 => "0001010000101100",
25904 => "0001010000110000",
25905 => "0001010000110000",
25906 => "0001010000110000",
25907 => "0001010000110000",
25908 => "0001010000110100",
25909 => "0001010000110100",
25910 => "0001010000110100",
25911 => "0001010000110100",
25912 => "0001010000111000",
25913 => "0001010000111000",
25914 => "0001010000111000",
25915 => "0001010000111100",
25916 => "0001010000111100",
25917 => "0001010000111100",
25918 => "0001010000111100",
25919 => "0001010001000000",
25920 => "0001010001000000",
25921 => "0001010001000000",
25922 => "0001010001000000",
25923 => "0001010001000100",
25924 => "0001010001000100",
25925 => "0001010001000100",
25926 => "0001010001000100",
25927 => "0001010001001000",
25928 => "0001010001001000",
25929 => "0001010001001000",
25930 => "0001010001001100",
25931 => "0001010001001100",
25932 => "0001010001001100",
25933 => "0001010001001100",
25934 => "0001010001010000",
25935 => "0001010001010000",
25936 => "0001010001010000",
25937 => "0001010001010000",
25938 => "0001010001010100",
25939 => "0001010001010100",
25940 => "0001010001010100",
25941 => "0001010001010100",
25942 => "0001010001011000",
25943 => "0001010001011000",
25944 => "0001010001011000",
25945 => "0001010001011100",
25946 => "0001010001011100",
25947 => "0001010001011100",
25948 => "0001010001011100",
25949 => "0001010001100000",
25950 => "0001010001100000",
25951 => "0001010001100000",
25952 => "0001010001100000",
25953 => "0001010001100100",
25954 => "0001010001100100",
25955 => "0001010001100100",
25956 => "0001010001100100",
25957 => "0001010001101000",
25958 => "0001010001101000",
25959 => "0001010001101000",
25960 => "0001010001101100",
25961 => "0001010001101100",
25962 => "0001010001101100",
25963 => "0001010001101100",
25964 => "0001010001110000",
25965 => "0001010001110000",
25966 => "0001010001110000",
25967 => "0001010001110000",
25968 => "0001010001110100",
25969 => "0001010001110100",
25970 => "0001010001110100",
25971 => "0001010001111000",
25972 => "0001010001111000",
25973 => "0001010001111000",
25974 => "0001010001111000",
25975 => "0001010001111100",
25976 => "0001010001111100",
25977 => "0001010001111100",
25978 => "0001010001111100",
25979 => "0001010010000000",
25980 => "0001010010000000",
25981 => "0001010010000000",
25982 => "0001010010000000",
25983 => "0001010010000100",
25984 => "0001010010000100",
25985 => "0001010010000100",
25986 => "0001010010001000",
25987 => "0001010010001000",
25988 => "0001010010001000",
25989 => "0001010010001000",
25990 => "0001010010001100",
25991 => "0001010010001100",
25992 => "0001010010001100",
25993 => "0001010010001100",
25994 => "0001010010010000",
25995 => "0001010010010000",
25996 => "0001010010010000",
25997 => "0001010010010100",
25998 => "0001010010010100",
25999 => "0001010010010100",
26000 => "0001010010010100",
26001 => "0001010010011000",
26002 => "0001010010011000",
26003 => "0001010010011000",
26004 => "0001010010011000",
26005 => "0001010010011100",
26006 => "0001010010011100",
26007 => "0001010010011100",
26008 => "0001010010011100",
26009 => "0001010010100000",
26010 => "0001010010100000",
26011 => "0001010010100000",
26012 => "0001010010100100",
26013 => "0001010010100100",
26014 => "0001010010100100",
26015 => "0001010010100100",
26016 => "0001010010101000",
26017 => "0001010010101000",
26018 => "0001010010101000",
26019 => "0001010010101000",
26020 => "0001010010101100",
26021 => "0001010010101100",
26022 => "0001010010101100",
26023 => "0001010010110000",
26024 => "0001010010110000",
26025 => "0001010010110000",
26026 => "0001010010110000",
26027 => "0001010010110100",
26028 => "0001010010110100",
26029 => "0001010010110100",
26030 => "0001010010110100",
26031 => "0001010010111000",
26032 => "0001010010111000",
26033 => "0001010010111000",
26034 => "0001010010111100",
26035 => "0001010010111100",
26036 => "0001010010111100",
26037 => "0001010010111100",
26038 => "0001010011000000",
26039 => "0001010011000000",
26040 => "0001010011000000",
26041 => "0001010011000000",
26042 => "0001010011000100",
26043 => "0001010011000100",
26044 => "0001010011000100",
26045 => "0001010011001000",
26046 => "0001010011001000",
26047 => "0001010011001000",
26048 => "0001010011001000",
26049 => "0001010011001100",
26050 => "0001010011001100",
26051 => "0001010011001100",
26052 => "0001010011001100",
26053 => "0001010011010000",
26054 => "0001010011010000",
26055 => "0001010011010000",
26056 => "0001010011010100",
26057 => "0001010011010100",
26058 => "0001010011010100",
26059 => "0001010011010100",
26060 => "0001010011011000",
26061 => "0001010011011000",
26062 => "0001010011011000",
26063 => "0001010011011000",
26064 => "0001010011011100",
26065 => "0001010011011100",
26066 => "0001010011011100",
26067 => "0001010011100000",
26068 => "0001010011100000",
26069 => "0001010011100000",
26070 => "0001010011100000",
26071 => "0001010011100100",
26072 => "0001010011100100",
26073 => "0001010011100100",
26074 => "0001010011100100",
26075 => "0001010011101000",
26076 => "0001010011101000",
26077 => "0001010011101000",
26078 => "0001010011101100",
26079 => "0001010011101100",
26080 => "0001010011101100",
26081 => "0001010011101100",
26082 => "0001010011110000",
26083 => "0001010011110000",
26084 => "0001010011110000",
26085 => "0001010011110000",
26086 => "0001010011110100",
26087 => "0001010011110100",
26088 => "0001010011110100",
26089 => "0001010011111000",
26090 => "0001010011111000",
26091 => "0001010011111000",
26092 => "0001010011111000",
26093 => "0001010011111100",
26094 => "0001010011111100",
26095 => "0001010011111100",
26096 => "0001010011111100",
26097 => "0001010100000000",
26098 => "0001010100000000",
26099 => "0001010100000000",
26100 => "0001010100000100",
26101 => "0001010100000100",
26102 => "0001010100000100",
26103 => "0001010100000100",
26104 => "0001010100001000",
26105 => "0001010100001000",
26106 => "0001010100001000",
26107 => "0001010100001000",
26108 => "0001010100001100",
26109 => "0001010100001100",
26110 => "0001010100001100",
26111 => "0001010100010000",
26112 => "0001010100010000",
26113 => "0001010100010000",
26114 => "0001010100010000",
26115 => "0001010100010100",
26116 => "0001010100010100",
26117 => "0001010100010100",
26118 => "0001010100010100",
26119 => "0001010100011000",
26120 => "0001010100011000",
26121 => "0001010100011000",
26122 => "0001010100011100",
26123 => "0001010100011100",
26124 => "0001010100011100",
26125 => "0001010100011100",
26126 => "0001010100100000",
26127 => "0001010100100000",
26128 => "0001010100100000",
26129 => "0001010100100100",
26130 => "0001010100100100",
26131 => "0001010100100100",
26132 => "0001010100100100",
26133 => "0001010100101000",
26134 => "0001010100101000",
26135 => "0001010100101000",
26136 => "0001010100101000",
26137 => "0001010100101100",
26138 => "0001010100101100",
26139 => "0001010100101100",
26140 => "0001010100110000",
26141 => "0001010100110000",
26142 => "0001010100110000",
26143 => "0001010100110000",
26144 => "0001010100110100",
26145 => "0001010100110100",
26146 => "0001010100110100",
26147 => "0001010100110100",
26148 => "0001010100111000",
26149 => "0001010100111000",
26150 => "0001010100111000",
26151 => "0001010100111100",
26152 => "0001010100111100",
26153 => "0001010100111100",
26154 => "0001010100111100",
26155 => "0001010101000000",
26156 => "0001010101000000",
26157 => "0001010101000000",
26158 => "0001010101000100",
26159 => "0001010101000100",
26160 => "0001010101000100",
26161 => "0001010101000100",
26162 => "0001010101001000",
26163 => "0001010101001000",
26164 => "0001010101001000",
26165 => "0001010101001000",
26166 => "0001010101001100",
26167 => "0001010101001100",
26168 => "0001010101001100",
26169 => "0001010101010000",
26170 => "0001010101010000",
26171 => "0001010101010000",
26172 => "0001010101010000",
26173 => "0001010101010100",
26174 => "0001010101010100",
26175 => "0001010101010100",
26176 => "0001010101011000",
26177 => "0001010101011000",
26178 => "0001010101011000",
26179 => "0001010101011000",
26180 => "0001010101011100",
26181 => "0001010101011100",
26182 => "0001010101011100",
26183 => "0001010101011100",
26184 => "0001010101100000",
26185 => "0001010101100000",
26186 => "0001010101100000",
26187 => "0001010101100100",
26188 => "0001010101100100",
26189 => "0001010101100100",
26190 => "0001010101100100",
26191 => "0001010101101000",
26192 => "0001010101101000",
26193 => "0001010101101000",
26194 => "0001010101101100",
26195 => "0001010101101100",
26196 => "0001010101101100",
26197 => "0001010101101100",
26198 => "0001010101110000",
26199 => "0001010101110000",
26200 => "0001010101110000",
26201 => "0001010101110000",
26202 => "0001010101110100",
26203 => "0001010101110100",
26204 => "0001010101110100",
26205 => "0001010101111000",
26206 => "0001010101111000",
26207 => "0001010101111000",
26208 => "0001010101111000",
26209 => "0001010101111100",
26210 => "0001010101111100",
26211 => "0001010101111100",
26212 => "0001010110000000",
26213 => "0001010110000000",
26214 => "0001010110000000",
26215 => "0001010110000000",
26216 => "0001010110000100",
26217 => "0001010110000100",
26218 => "0001010110000100",
26219 => "0001010110001000",
26220 => "0001010110001000",
26221 => "0001010110001000",
26222 => "0001010110001000",
26223 => "0001010110001100",
26224 => "0001010110001100",
26225 => "0001010110001100",
26226 => "0001010110001100",
26227 => "0001010110010000",
26228 => "0001010110010000",
26229 => "0001010110010000",
26230 => "0001010110010100",
26231 => "0001010110010100",
26232 => "0001010110010100",
26233 => "0001010110010100",
26234 => "0001010110011000",
26235 => "0001010110011000",
26236 => "0001010110011000",
26237 => "0001010110011100",
26238 => "0001010110011100",
26239 => "0001010110011100",
26240 => "0001010110011100",
26241 => "0001010110100000",
26242 => "0001010110100000",
26243 => "0001010110100000",
26244 => "0001010110100100",
26245 => "0001010110100100",
26246 => "0001010110100100",
26247 => "0001010110100100",
26248 => "0001010110101000",
26249 => "0001010110101000",
26250 => "0001010110101000",
26251 => "0001010110101000",
26252 => "0001010110101100",
26253 => "0001010110101100",
26254 => "0001010110101100",
26255 => "0001010110110000",
26256 => "0001010110110000",
26257 => "0001010110110000",
26258 => "0001010110110000",
26259 => "0001010110110100",
26260 => "0001010110110100",
26261 => "0001010110110100",
26262 => "0001010110111000",
26263 => "0001010110111000",
26264 => "0001010110111000",
26265 => "0001010110111000",
26266 => "0001010110111100",
26267 => "0001010110111100",
26268 => "0001010110111100",
26269 => "0001010111000000",
26270 => "0001010111000000",
26271 => "0001010111000000",
26272 => "0001010111000000",
26273 => "0001010111000100",
26274 => "0001010111000100",
26275 => "0001010111000100",
26276 => "0001010111001000",
26277 => "0001010111001000",
26278 => "0001010111001000",
26279 => "0001010111001000",
26280 => "0001010111001100",
26281 => "0001010111001100",
26282 => "0001010111001100",
26283 => "0001010111010000",
26284 => "0001010111010000",
26285 => "0001010111010000",
26286 => "0001010111010000",
26287 => "0001010111010100",
26288 => "0001010111010100",
26289 => "0001010111010100",
26290 => "0001010111010100",
26291 => "0001010111011000",
26292 => "0001010111011000",
26293 => "0001010111011000",
26294 => "0001010111011100",
26295 => "0001010111011100",
26296 => "0001010111011100",
26297 => "0001010111011100",
26298 => "0001010111100000",
26299 => "0001010111100000",
26300 => "0001010111100000",
26301 => "0001010111100100",
26302 => "0001010111100100",
26303 => "0001010111100100",
26304 => "0001010111100100",
26305 => "0001010111101000",
26306 => "0001010111101000",
26307 => "0001010111101000",
26308 => "0001010111101100",
26309 => "0001010111101100",
26310 => "0001010111101100",
26311 => "0001010111101100",
26312 => "0001010111110000",
26313 => "0001010111110000",
26314 => "0001010111110000",
26315 => "0001010111110100",
26316 => "0001010111110100",
26317 => "0001010111110100",
26318 => "0001010111110100",
26319 => "0001010111111000",
26320 => "0001010111111000",
26321 => "0001010111111000",
26322 => "0001010111111100",
26323 => "0001010111111100",
26324 => "0001010111111100",
26325 => "0001010111111100",
26326 => "0001011000000000",
26327 => "0001011000000000",
26328 => "0001011000000000",
26329 => "0001011000000100",
26330 => "0001011000000100",
26331 => "0001011000000100",
26332 => "0001011000000100",
26333 => "0001011000001000",
26334 => "0001011000001000",
26335 => "0001011000001000",
26336 => "0001011000001100",
26337 => "0001011000001100",
26338 => "0001011000001100",
26339 => "0001011000001100",
26340 => "0001011000010000",
26341 => "0001011000010000",
26342 => "0001011000010000",
26343 => "0001011000010100",
26344 => "0001011000010100",
26345 => "0001011000010100",
26346 => "0001011000010100",
26347 => "0001011000011000",
26348 => "0001011000011000",
26349 => "0001011000011000",
26350 => "0001011000011100",
26351 => "0001011000011100",
26352 => "0001011000011100",
26353 => "0001011000011100",
26354 => "0001011000100000",
26355 => "0001011000100000",
26356 => "0001011000100000",
26357 => "0001011000100100",
26358 => "0001011000100100",
26359 => "0001011000100100",
26360 => "0001011000100100",
26361 => "0001011000101000",
26362 => "0001011000101000",
26363 => "0001011000101000",
26364 => "0001011000101100",
26365 => "0001011000101100",
26366 => "0001011000101100",
26367 => "0001011000101100",
26368 => "0001011000110000",
26369 => "0001011000110000",
26370 => "0001011000110000",
26371 => "0001011000110100",
26372 => "0001011000110100",
26373 => "0001011000110100",
26374 => "0001011000110100",
26375 => "0001011000111000",
26376 => "0001011000111000",
26377 => "0001011000111000",
26378 => "0001011000111100",
26379 => "0001011000111100",
26380 => "0001011000111100",
26381 => "0001011000111100",
26382 => "0001011001000000",
26383 => "0001011001000000",
26384 => "0001011001000000",
26385 => "0001011001000100",
26386 => "0001011001000100",
26387 => "0001011001000100",
26388 => "0001011001000100",
26389 => "0001011001001000",
26390 => "0001011001001000",
26391 => "0001011001001000",
26392 => "0001011001001100",
26393 => "0001011001001100",
26394 => "0001011001001100",
26395 => "0001011001001100",
26396 => "0001011001010000",
26397 => "0001011001010000",
26398 => "0001011001010000",
26399 => "0001011001010100",
26400 => "0001011001010100",
26401 => "0001011001010100",
26402 => "0001011001010100",
26403 => "0001011001011000",
26404 => "0001011001011000",
26405 => "0001011001011000",
26406 => "0001011001011100",
26407 => "0001011001011100",
26408 => "0001011001011100",
26409 => "0001011001011100",
26410 => "0001011001100000",
26411 => "0001011001100000",
26412 => "0001011001100000",
26413 => "0001011001100100",
26414 => "0001011001100100",
26415 => "0001011001100100",
26416 => "0001011001100100",
26417 => "0001011001101000",
26418 => "0001011001101000",
26419 => "0001011001101000",
26420 => "0001011001101100",
26421 => "0001011001101100",
26422 => "0001011001101100",
26423 => "0001011001110000",
26424 => "0001011001110000",
26425 => "0001011001110000",
26426 => "0001011001110000",
26427 => "0001011001110100",
26428 => "0001011001110100",
26429 => "0001011001110100",
26430 => "0001011001111000",
26431 => "0001011001111000",
26432 => "0001011001111000",
26433 => "0001011001111000",
26434 => "0001011001111100",
26435 => "0001011001111100",
26436 => "0001011001111100",
26437 => "0001011010000000",
26438 => "0001011010000000",
26439 => "0001011010000000",
26440 => "0001011010000000",
26441 => "0001011010000100",
26442 => "0001011010000100",
26443 => "0001011010000100",
26444 => "0001011010001000",
26445 => "0001011010001000",
26446 => "0001011010001000",
26447 => "0001011010001000",
26448 => "0001011010001100",
26449 => "0001011010001100",
26450 => "0001011010001100",
26451 => "0001011010010000",
26452 => "0001011010010000",
26453 => "0001011010010000",
26454 => "0001011010010100",
26455 => "0001011010010100",
26456 => "0001011010010100",
26457 => "0001011010010100",
26458 => "0001011010011000",
26459 => "0001011010011000",
26460 => "0001011010011000",
26461 => "0001011010011100",
26462 => "0001011010011100",
26463 => "0001011010011100",
26464 => "0001011010011100",
26465 => "0001011010100000",
26466 => "0001011010100000",
26467 => "0001011010100000",
26468 => "0001011010100100",
26469 => "0001011010100100",
26470 => "0001011010100100",
26471 => "0001011010100100",
26472 => "0001011010101000",
26473 => "0001011010101000",
26474 => "0001011010101000",
26475 => "0001011010101100",
26476 => "0001011010101100",
26477 => "0001011010101100",
26478 => "0001011010101100",
26479 => "0001011010110000",
26480 => "0001011010110000",
26481 => "0001011010110000",
26482 => "0001011010110100",
26483 => "0001011010110100",
26484 => "0001011010110100",
26485 => "0001011010111000",
26486 => "0001011010111000",
26487 => "0001011010111000",
26488 => "0001011010111000",
26489 => "0001011010111100",
26490 => "0001011010111100",
26491 => "0001011010111100",
26492 => "0001011011000000",
26493 => "0001011011000000",
26494 => "0001011011000000",
26495 => "0001011011000000",
26496 => "0001011011000100",
26497 => "0001011011000100",
26498 => "0001011011000100",
26499 => "0001011011001000",
26500 => "0001011011001000",
26501 => "0001011011001000",
26502 => "0001011011001100",
26503 => "0001011011001100",
26504 => "0001011011001100",
26505 => "0001011011001100",
26506 => "0001011011010000",
26507 => "0001011011010000",
26508 => "0001011011010000",
26509 => "0001011011010100",
26510 => "0001011011010100",
26511 => "0001011011010100",
26512 => "0001011011010100",
26513 => "0001011011011000",
26514 => "0001011011011000",
26515 => "0001011011011000",
26516 => "0001011011011100",
26517 => "0001011011011100",
26518 => "0001011011011100",
26519 => "0001011011011100",
26520 => "0001011011100000",
26521 => "0001011011100000",
26522 => "0001011011100000",
26523 => "0001011011100100",
26524 => "0001011011100100",
26525 => "0001011011100100",
26526 => "0001011011101000",
26527 => "0001011011101000",
26528 => "0001011011101000",
26529 => "0001011011101000",
26530 => "0001011011101100",
26531 => "0001011011101100",
26532 => "0001011011101100",
26533 => "0001011011110000",
26534 => "0001011011110000",
26535 => "0001011011110000",
26536 => "0001011011110000",
26537 => "0001011011110100",
26538 => "0001011011110100",
26539 => "0001011011110100",
26540 => "0001011011111000",
26541 => "0001011011111000",
26542 => "0001011011111000",
26543 => "0001011011111100",
26544 => "0001011011111100",
26545 => "0001011011111100",
26546 => "0001011011111100",
26547 => "0001011100000000",
26548 => "0001011100000000",
26549 => "0001011100000000",
26550 => "0001011100000100",
26551 => "0001011100000100",
26552 => "0001011100000100",
26553 => "0001011100000100",
26554 => "0001011100001000",
26555 => "0001011100001000",
26556 => "0001011100001000",
26557 => "0001011100001100",
26558 => "0001011100001100",
26559 => "0001011100001100",
26560 => "0001011100010000",
26561 => "0001011100010000",
26562 => "0001011100010000",
26563 => "0001011100010000",
26564 => "0001011100010100",
26565 => "0001011100010100",
26566 => "0001011100010100",
26567 => "0001011100011000",
26568 => "0001011100011000",
26569 => "0001011100011000",
26570 => "0001011100011100",
26571 => "0001011100011100",
26572 => "0001011100011100",
26573 => "0001011100011100",
26574 => "0001011100100000",
26575 => "0001011100100000",
26576 => "0001011100100000",
26577 => "0001011100100100",
26578 => "0001011100100100",
26579 => "0001011100100100",
26580 => "0001011100100100",
26581 => "0001011100101000",
26582 => "0001011100101000",
26583 => "0001011100101000",
26584 => "0001011100101100",
26585 => "0001011100101100",
26586 => "0001011100101100",
26587 => "0001011100110000",
26588 => "0001011100110000",
26589 => "0001011100110000",
26590 => "0001011100110000",
26591 => "0001011100110100",
26592 => "0001011100110100",
26593 => "0001011100110100",
26594 => "0001011100111000",
26595 => "0001011100111000",
26596 => "0001011100111000",
26597 => "0001011100111100",
26598 => "0001011100111100",
26599 => "0001011100111100",
26600 => "0001011100111100",
26601 => "0001011101000000",
26602 => "0001011101000000",
26603 => "0001011101000000",
26604 => "0001011101000100",
26605 => "0001011101000100",
26606 => "0001011101000100",
26607 => "0001011101000100",
26608 => "0001011101001000",
26609 => "0001011101001000",
26610 => "0001011101001000",
26611 => "0001011101001100",
26612 => "0001011101001100",
26613 => "0001011101001100",
26614 => "0001011101010000",
26615 => "0001011101010000",
26616 => "0001011101010000",
26617 => "0001011101010000",
26618 => "0001011101010100",
26619 => "0001011101010100",
26620 => "0001011101010100",
26621 => "0001011101011000",
26622 => "0001011101011000",
26623 => "0001011101011000",
26624 => "0001011101011100",
26625 => "0001011101011100",
26626 => "0001011101011100",
26627 => "0001011101011100",
26628 => "0001011101100000",
26629 => "0001011101100000",
26630 => "0001011101100000",
26631 => "0001011101100100",
26632 => "0001011101100100",
26633 => "0001011101100100",
26634 => "0001011101101000",
26635 => "0001011101101000",
26636 => "0001011101101000",
26637 => "0001011101101000",
26638 => "0001011101101100",
26639 => "0001011101101100",
26640 => "0001011101101100",
26641 => "0001011101110000",
26642 => "0001011101110000",
26643 => "0001011101110000",
26644 => "0001011101110100",
26645 => "0001011101110100",
26646 => "0001011101110100",
26647 => "0001011101110100",
26648 => "0001011101111000",
26649 => "0001011101111000",
26650 => "0001011101111000",
26651 => "0001011101111100",
26652 => "0001011101111100",
26653 => "0001011101111100",
26654 => "0001011110000000",
26655 => "0001011110000000",
26656 => "0001011110000000",
26657 => "0001011110000000",
26658 => "0001011110000100",
26659 => "0001011110000100",
26660 => "0001011110000100",
26661 => "0001011110001000",
26662 => "0001011110001000",
26663 => "0001011110001000",
26664 => "0001011110001100",
26665 => "0001011110001100",
26666 => "0001011110001100",
26667 => "0001011110001100",
26668 => "0001011110010000",
26669 => "0001011110010000",
26670 => "0001011110010000",
26671 => "0001011110010100",
26672 => "0001011110010100",
26673 => "0001011110010100",
26674 => "0001011110011000",
26675 => "0001011110011000",
26676 => "0001011110011000",
26677 => "0001011110011000",
26678 => "0001011110011100",
26679 => "0001011110011100",
26680 => "0001011110011100",
26681 => "0001011110100000",
26682 => "0001011110100000",
26683 => "0001011110100000",
26684 => "0001011110100100",
26685 => "0001011110100100",
26686 => "0001011110100100",
26687 => "0001011110100100",
26688 => "0001011110101000",
26689 => "0001011110101000",
26690 => "0001011110101000",
26691 => "0001011110101100",
26692 => "0001011110101100",
26693 => "0001011110101100",
26694 => "0001011110110000",
26695 => "0001011110110000",
26696 => "0001011110110000",
26697 => "0001011110110000",
26698 => "0001011110110100",
26699 => "0001011110110100",
26700 => "0001011110110100",
26701 => "0001011110111000",
26702 => "0001011110111000",
26703 => "0001011110111000",
26704 => "0001011110111100",
26705 => "0001011110111100",
26706 => "0001011110111100",
26707 => "0001011110111100",
26708 => "0001011111000000",
26709 => "0001011111000000",
26710 => "0001011111000000",
26711 => "0001011111000100",
26712 => "0001011111000100",
26713 => "0001011111000100",
26714 => "0001011111001000",
26715 => "0001011111001000",
26716 => "0001011111001000",
26717 => "0001011111001000",
26718 => "0001011111001100",
26719 => "0001011111001100",
26720 => "0001011111001100",
26721 => "0001011111010000",
26722 => "0001011111010000",
26723 => "0001011111010000",
26724 => "0001011111010100",
26725 => "0001011111010100",
26726 => "0001011111010100",
26727 => "0001011111011000",
26728 => "0001011111011000",
26729 => "0001011111011000",
26730 => "0001011111011000",
26731 => "0001011111011100",
26732 => "0001011111011100",
26733 => "0001011111011100",
26734 => "0001011111100000",
26735 => "0001011111100000",
26736 => "0001011111100000",
26737 => "0001011111100100",
26738 => "0001011111100100",
26739 => "0001011111100100",
26740 => "0001011111100100",
26741 => "0001011111101000",
26742 => "0001011111101000",
26743 => "0001011111101000",
26744 => "0001011111101100",
26745 => "0001011111101100",
26746 => "0001011111101100",
26747 => "0001011111110000",
26748 => "0001011111110000",
26749 => "0001011111110000",
26750 => "0001011111110100",
26751 => "0001011111110100",
26752 => "0001011111110100",
26753 => "0001011111110100",
26754 => "0001011111111000",
26755 => "0001011111111000",
26756 => "0001011111111000",
26757 => "0001011111111100",
26758 => "0001011111111100",
26759 => "0001011111111100",
26760 => "0001100000000000",
26761 => "0001100000000000",
26762 => "0001100000000000",
26763 => "0001100000000000",
26764 => "0001100000000100",
26765 => "0001100000000100",
26766 => "0001100000000100",
26767 => "0001100000001000",
26768 => "0001100000001000",
26769 => "0001100000001000",
26770 => "0001100000001100",
26771 => "0001100000001100",
26772 => "0001100000001100",
26773 => "0001100000010000",
26774 => "0001100000010000",
26775 => "0001100000010000",
26776 => "0001100000010000",
26777 => "0001100000010100",
26778 => "0001100000010100",
26779 => "0001100000010100",
26780 => "0001100000011000",
26781 => "0001100000011000",
26782 => "0001100000011000",
26783 => "0001100000011100",
26784 => "0001100000011100",
26785 => "0001100000011100",
26786 => "0001100000011100",
26787 => "0001100000100000",
26788 => "0001100000100000",
26789 => "0001100000100000",
26790 => "0001100000100100",
26791 => "0001100000100100",
26792 => "0001100000100100",
26793 => "0001100000101000",
26794 => "0001100000101000",
26795 => "0001100000101000",
26796 => "0001100000101100",
26797 => "0001100000101100",
26798 => "0001100000101100",
26799 => "0001100000101100",
26800 => "0001100000110000",
26801 => "0001100000110000",
26802 => "0001100000110000",
26803 => "0001100000110100",
26804 => "0001100000110100",
26805 => "0001100000110100",
26806 => "0001100000111000",
26807 => "0001100000111000",
26808 => "0001100000111000",
26809 => "0001100000111100",
26810 => "0001100000111100",
26811 => "0001100000111100",
26812 => "0001100000111100",
26813 => "0001100001000000",
26814 => "0001100001000000",
26815 => "0001100001000000",
26816 => "0001100001000100",
26817 => "0001100001000100",
26818 => "0001100001000100",
26819 => "0001100001001000",
26820 => "0001100001001000",
26821 => "0001100001001000",
26822 => "0001100001001100",
26823 => "0001100001001100",
26824 => "0001100001001100",
26825 => "0001100001001100",
26826 => "0001100001010000",
26827 => "0001100001010000",
26828 => "0001100001010000",
26829 => "0001100001010100",
26830 => "0001100001010100",
26831 => "0001100001010100",
26832 => "0001100001011000",
26833 => "0001100001011000",
26834 => "0001100001011000",
26835 => "0001100001011100",
26836 => "0001100001011100",
26837 => "0001100001011100",
26838 => "0001100001011100",
26839 => "0001100001100000",
26840 => "0001100001100000",
26841 => "0001100001100000",
26842 => "0001100001100100",
26843 => "0001100001100100",
26844 => "0001100001100100",
26845 => "0001100001101000",
26846 => "0001100001101000",
26847 => "0001100001101000",
26848 => "0001100001101100",
26849 => "0001100001101100",
26850 => "0001100001101100",
26851 => "0001100001101100",
26852 => "0001100001110000",
26853 => "0001100001110000",
26854 => "0001100001110000",
26855 => "0001100001110100",
26856 => "0001100001110100",
26857 => "0001100001110100",
26858 => "0001100001111000",
26859 => "0001100001111000",
26860 => "0001100001111000",
26861 => "0001100001111100",
26862 => "0001100001111100",
26863 => "0001100001111100",
26864 => "0001100001111100",
26865 => "0001100010000000",
26866 => "0001100010000000",
26867 => "0001100010000000",
26868 => "0001100010000100",
26869 => "0001100010000100",
26870 => "0001100010000100",
26871 => "0001100010001000",
26872 => "0001100010001000",
26873 => "0001100010001000",
26874 => "0001100010001100",
26875 => "0001100010001100",
26876 => "0001100010001100",
26877 => "0001100010010000",
26878 => "0001100010010000",
26879 => "0001100010010000",
26880 => "0001100010010000",
26881 => "0001100010010100",
26882 => "0001100010010100",
26883 => "0001100010010100",
26884 => "0001100010011000",
26885 => "0001100010011000",
26886 => "0001100010011000",
26887 => "0001100010011100",
26888 => "0001100010011100",
26889 => "0001100010011100",
26890 => "0001100010100000",
26891 => "0001100010100000",
26892 => "0001100010100000",
26893 => "0001100010100000",
26894 => "0001100010100100",
26895 => "0001100010100100",
26896 => "0001100010100100",
26897 => "0001100010101000",
26898 => "0001100010101000",
26899 => "0001100010101000",
26900 => "0001100010101100",
26901 => "0001100010101100",
26902 => "0001100010101100",
26903 => "0001100010110000",
26904 => "0001100010110000",
26905 => "0001100010110000",
26906 => "0001100010110100",
26907 => "0001100010110100",
26908 => "0001100010110100",
26909 => "0001100010110100",
26910 => "0001100010111000",
26911 => "0001100010111000",
26912 => "0001100010111000",
26913 => "0001100010111100",
26914 => "0001100010111100",
26915 => "0001100010111100",
26916 => "0001100011000000",
26917 => "0001100011000000",
26918 => "0001100011000000",
26919 => "0001100011000100",
26920 => "0001100011000100",
26921 => "0001100011000100",
26922 => "0001100011001000",
26923 => "0001100011001000",
26924 => "0001100011001000",
26925 => "0001100011001000",
26926 => "0001100011001100",
26927 => "0001100011001100",
26928 => "0001100011001100",
26929 => "0001100011010000",
26930 => "0001100011010000",
26931 => "0001100011010000",
26932 => "0001100011010100",
26933 => "0001100011010100",
26934 => "0001100011010100",
26935 => "0001100011011000",
26936 => "0001100011011000",
26937 => "0001100011011000",
26938 => "0001100011011100",
26939 => "0001100011011100",
26940 => "0001100011011100",
26941 => "0001100011011100",
26942 => "0001100011100000",
26943 => "0001100011100000",
26944 => "0001100011100000",
26945 => "0001100011100100",
26946 => "0001100011100100",
26947 => "0001100011100100",
26948 => "0001100011101000",
26949 => "0001100011101000",
26950 => "0001100011101000",
26951 => "0001100011101100",
26952 => "0001100011101100",
26953 => "0001100011101100",
26954 => "0001100011110000",
26955 => "0001100011110000",
26956 => "0001100011110000",
26957 => "0001100011110000",
26958 => "0001100011110100",
26959 => "0001100011110100",
26960 => "0001100011110100",
26961 => "0001100011111000",
26962 => "0001100011111000",
26963 => "0001100011111000",
26964 => "0001100011111100",
26965 => "0001100011111100",
26966 => "0001100011111100",
26967 => "0001100100000000",
26968 => "0001100100000000",
26969 => "0001100100000000",
26970 => "0001100100000100",
26971 => "0001100100000100",
26972 => "0001100100000100",
26973 => "0001100100000100",
26974 => "0001100100001000",
26975 => "0001100100001000",
26976 => "0001100100001000",
26977 => "0001100100001100",
26978 => "0001100100001100",
26979 => "0001100100001100",
26980 => "0001100100010000",
26981 => "0001100100010000",
26982 => "0001100100010000",
26983 => "0001100100010100",
26984 => "0001100100010100",
26985 => "0001100100010100",
26986 => "0001100100011000",
26987 => "0001100100011000",
26988 => "0001100100011000",
26989 => "0001100100011100",
26990 => "0001100100011100",
26991 => "0001100100011100",
26992 => "0001100100011100",
26993 => "0001100100100000",
26994 => "0001100100100000",
26995 => "0001100100100000",
26996 => "0001100100100100",
26997 => "0001100100100100",
26998 => "0001100100100100",
26999 => "0001100100101000",
27000 => "0001100100101000",
27001 => "0001100100101000",
27002 => "0001100100101100",
27003 => "0001100100101100",
27004 => "0001100100101100",
27005 => "0001100100110000",
27006 => "0001100100110000",
27007 => "0001100100110000",
27008 => "0001100100110100",
27009 => "0001100100110100",
27010 => "0001100100110100",
27011 => "0001100100110100",
27012 => "0001100100111000",
27013 => "0001100100111000",
27014 => "0001100100111000",
27015 => "0001100100111100",
27016 => "0001100100111100",
27017 => "0001100100111100",
27018 => "0001100101000000",
27019 => "0001100101000000",
27020 => "0001100101000000",
27021 => "0001100101000100",
27022 => "0001100101000100",
27023 => "0001100101000100",
27024 => "0001100101001000",
27025 => "0001100101001000",
27026 => "0001100101001000",
27027 => "0001100101001100",
27028 => "0001100101001100",
27029 => "0001100101001100",
27030 => "0001100101001100",
27031 => "0001100101010000",
27032 => "0001100101010000",
27033 => "0001100101010000",
27034 => "0001100101010100",
27035 => "0001100101010100",
27036 => "0001100101010100",
27037 => "0001100101011000",
27038 => "0001100101011000",
27039 => "0001100101011000",
27040 => "0001100101011100",
27041 => "0001100101011100",
27042 => "0001100101011100",
27043 => "0001100101100000",
27044 => "0001100101100000",
27045 => "0001100101100000",
27046 => "0001100101100100",
27047 => "0001100101100100",
27048 => "0001100101100100",
27049 => "0001100101101000",
27050 => "0001100101101000",
27051 => "0001100101101000",
27052 => "0001100101101000",
27053 => "0001100101101100",
27054 => "0001100101101100",
27055 => "0001100101101100",
27056 => "0001100101110000",
27057 => "0001100101110000",
27058 => "0001100101110000",
27059 => "0001100101110100",
27060 => "0001100101110100",
27061 => "0001100101110100",
27062 => "0001100101111000",
27063 => "0001100101111000",
27064 => "0001100101111000",
27065 => "0001100101111100",
27066 => "0001100101111100",
27067 => "0001100101111100",
27068 => "0001100110000000",
27069 => "0001100110000000",
27070 => "0001100110000000",
27071 => "0001100110000100",
27072 => "0001100110000100",
27073 => "0001100110000100",
27074 => "0001100110001000",
27075 => "0001100110001000",
27076 => "0001100110001000",
27077 => "0001100110001000",
27078 => "0001100110001100",
27079 => "0001100110001100",
27080 => "0001100110001100",
27081 => "0001100110010000",
27082 => "0001100110010000",
27083 => "0001100110010000",
27084 => "0001100110010100",
27085 => "0001100110010100",
27086 => "0001100110010100",
27087 => "0001100110011000",
27088 => "0001100110011000",
27089 => "0001100110011000",
27090 => "0001100110011100",
27091 => "0001100110011100",
27092 => "0001100110011100",
27093 => "0001100110100000",
27094 => "0001100110100000",
27095 => "0001100110100000",
27096 => "0001100110100100",
27097 => "0001100110100100",
27098 => "0001100110100100",
27099 => "0001100110100100",
27100 => "0001100110101000",
27101 => "0001100110101000",
27102 => "0001100110101000",
27103 => "0001100110101100",
27104 => "0001100110101100",
27105 => "0001100110101100",
27106 => "0001100110110000",
27107 => "0001100110110000",
27108 => "0001100110110000",
27109 => "0001100110110100",
27110 => "0001100110110100",
27111 => "0001100110110100",
27112 => "0001100110111000",
27113 => "0001100110111000",
27114 => "0001100110111000",
27115 => "0001100110111100",
27116 => "0001100110111100",
27117 => "0001100110111100",
27118 => "0001100111000000",
27119 => "0001100111000000",
27120 => "0001100111000000",
27121 => "0001100111000100",
27122 => "0001100111000100",
27123 => "0001100111000100",
27124 => "0001100111001000",
27125 => "0001100111001000",
27126 => "0001100111001000",
27127 => "0001100111001000",
27128 => "0001100111001100",
27129 => "0001100111001100",
27130 => "0001100111001100",
27131 => "0001100111010000",
27132 => "0001100111010000",
27133 => "0001100111010000",
27134 => "0001100111010100",
27135 => "0001100111010100",
27136 => "0001100111010100",
27137 => "0001100111011000",
27138 => "0001100111011000",
27139 => "0001100111011000",
27140 => "0001100111011100",
27141 => "0001100111011100",
27142 => "0001100111011100",
27143 => "0001100111100000",
27144 => "0001100111100000",
27145 => "0001100111100000",
27146 => "0001100111100100",
27147 => "0001100111100100",
27148 => "0001100111100100",
27149 => "0001100111101000",
27150 => "0001100111101000",
27151 => "0001100111101000",
27152 => "0001100111101100",
27153 => "0001100111101100",
27154 => "0001100111101100",
27155 => "0001100111110000",
27156 => "0001100111110000",
27157 => "0001100111110000",
27158 => "0001100111110000",
27159 => "0001100111110100",
27160 => "0001100111110100",
27161 => "0001100111110100",
27162 => "0001100111111000",
27163 => "0001100111111000",
27164 => "0001100111111000",
27165 => "0001100111111100",
27166 => "0001100111111100",
27167 => "0001100111111100",
27168 => "0001101000000000",
27169 => "0001101000000000",
27170 => "0001101000000000",
27171 => "0001101000000100",
27172 => "0001101000000100",
27173 => "0001101000000100",
27174 => "0001101000001000",
27175 => "0001101000001000",
27176 => "0001101000001000",
27177 => "0001101000001100",
27178 => "0001101000001100",
27179 => "0001101000001100",
27180 => "0001101000010000",
27181 => "0001101000010000",
27182 => "0001101000010000",
27183 => "0001101000010100",
27184 => "0001101000010100",
27185 => "0001101000010100",
27186 => "0001101000011000",
27187 => "0001101000011000",
27188 => "0001101000011000",
27189 => "0001101000011100",
27190 => "0001101000011100",
27191 => "0001101000011100",
27192 => "0001101000100000",
27193 => "0001101000100000",
27194 => "0001101000100000",
27195 => "0001101000100000",
27196 => "0001101000100100",
27197 => "0001101000100100",
27198 => "0001101000100100",
27199 => "0001101000101000",
27200 => "0001101000101000",
27201 => "0001101000101000",
27202 => "0001101000101100",
27203 => "0001101000101100",
27204 => "0001101000101100",
27205 => "0001101000110000",
27206 => "0001101000110000",
27207 => "0001101000110000",
27208 => "0001101000110100",
27209 => "0001101000110100",
27210 => "0001101000110100",
27211 => "0001101000111000",
27212 => "0001101000111000",
27213 => "0001101000111000",
27214 => "0001101000111100",
27215 => "0001101000111100",
27216 => "0001101000111100",
27217 => "0001101001000000",
27218 => "0001101001000000",
27219 => "0001101001000000",
27220 => "0001101001000100",
27221 => "0001101001000100",
27222 => "0001101001000100",
27223 => "0001101001001000",
27224 => "0001101001001000",
27225 => "0001101001001000",
27226 => "0001101001001100",
27227 => "0001101001001100",
27228 => "0001101001001100",
27229 => "0001101001010000",
27230 => "0001101001010000",
27231 => "0001101001010000",
27232 => "0001101001010100",
27233 => "0001101001010100",
27234 => "0001101001010100",
27235 => "0001101001011000",
27236 => "0001101001011000",
27237 => "0001101001011000",
27238 => "0001101001011000",
27239 => "0001101001011100",
27240 => "0001101001011100",
27241 => "0001101001011100",
27242 => "0001101001100000",
27243 => "0001101001100000",
27244 => "0001101001100000",
27245 => "0001101001100100",
27246 => "0001101001100100",
27247 => "0001101001100100",
27248 => "0001101001101000",
27249 => "0001101001101000",
27250 => "0001101001101000",
27251 => "0001101001101100",
27252 => "0001101001101100",
27253 => "0001101001101100",
27254 => "0001101001110000",
27255 => "0001101001110000",
27256 => "0001101001110000",
27257 => "0001101001110100",
27258 => "0001101001110100",
27259 => "0001101001110100",
27260 => "0001101001111000",
27261 => "0001101001111000",
27262 => "0001101001111000",
27263 => "0001101001111100",
27264 => "0001101001111100",
27265 => "0001101001111100",
27266 => "0001101010000000",
27267 => "0001101010000000",
27268 => "0001101010000000",
27269 => "0001101010000100",
27270 => "0001101010000100",
27271 => "0001101010000100",
27272 => "0001101010001000",
27273 => "0001101010001000",
27274 => "0001101010001000",
27275 => "0001101010001100",
27276 => "0001101010001100",
27277 => "0001101010001100",
27278 => "0001101010010000",
27279 => "0001101010010000",
27280 => "0001101010010000",
27281 => "0001101010010100",
27282 => "0001101010010100",
27283 => "0001101010010100",
27284 => "0001101010011000",
27285 => "0001101010011000",
27286 => "0001101010011000",
27287 => "0001101010011100",
27288 => "0001101010011100",
27289 => "0001101010011100",
27290 => "0001101010100000",
27291 => "0001101010100000",
27292 => "0001101010100000",
27293 => "0001101010100100",
27294 => "0001101010100100",
27295 => "0001101010100100",
27296 => "0001101010101000",
27297 => "0001101010101000",
27298 => "0001101010101000",
27299 => "0001101010101100",
27300 => "0001101010101100",
27301 => "0001101010101100",
27302 => "0001101010110000",
27303 => "0001101010110000",
27304 => "0001101010110000",
27305 => "0001101010110100",
27306 => "0001101010110100",
27307 => "0001101010110100",
27308 => "0001101010110100",
27309 => "0001101010111000",
27310 => "0001101010111000",
27311 => "0001101010111000",
27312 => "0001101010111100",
27313 => "0001101010111100",
27314 => "0001101010111100",
27315 => "0001101011000000",
27316 => "0001101011000000",
27317 => "0001101011000000",
27318 => "0001101011000100",
27319 => "0001101011000100",
27320 => "0001101011000100",
27321 => "0001101011001000",
27322 => "0001101011001000",
27323 => "0001101011001000",
27324 => "0001101011001100",
27325 => "0001101011001100",
27326 => "0001101011001100",
27327 => "0001101011010000",
27328 => "0001101011010000",
27329 => "0001101011010000",
27330 => "0001101011010100",
27331 => "0001101011010100",
27332 => "0001101011010100",
27333 => "0001101011011000",
27334 => "0001101011011000",
27335 => "0001101011011000",
27336 => "0001101011011100",
27337 => "0001101011011100",
27338 => "0001101011011100",
27339 => "0001101011100000",
27340 => "0001101011100000",
27341 => "0001101011100000",
27342 => "0001101011100100",
27343 => "0001101011100100",
27344 => "0001101011100100",
27345 => "0001101011101000",
27346 => "0001101011101000",
27347 => "0001101011101000",
27348 => "0001101011101100",
27349 => "0001101011101100",
27350 => "0001101011101100",
27351 => "0001101011110000",
27352 => "0001101011110000",
27353 => "0001101011110000",
27354 => "0001101011110100",
27355 => "0001101011110100",
27356 => "0001101011110100",
27357 => "0001101011111000",
27358 => "0001101011111000",
27359 => "0001101011111000",
27360 => "0001101011111100",
27361 => "0001101011111100",
27362 => "0001101011111100",
27363 => "0001101100000000",
27364 => "0001101100000000",
27365 => "0001101100000000",
27366 => "0001101100000100",
27367 => "0001101100000100",
27368 => "0001101100000100",
27369 => "0001101100001000",
27370 => "0001101100001000",
27371 => "0001101100001000",
27372 => "0001101100001100",
27373 => "0001101100001100",
27374 => "0001101100001100",
27375 => "0001101100010000",
27376 => "0001101100010000",
27377 => "0001101100010000",
27378 => "0001101100010100",
27379 => "0001101100010100",
27380 => "0001101100010100",
27381 => "0001101100011000",
27382 => "0001101100011000",
27383 => "0001101100011000",
27384 => "0001101100011100",
27385 => "0001101100011100",
27386 => "0001101100011100",
27387 => "0001101100100000",
27388 => "0001101100100000",
27389 => "0001101100100000",
27390 => "0001101100100100",
27391 => "0001101100100100",
27392 => "0001101100100100",
27393 => "0001101100101000",
27394 => "0001101100101000",
27395 => "0001101100101000",
27396 => "0001101100101100",
27397 => "0001101100101100",
27398 => "0001101100101100",
27399 => "0001101100110000",
27400 => "0001101100110000",
27401 => "0001101100110000",
27402 => "0001101100110100",
27403 => "0001101100110100",
27404 => "0001101100110100",
27405 => "0001101100111000",
27406 => "0001101100111000",
27407 => "0001101100111000",
27408 => "0001101100111100",
27409 => "0001101100111100",
27410 => "0001101100111100",
27411 => "0001101101000000",
27412 => "0001101101000000",
27413 => "0001101101000000",
27414 => "0001101101000100",
27415 => "0001101101000100",
27416 => "0001101101000100",
27417 => "0001101101001000",
27418 => "0001101101001000",
27419 => "0001101101001000",
27420 => "0001101101001100",
27421 => "0001101101001100",
27422 => "0001101101001100",
27423 => "0001101101010000",
27424 => "0001101101010000",
27425 => "0001101101010000",
27426 => "0001101101010100",
27427 => "0001101101010100",
27428 => "0001101101010100",
27429 => "0001101101011000",
27430 => "0001101101011000",
27431 => "0001101101011000",
27432 => "0001101101011100",
27433 => "0001101101011100",
27434 => "0001101101011100",
27435 => "0001101101100000",
27436 => "0001101101100000",
27437 => "0001101101100000",
27438 => "0001101101100100",
27439 => "0001101101100100",
27440 => "0001101101101000",
27441 => "0001101101101000",
27442 => "0001101101101000",
27443 => "0001101101101100",
27444 => "0001101101101100",
27445 => "0001101101101100",
27446 => "0001101101110000",
27447 => "0001101101110000",
27448 => "0001101101110000",
27449 => "0001101101110100",
27450 => "0001101101110100",
27451 => "0001101101110100",
27452 => "0001101101111000",
27453 => "0001101101111000",
27454 => "0001101101111000",
27455 => "0001101101111100",
27456 => "0001101101111100",
27457 => "0001101101111100",
27458 => "0001101110000000",
27459 => "0001101110000000",
27460 => "0001101110000000",
27461 => "0001101110000100",
27462 => "0001101110000100",
27463 => "0001101110000100",
27464 => "0001101110001000",
27465 => "0001101110001000",
27466 => "0001101110001000",
27467 => "0001101110001100",
27468 => "0001101110001100",
27469 => "0001101110001100",
27470 => "0001101110010000",
27471 => "0001101110010000",
27472 => "0001101110010000",
27473 => "0001101110010100",
27474 => "0001101110010100",
27475 => "0001101110010100",
27476 => "0001101110011000",
27477 => "0001101110011000",
27478 => "0001101110011000",
27479 => "0001101110011100",
27480 => "0001101110011100",
27481 => "0001101110011100",
27482 => "0001101110100000",
27483 => "0001101110100000",
27484 => "0001101110100000",
27485 => "0001101110100100",
27486 => "0001101110100100",
27487 => "0001101110100100",
27488 => "0001101110101000",
27489 => "0001101110101000",
27490 => "0001101110101000",
27491 => "0001101110101100",
27492 => "0001101110101100",
27493 => "0001101110101100",
27494 => "0001101110110000",
27495 => "0001101110110000",
27496 => "0001101110110000",
27497 => "0001101110110100",
27498 => "0001101110110100",
27499 => "0001101110110100",
27500 => "0001101110111000",
27501 => "0001101110111000",
27502 => "0001101110111000",
27503 => "0001101110111100",
27504 => "0001101110111100",
27505 => "0001101110111100",
27506 => "0001101111000000",
27507 => "0001101111000000",
27508 => "0001101111000000",
27509 => "0001101111000100",
27510 => "0001101111000100",
27511 => "0001101111001000",
27512 => "0001101111001000",
27513 => "0001101111001000",
27514 => "0001101111001100",
27515 => "0001101111001100",
27516 => "0001101111001100",
27517 => "0001101111010000",
27518 => "0001101111010000",
27519 => "0001101111010000",
27520 => "0001101111010100",
27521 => "0001101111010100",
27522 => "0001101111010100",
27523 => "0001101111011000",
27524 => "0001101111011000",
27525 => "0001101111011000",
27526 => "0001101111011100",
27527 => "0001101111011100",
27528 => "0001101111011100",
27529 => "0001101111100000",
27530 => "0001101111100000",
27531 => "0001101111100000",
27532 => "0001101111100100",
27533 => "0001101111100100",
27534 => "0001101111100100",
27535 => "0001101111101000",
27536 => "0001101111101000",
27537 => "0001101111101000",
27538 => "0001101111101100",
27539 => "0001101111101100",
27540 => "0001101111101100",
27541 => "0001101111110000",
27542 => "0001101111110000",
27543 => "0001101111110000",
27544 => "0001101111110100",
27545 => "0001101111110100",
27546 => "0001101111110100",
27547 => "0001101111111000",
27548 => "0001101111111000",
27549 => "0001101111111000",
27550 => "0001101111111100",
27551 => "0001101111111100",
27552 => "0001101111111100",
27553 => "0001110000000000",
27554 => "0001110000000000",
27555 => "0001110000000100",
27556 => "0001110000000100",
27557 => "0001110000000100",
27558 => "0001110000001000",
27559 => "0001110000001000",
27560 => "0001110000001000",
27561 => "0001110000001100",
27562 => "0001110000001100",
27563 => "0001110000001100",
27564 => "0001110000010000",
27565 => "0001110000010000",
27566 => "0001110000010000",
27567 => "0001110000010100",
27568 => "0001110000010100",
27569 => "0001110000010100",
27570 => "0001110000011000",
27571 => "0001110000011000",
27572 => "0001110000011000",
27573 => "0001110000011100",
27574 => "0001110000011100",
27575 => "0001110000011100",
27576 => "0001110000100000",
27577 => "0001110000100000",
27578 => "0001110000100000",
27579 => "0001110000100100",
27580 => "0001110000100100",
27581 => "0001110000100100",
27582 => "0001110000101000",
27583 => "0001110000101000",
27584 => "0001110000101000",
27585 => "0001110000101100",
27586 => "0001110000101100",
27587 => "0001110000101100",
27588 => "0001110000110000",
27589 => "0001110000110000",
27590 => "0001110000110100",
27591 => "0001110000110100",
27592 => "0001110000110100",
27593 => "0001110000111000",
27594 => "0001110000111000",
27595 => "0001110000111000",
27596 => "0001110000111100",
27597 => "0001110000111100",
27598 => "0001110000111100",
27599 => "0001110001000000",
27600 => "0001110001000000",
27601 => "0001110001000000",
27602 => "0001110001000100",
27603 => "0001110001000100",
27604 => "0001110001000100",
27605 => "0001110001001000",
27606 => "0001110001001000",
27607 => "0001110001001000",
27608 => "0001110001001100",
27609 => "0001110001001100",
27610 => "0001110001001100",
27611 => "0001110001010000",
27612 => "0001110001010000",
27613 => "0001110001010000",
27614 => "0001110001010100",
27615 => "0001110001010100",
27616 => "0001110001010100",
27617 => "0001110001011000",
27618 => "0001110001011000",
27619 => "0001110001011000",
27620 => "0001110001011100",
27621 => "0001110001011100",
27622 => "0001110001100000",
27623 => "0001110001100000",
27624 => "0001110001100000",
27625 => "0001110001100100",
27626 => "0001110001100100",
27627 => "0001110001100100",
27628 => "0001110001101000",
27629 => "0001110001101000",
27630 => "0001110001101000",
27631 => "0001110001101100",
27632 => "0001110001101100",
27633 => "0001110001101100",
27634 => "0001110001110000",
27635 => "0001110001110000",
27636 => "0001110001110000",
27637 => "0001110001110100",
27638 => "0001110001110100",
27639 => "0001110001110100",
27640 => "0001110001111000",
27641 => "0001110001111000",
27642 => "0001110001111000",
27643 => "0001110001111100",
27644 => "0001110001111100",
27645 => "0001110001111100",
27646 => "0001110010000000",
27647 => "0001110010000000",
27648 => "0001110010000100",
27649 => "0001110010000100",
27650 => "0001110010000100",
27651 => "0001110010001000",
27652 => "0001110010001000",
27653 => "0001110010001000",
27654 => "0001110010001100",
27655 => "0001110010001100",
27656 => "0001110010001100",
27657 => "0001110010010000",
27658 => "0001110010010000",
27659 => "0001110010010000",
27660 => "0001110010010100",
27661 => "0001110010010100",
27662 => "0001110010010100",
27663 => "0001110010011000",
27664 => "0001110010011000",
27665 => "0001110010011000",
27666 => "0001110010011100",
27667 => "0001110010011100",
27668 => "0001110010011100",
27669 => "0001110010100000",
27670 => "0001110010100000",
27671 => "0001110010100000",
27672 => "0001110010100100",
27673 => "0001110010100100",
27674 => "0001110010101000",
27675 => "0001110010101000",
27676 => "0001110010101000",
27677 => "0001110010101100",
27678 => "0001110010101100",
27679 => "0001110010101100",
27680 => "0001110010110000",
27681 => "0001110010110000",
27682 => "0001110010110000",
27683 => "0001110010110100",
27684 => "0001110010110100",
27685 => "0001110010110100",
27686 => "0001110010111000",
27687 => "0001110010111000",
27688 => "0001110010111000",
27689 => "0001110010111100",
27690 => "0001110010111100",
27691 => "0001110010111100",
27692 => "0001110011000000",
27693 => "0001110011000000",
27694 => "0001110011000000",
27695 => "0001110011000100",
27696 => "0001110011000100",
27697 => "0001110011001000",
27698 => "0001110011001000",
27699 => "0001110011001000",
27700 => "0001110011001100",
27701 => "0001110011001100",
27702 => "0001110011001100",
27703 => "0001110011010000",
27704 => "0001110011010000",
27705 => "0001110011010000",
27706 => "0001110011010100",
27707 => "0001110011010100",
27708 => "0001110011010100",
27709 => "0001110011011000",
27710 => "0001110011011000",
27711 => "0001110011011000",
27712 => "0001110011011100",
27713 => "0001110011011100",
27714 => "0001110011011100",
27715 => "0001110011100000",
27716 => "0001110011100000",
27717 => "0001110011100100",
27718 => "0001110011100100",
27719 => "0001110011100100",
27720 => "0001110011101000",
27721 => "0001110011101000",
27722 => "0001110011101000",
27723 => "0001110011101100",
27724 => "0001110011101100",
27725 => "0001110011101100",
27726 => "0001110011110000",
27727 => "0001110011110000",
27728 => "0001110011110000",
27729 => "0001110011110100",
27730 => "0001110011110100",
27731 => "0001110011110100",
27732 => "0001110011111000",
27733 => "0001110011111000",
27734 => "0001110011111000",
27735 => "0001110011111100",
27736 => "0001110011111100",
27737 => "0001110100000000",
27738 => "0001110100000000",
27739 => "0001110100000000",
27740 => "0001110100000100",
27741 => "0001110100000100",
27742 => "0001110100000100",
27743 => "0001110100001000",
27744 => "0001110100001000",
27745 => "0001110100001000",
27746 => "0001110100001100",
27747 => "0001110100001100",
27748 => "0001110100001100",
27749 => "0001110100010000",
27750 => "0001110100010000",
27751 => "0001110100010000",
27752 => "0001110100010100",
27753 => "0001110100010100",
27754 => "0001110100010100",
27755 => "0001110100011000",
27756 => "0001110100011000",
27757 => "0001110100011100",
27758 => "0001110100011100",
27759 => "0001110100011100",
27760 => "0001110100100000",
27761 => "0001110100100000",
27762 => "0001110100100000",
27763 => "0001110100100100",
27764 => "0001110100100100",
27765 => "0001110100100100",
27766 => "0001110100101000",
27767 => "0001110100101000",
27768 => "0001110100101000",
27769 => "0001110100101100",
27770 => "0001110100101100",
27771 => "0001110100101100",
27772 => "0001110100110000",
27773 => "0001110100110000",
27774 => "0001110100110100",
27775 => "0001110100110100",
27776 => "0001110100110100",
27777 => "0001110100111000",
27778 => "0001110100111000",
27779 => "0001110100111000",
27780 => "0001110100111100",
27781 => "0001110100111100",
27782 => "0001110100111100",
27783 => "0001110101000000",
27784 => "0001110101000000",
27785 => "0001110101000000",
27786 => "0001110101000100",
27787 => "0001110101000100",
27788 => "0001110101000100",
27789 => "0001110101001000",
27790 => "0001110101001000",
27791 => "0001110101001000",
27792 => "0001110101001100",
27793 => "0001110101001100",
27794 => "0001110101010000",
27795 => "0001110101010000",
27796 => "0001110101010000",
27797 => "0001110101010100",
27798 => "0001110101010100",
27799 => "0001110101010100",
27800 => "0001110101011000",
27801 => "0001110101011000",
27802 => "0001110101011000",
27803 => "0001110101011100",
27804 => "0001110101011100",
27805 => "0001110101011100",
27806 => "0001110101100000",
27807 => "0001110101100000",
27808 => "0001110101100100",
27809 => "0001110101100100",
27810 => "0001110101100100",
27811 => "0001110101101000",
27812 => "0001110101101000",
27813 => "0001110101101000",
27814 => "0001110101101100",
27815 => "0001110101101100",
27816 => "0001110101101100",
27817 => "0001110101110000",
27818 => "0001110101110000",
27819 => "0001110101110000",
27820 => "0001110101110100",
27821 => "0001110101110100",
27822 => "0001110101110100",
27823 => "0001110101111000",
27824 => "0001110101111000",
27825 => "0001110101111100",
27826 => "0001110101111100",
27827 => "0001110101111100",
27828 => "0001110110000000",
27829 => "0001110110000000",
27830 => "0001110110000000",
27831 => "0001110110000100",
27832 => "0001110110000100",
27833 => "0001110110000100",
27834 => "0001110110001000",
27835 => "0001110110001000",
27836 => "0001110110001000",
27837 => "0001110110001100",
27838 => "0001110110001100",
27839 => "0001110110001100",
27840 => "0001110110010000",
27841 => "0001110110010000",
27842 => "0001110110010100",
27843 => "0001110110010100",
27844 => "0001110110010100",
27845 => "0001110110011000",
27846 => "0001110110011000",
27847 => "0001110110011000",
27848 => "0001110110011100",
27849 => "0001110110011100",
27850 => "0001110110011100",
27851 => "0001110110100000",
27852 => "0001110110100000",
27853 => "0001110110100000",
27854 => "0001110110100100",
27855 => "0001110110100100",
27856 => "0001110110101000",
27857 => "0001110110101000",
27858 => "0001110110101000",
27859 => "0001110110101100",
27860 => "0001110110101100",
27861 => "0001110110101100",
27862 => "0001110110110000",
27863 => "0001110110110000",
27864 => "0001110110110000",
27865 => "0001110110110100",
27866 => "0001110110110100",
27867 => "0001110110110100",
27868 => "0001110110111000",
27869 => "0001110110111000",
27870 => "0001110110111100",
27871 => "0001110110111100",
27872 => "0001110110111100",
27873 => "0001110111000000",
27874 => "0001110111000000",
27875 => "0001110111000000",
27876 => "0001110111000100",
27877 => "0001110111000100",
27878 => "0001110111000100",
27879 => "0001110111001000",
27880 => "0001110111001000",
27881 => "0001110111001000",
27882 => "0001110111001100",
27883 => "0001110111001100",
27884 => "0001110111010000",
27885 => "0001110111010000",
27886 => "0001110111010000",
27887 => "0001110111010100",
27888 => "0001110111010100",
27889 => "0001110111010100",
27890 => "0001110111011000",
27891 => "0001110111011000",
27892 => "0001110111011000",
27893 => "0001110111011100",
27894 => "0001110111011100",
27895 => "0001110111011100",
27896 => "0001110111100000",
27897 => "0001110111100000",
27898 => "0001110111100100",
27899 => "0001110111100100",
27900 => "0001110111100100",
27901 => "0001110111101000",
27902 => "0001110111101000",
27903 => "0001110111101000",
27904 => "0001110111101100",
27905 => "0001110111101100",
27906 => "0001110111101100",
27907 => "0001110111110000",
27908 => "0001110111110000",
27909 => "0001110111110000",
27910 => "0001110111110100",
27911 => "0001110111110100",
27912 => "0001110111111000",
27913 => "0001110111111000",
27914 => "0001110111111000",
27915 => "0001110111111100",
27916 => "0001110111111100",
27917 => "0001110111111100",
27918 => "0001111000000000",
27919 => "0001111000000000",
27920 => "0001111000000000",
27921 => "0001111000000100",
27922 => "0001111000000100",
27923 => "0001111000000100",
27924 => "0001111000001000",
27925 => "0001111000001000",
27926 => "0001111000001100",
27927 => "0001111000001100",
27928 => "0001111000001100",
27929 => "0001111000010000",
27930 => "0001111000010000",
27931 => "0001111000010000",
27932 => "0001111000010100",
27933 => "0001111000010100",
27934 => "0001111000010100",
27935 => "0001111000011000",
27936 => "0001111000011000",
27937 => "0001111000011100",
27938 => "0001111000011100",
27939 => "0001111000011100",
27940 => "0001111000100000",
27941 => "0001111000100000",
27942 => "0001111000100000",
27943 => "0001111000100100",
27944 => "0001111000100100",
27945 => "0001111000100100",
27946 => "0001111000101000",
27947 => "0001111000101000",
27948 => "0001111000101000",
27949 => "0001111000101100",
27950 => "0001111000101100",
27951 => "0001111000110000",
27952 => "0001111000110000",
27953 => "0001111000110000",
27954 => "0001111000110100",
27955 => "0001111000110100",
27956 => "0001111000110100",
27957 => "0001111000111000",
27958 => "0001111000111000",
27959 => "0001111000111000",
27960 => "0001111000111100",
27961 => "0001111000111100",
27962 => "0001111001000000",
27963 => "0001111001000000",
27964 => "0001111001000000",
27965 => "0001111001000100",
27966 => "0001111001000100",
27967 => "0001111001000100",
27968 => "0001111001001000",
27969 => "0001111001001000",
27970 => "0001111001001000",
27971 => "0001111001001100",
27972 => "0001111001001100",
27973 => "0001111001010000",
27974 => "0001111001010000",
27975 => "0001111001010000",
27976 => "0001111001010100",
27977 => "0001111001010100",
27978 => "0001111001010100",
27979 => "0001111001011000",
27980 => "0001111001011000",
27981 => "0001111001011000",
27982 => "0001111001011100",
27983 => "0001111001011100",
27984 => "0001111001011100",
27985 => "0001111001100000",
27986 => "0001111001100000",
27987 => "0001111001100100",
27988 => "0001111001100100",
27989 => "0001111001100100",
27990 => "0001111001101000",
27991 => "0001111001101000",
27992 => "0001111001101000",
27993 => "0001111001101100",
27994 => "0001111001101100",
27995 => "0001111001101100",
27996 => "0001111001110000",
27997 => "0001111001110000",
27998 => "0001111001110100",
27999 => "0001111001110100",
28000 => "0001111001110100",
28001 => "0001111001111000",
28002 => "0001111001111000",
28003 => "0001111001111000",
28004 => "0001111001111100",
28005 => "0001111001111100",
28006 => "0001111001111100",
28007 => "0001111010000000",
28008 => "0001111010000000",
28009 => "0001111010000100",
28010 => "0001111010000100",
28011 => "0001111010000100",
28012 => "0001111010001000",
28013 => "0001111010001000",
28014 => "0001111010001000",
28015 => "0001111010001100",
28016 => "0001111010001100",
28017 => "0001111010001100",
28018 => "0001111010010000",
28019 => "0001111010010000",
28020 => "0001111010010100",
28021 => "0001111010010100",
28022 => "0001111010010100",
28023 => "0001111010011000",
28024 => "0001111010011000",
28025 => "0001111010011000",
28026 => "0001111010011100",
28027 => "0001111010011100",
28028 => "0001111010011100",
28029 => "0001111010100000",
28030 => "0001111010100000",
28031 => "0001111010100100",
28032 => "0001111010100100",
28033 => "0001111010100100",
28034 => "0001111010101000",
28035 => "0001111010101000",
28036 => "0001111010101000",
28037 => "0001111010101100",
28038 => "0001111010101100",
28039 => "0001111010101100",
28040 => "0001111010110000",
28041 => "0001111010110000",
28042 => "0001111010110100",
28043 => "0001111010110100",
28044 => "0001111010110100",
28045 => "0001111010111000",
28046 => "0001111010111000",
28047 => "0001111010111000",
28048 => "0001111010111100",
28049 => "0001111010111100",
28050 => "0001111010111100",
28051 => "0001111011000000",
28052 => "0001111011000000",
28053 => "0001111011000100",
28054 => "0001111011000100",
28055 => "0001111011000100",
28056 => "0001111011001000",
28057 => "0001111011001000",
28058 => "0001111011001000",
28059 => "0001111011001100",
28060 => "0001111011001100",
28061 => "0001111011001100",
28062 => "0001111011010000",
28063 => "0001111011010000",
28064 => "0001111011010100",
28065 => "0001111011010100",
28066 => "0001111011010100",
28067 => "0001111011011000",
28068 => "0001111011011000",
28069 => "0001111011011000",
28070 => "0001111011011100",
28071 => "0001111011011100",
28072 => "0001111011100000",
28073 => "0001111011100000",
28074 => "0001111011100000",
28075 => "0001111011100100",
28076 => "0001111011100100",
28077 => "0001111011100100",
28078 => "0001111011101000",
28079 => "0001111011101000",
28080 => "0001111011101000",
28081 => "0001111011101100",
28082 => "0001111011101100",
28083 => "0001111011110000",
28084 => "0001111011110000",
28085 => "0001111011110000",
28086 => "0001111011110100",
28087 => "0001111011110100",
28088 => "0001111011110100",
28089 => "0001111011111000",
28090 => "0001111011111000",
28091 => "0001111011111000",
28092 => "0001111011111100",
28093 => "0001111011111100",
28094 => "0001111100000000",
28095 => "0001111100000000",
28096 => "0001111100000000",
28097 => "0001111100000100",
28098 => "0001111100000100",
28099 => "0001111100000100",
28100 => "0001111100001000",
28101 => "0001111100001000",
28102 => "0001111100001100",
28103 => "0001111100001100",
28104 => "0001111100001100",
28105 => "0001111100010000",
28106 => "0001111100010000",
28107 => "0001111100010000",
28108 => "0001111100010100",
28109 => "0001111100010100",
28110 => "0001111100010100",
28111 => "0001111100011000",
28112 => "0001111100011000",
28113 => "0001111100011100",
28114 => "0001111100011100",
28115 => "0001111100011100",
28116 => "0001111100100000",
28117 => "0001111100100000",
28118 => "0001111100100000",
28119 => "0001111100100100",
28120 => "0001111100100100",
28121 => "0001111100100100",
28122 => "0001111100101000",
28123 => "0001111100101000",
28124 => "0001111100101100",
28125 => "0001111100101100",
28126 => "0001111100101100",
28127 => "0001111100110000",
28128 => "0001111100110000",
28129 => "0001111100110000",
28130 => "0001111100110100",
28131 => "0001111100110100",
28132 => "0001111100111000",
28133 => "0001111100111000",
28134 => "0001111100111000",
28135 => "0001111100111100",
28136 => "0001111100111100",
28137 => "0001111100111100",
28138 => "0001111101000000",
28139 => "0001111101000000",
28140 => "0001111101000100",
28141 => "0001111101000100",
28142 => "0001111101000100",
28143 => "0001111101001000",
28144 => "0001111101001000",
28145 => "0001111101001000",
28146 => "0001111101001100",
28147 => "0001111101001100",
28148 => "0001111101001100",
28149 => "0001111101010000",
28150 => "0001111101010000",
28151 => "0001111101010100",
28152 => "0001111101010100",
28153 => "0001111101010100",
28154 => "0001111101011000",
28155 => "0001111101011000",
28156 => "0001111101011000",
28157 => "0001111101011100",
28158 => "0001111101011100",
28159 => "0001111101100000",
28160 => "0001111101100000",
28161 => "0001111101100000",
28162 => "0001111101100100",
28163 => "0001111101100100",
28164 => "0001111101100100",
28165 => "0001111101101000",
28166 => "0001111101101000",
28167 => "0001111101101000",
28168 => "0001111101101100",
28169 => "0001111101101100",
28170 => "0001111101110000",
28171 => "0001111101110000",
28172 => "0001111101110000",
28173 => "0001111101110100",
28174 => "0001111101110100",
28175 => "0001111101110100",
28176 => "0001111101111000",
28177 => "0001111101111000",
28178 => "0001111101111100",
28179 => "0001111101111100",
28180 => "0001111101111100",
28181 => "0001111110000000",
28182 => "0001111110000000",
28183 => "0001111110000000",
28184 => "0001111110000100",
28185 => "0001111110000100",
28186 => "0001111110001000",
28187 => "0001111110001000",
28188 => "0001111110001000",
28189 => "0001111110001100",
28190 => "0001111110001100",
28191 => "0001111110001100",
28192 => "0001111110010000",
28193 => "0001111110010000",
28194 => "0001111110010100",
28195 => "0001111110010100",
28196 => "0001111110010100",
28197 => "0001111110011000",
28198 => "0001111110011000",
28199 => "0001111110011000",
28200 => "0001111110011100",
28201 => "0001111110011100",
28202 => "0001111110011100",
28203 => "0001111110100000",
28204 => "0001111110100000",
28205 => "0001111110100100",
28206 => "0001111110100100",
28207 => "0001111110100100",
28208 => "0001111110101000",
28209 => "0001111110101000",
28210 => "0001111110101000",
28211 => "0001111110101100",
28212 => "0001111110101100",
28213 => "0001111110110000",
28214 => "0001111110110000",
28215 => "0001111110110000",
28216 => "0001111110110100",
28217 => "0001111110110100",
28218 => "0001111110110100",
28219 => "0001111110111000",
28220 => "0001111110111000",
28221 => "0001111110111100",
28222 => "0001111110111100",
28223 => "0001111110111100",
28224 => "0001111111000000",
28225 => "0001111111000000",
28226 => "0001111111000000",
28227 => "0001111111000100",
28228 => "0001111111000100",
28229 => "0001111111001000",
28230 => "0001111111001000",
28231 => "0001111111001000",
28232 => "0001111111001100",
28233 => "0001111111001100",
28234 => "0001111111001100",
28235 => "0001111111010000",
28236 => "0001111111010000",
28237 => "0001111111010100",
28238 => "0001111111010100",
28239 => "0001111111010100",
28240 => "0001111111011000",
28241 => "0001111111011000",
28242 => "0001111111011000",
28243 => "0001111111011100",
28244 => "0001111111011100",
28245 => "0001111111100000",
28246 => "0001111111100000",
28247 => "0001111111100000",
28248 => "0001111111100100",
28249 => "0001111111100100",
28250 => "0001111111100100",
28251 => "0001111111101000",
28252 => "0001111111101000",
28253 => "0001111111101100",
28254 => "0001111111101100",
28255 => "0001111111101100",
28256 => "0001111111110000",
28257 => "0001111111110000",
28258 => "0001111111110000",
28259 => "0001111111110100",
28260 => "0001111111110100",
28261 => "0001111111111000",
28262 => "0001111111111000",
28263 => "0001111111111000",
28264 => "0001111111111100",
28265 => "0001111111111100",
28266 => "0001111111111100",
28267 => "0010000000000000",
28268 => "0010000000000000",
28269 => "0010000000000000",
28270 => "0010000000000000",
28271 => "0010000000001000",
28272 => "0010000000001000",
28273 => "0010000000001000",
28274 => "0010000000001000",
28275 => "0010000000001000",
28276 => "0010000000010000",
28277 => "0010000000010000",
28278 => "0010000000010000",
28279 => "0010000000010000",
28280 => "0010000000010000",
28281 => "0010000000011000",
28282 => "0010000000011000",
28283 => "0010000000011000",
28284 => "0010000000011000",
28285 => "0010000000011000",
28286 => "0010000000011000",
28287 => "0010000000100000",
28288 => "0010000000100000",
28289 => "0010000000100000",
28290 => "0010000000100000",
28291 => "0010000000100000",
28292 => "0010000000101000",
28293 => "0010000000101000",
28294 => "0010000000101000",
28295 => "0010000000101000",
28296 => "0010000000101000",
28297 => "0010000000110000",
28298 => "0010000000110000",
28299 => "0010000000110000",
28300 => "0010000000110000",
28301 => "0010000000110000",
28302 => "0010000000110000",
28303 => "0010000000111000",
28304 => "0010000000111000",
28305 => "0010000000111000",
28306 => "0010000000111000",
28307 => "0010000000111000",
28308 => "0010000001000000",
28309 => "0010000001000000",
28310 => "0010000001000000",
28311 => "0010000001000000",
28312 => "0010000001000000",
28313 => "0010000001001000",
28314 => "0010000001001000",
28315 => "0010000001001000",
28316 => "0010000001001000",
28317 => "0010000001001000",
28318 => "0010000001001000",
28319 => "0010000001010000",
28320 => "0010000001010000",
28321 => "0010000001010000",
28322 => "0010000001010000",
28323 => "0010000001010000",
28324 => "0010000001011000",
28325 => "0010000001011000",
28326 => "0010000001011000",
28327 => "0010000001011000",
28328 => "0010000001011000",
28329 => "0010000001100000",
28330 => "0010000001100000",
28331 => "0010000001100000",
28332 => "0010000001100000",
28333 => "0010000001100000",
28334 => "0010000001100000",
28335 => "0010000001101000",
28336 => "0010000001101000",
28337 => "0010000001101000",
28338 => "0010000001101000",
28339 => "0010000001101000",
28340 => "0010000001110000",
28341 => "0010000001110000",
28342 => "0010000001110000",
28343 => "0010000001110000",
28344 => "0010000001110000",
28345 => "0010000001111000",
28346 => "0010000001111000",
28347 => "0010000001111000",
28348 => "0010000001111000",
28349 => "0010000001111000",
28350 => "0010000010000000",
28351 => "0010000010000000",
28352 => "0010000010000000",
28353 => "0010000010000000",
28354 => "0010000010000000",
28355 => "0010000010000000",
28356 => "0010000010001000",
28357 => "0010000010001000",
28358 => "0010000010001000",
28359 => "0010000010001000",
28360 => "0010000010001000",
28361 => "0010000010010000",
28362 => "0010000010010000",
28363 => "0010000010010000",
28364 => "0010000010010000",
28365 => "0010000010010000",
28366 => "0010000010011000",
28367 => "0010000010011000",
28368 => "0010000010011000",
28369 => "0010000010011000",
28370 => "0010000010011000",
28371 => "0010000010011000",
28372 => "0010000010100000",
28373 => "0010000010100000",
28374 => "0010000010100000",
28375 => "0010000010100000",
28376 => "0010000010100000",
28377 => "0010000010101000",
28378 => "0010000010101000",
28379 => "0010000010101000",
28380 => "0010000010101000",
28381 => "0010000010101000",
28382 => "0010000010110000",
28383 => "0010000010110000",
28384 => "0010000010110000",
28385 => "0010000010110000",
28386 => "0010000010110000",
28387 => "0010000010111000",
28388 => "0010000010111000",
28389 => "0010000010111000",
28390 => "0010000010111000",
28391 => "0010000010111000",
28392 => "0010000010111000",
28393 => "0010000011000000",
28394 => "0010000011000000",
28395 => "0010000011000000",
28396 => "0010000011000000",
28397 => "0010000011000000",
28398 => "0010000011001000",
28399 => "0010000011001000",
28400 => "0010000011001000",
28401 => "0010000011001000",
28402 => "0010000011001000",
28403 => "0010000011010000",
28404 => "0010000011010000",
28405 => "0010000011010000",
28406 => "0010000011010000",
28407 => "0010000011010000",
28408 => "0010000011011000",
28409 => "0010000011011000",
28410 => "0010000011011000",
28411 => "0010000011011000",
28412 => "0010000011011000",
28413 => "0010000011011000",
28414 => "0010000011100000",
28415 => "0010000011100000",
28416 => "0010000011100000",
28417 => "0010000011100000",
28418 => "0010000011100000",
28419 => "0010000011101000",
28420 => "0010000011101000",
28421 => "0010000011101000",
28422 => "0010000011101000",
28423 => "0010000011101000",
28424 => "0010000011110000",
28425 => "0010000011110000",
28426 => "0010000011110000",
28427 => "0010000011110000",
28428 => "0010000011110000",
28429 => "0010000011111000",
28430 => "0010000011111000",
28431 => "0010000011111000",
28432 => "0010000011111000",
28433 => "0010000011111000",
28434 => "0010000100000000",
28435 => "0010000100000000",
28436 => "0010000100000000",
28437 => "0010000100000000",
28438 => "0010000100000000",
28439 => "0010000100000000",
28440 => "0010000100001000",
28441 => "0010000100001000",
28442 => "0010000100001000",
28443 => "0010000100001000",
28444 => "0010000100001000",
28445 => "0010000100010000",
28446 => "0010000100010000",
28447 => "0010000100010000",
28448 => "0010000100010000",
28449 => "0010000100010000",
28450 => "0010000100011000",
28451 => "0010000100011000",
28452 => "0010000100011000",
28453 => "0010000100011000",
28454 => "0010000100011000",
28455 => "0010000100100000",
28456 => "0010000100100000",
28457 => "0010000100100000",
28458 => "0010000100100000",
28459 => "0010000100100000",
28460 => "0010000100100000",
28461 => "0010000100101000",
28462 => "0010000100101000",
28463 => "0010000100101000",
28464 => "0010000100101000",
28465 => "0010000100101000",
28466 => "0010000100110000",
28467 => "0010000100110000",
28468 => "0010000100110000",
28469 => "0010000100110000",
28470 => "0010000100110000",
28471 => "0010000100111000",
28472 => "0010000100111000",
28473 => "0010000100111000",
28474 => "0010000100111000",
28475 => "0010000100111000",
28476 => "0010000101000000",
28477 => "0010000101000000",
28478 => "0010000101000000",
28479 => "0010000101000000",
28480 => "0010000101000000",
28481 => "0010000101001000",
28482 => "0010000101001000",
28483 => "0010000101001000",
28484 => "0010000101001000",
28485 => "0010000101001000",
28486 => "0010000101001000",
28487 => "0010000101010000",
28488 => "0010000101010000",
28489 => "0010000101010000",
28490 => "0010000101010000",
28491 => "0010000101010000",
28492 => "0010000101011000",
28493 => "0010000101011000",
28494 => "0010000101011000",
28495 => "0010000101011000",
28496 => "0010000101011000",
28497 => "0010000101100000",
28498 => "0010000101100000",
28499 => "0010000101100000",
28500 => "0010000101100000",
28501 => "0010000101100000",
28502 => "0010000101101000",
28503 => "0010000101101000",
28504 => "0010000101101000",
28505 => "0010000101101000",
28506 => "0010000101101000",
28507 => "0010000101110000",
28508 => "0010000101110000",
28509 => "0010000101110000",
28510 => "0010000101110000",
28511 => "0010000101110000",
28512 => "0010000101110000",
28513 => "0010000101111000",
28514 => "0010000101111000",
28515 => "0010000101111000",
28516 => "0010000101111000",
28517 => "0010000101111000",
28518 => "0010000110000000",
28519 => "0010000110000000",
28520 => "0010000110000000",
28521 => "0010000110000000",
28522 => "0010000110000000",
28523 => "0010000110001000",
28524 => "0010000110001000",
28525 => "0010000110001000",
28526 => "0010000110001000",
28527 => "0010000110001000",
28528 => "0010000110010000",
28529 => "0010000110010000",
28530 => "0010000110010000",
28531 => "0010000110010000",
28532 => "0010000110010000",
28533 => "0010000110011000",
28534 => "0010000110011000",
28535 => "0010000110011000",
28536 => "0010000110011000",
28537 => "0010000110011000",
28538 => "0010000110100000",
28539 => "0010000110100000",
28540 => "0010000110100000",
28541 => "0010000110100000",
28542 => "0010000110100000",
28543 => "0010000110100000",
28544 => "0010000110101000",
28545 => "0010000110101000",
28546 => "0010000110101000",
28547 => "0010000110101000",
28548 => "0010000110101000",
28549 => "0010000110110000",
28550 => "0010000110110000",
28551 => "0010000110110000",
28552 => "0010000110110000",
28553 => "0010000110110000",
28554 => "0010000110111000",
28555 => "0010000110111000",
28556 => "0010000110111000",
28557 => "0010000110111000",
28558 => "0010000110111000",
28559 => "0010000111000000",
28560 => "0010000111000000",
28561 => "0010000111000000",
28562 => "0010000111000000",
28563 => "0010000111000000",
28564 => "0010000111001000",
28565 => "0010000111001000",
28566 => "0010000111001000",
28567 => "0010000111001000",
28568 => "0010000111001000",
28569 => "0010000111010000",
28570 => "0010000111010000",
28571 => "0010000111010000",
28572 => "0010000111010000",
28573 => "0010000111010000",
28574 => "0010000111011000",
28575 => "0010000111011000",
28576 => "0010000111011000",
28577 => "0010000111011000",
28578 => "0010000111011000",
28579 => "0010000111011000",
28580 => "0010000111100000",
28581 => "0010000111100000",
28582 => "0010000111100000",
28583 => "0010000111100000",
28584 => "0010000111100000",
28585 => "0010000111101000",
28586 => "0010000111101000",
28587 => "0010000111101000",
28588 => "0010000111101000",
28589 => "0010000111101000",
28590 => "0010000111110000",
28591 => "0010000111110000",
28592 => "0010000111110000",
28593 => "0010000111110000",
28594 => "0010000111110000",
28595 => "0010000111111000",
28596 => "0010000111111000",
28597 => "0010000111111000",
28598 => "0010000111111000",
28599 => "0010000111111000",
28600 => "0010001000000000",
28601 => "0010001000000000",
28602 => "0010001000000000",
28603 => "0010001000000000",
28604 => "0010001000000000",
28605 => "0010001000001000",
28606 => "0010001000001000",
28607 => "0010001000001000",
28608 => "0010001000001000",
28609 => "0010001000001000",
28610 => "0010001000010000",
28611 => "0010001000010000",
28612 => "0010001000010000",
28613 => "0010001000010000",
28614 => "0010001000010000",
28615 => "0010001000010000",
28616 => "0010001000011000",
28617 => "0010001000011000",
28618 => "0010001000011000",
28619 => "0010001000011000",
28620 => "0010001000011000",
28621 => "0010001000100000",
28622 => "0010001000100000",
28623 => "0010001000100000",
28624 => "0010001000100000",
28625 => "0010001000100000",
28626 => "0010001000101000",
28627 => "0010001000101000",
28628 => "0010001000101000",
28629 => "0010001000101000",
28630 => "0010001000101000",
28631 => "0010001000110000",
28632 => "0010001000110000",
28633 => "0010001000110000",
28634 => "0010001000110000",
28635 => "0010001000110000",
28636 => "0010001000111000",
28637 => "0010001000111000",
28638 => "0010001000111000",
28639 => "0010001000111000",
28640 => "0010001000111000",
28641 => "0010001001000000",
28642 => "0010001001000000",
28643 => "0010001001000000",
28644 => "0010001001000000",
28645 => "0010001001000000",
28646 => "0010001001001000",
28647 => "0010001001001000",
28648 => "0010001001001000",
28649 => "0010001001001000",
28650 => "0010001001001000",
28651 => "0010001001010000",
28652 => "0010001001010000",
28653 => "0010001001010000",
28654 => "0010001001010000",
28655 => "0010001001010000",
28656 => "0010001001011000",
28657 => "0010001001011000",
28658 => "0010001001011000",
28659 => "0010001001011000",
28660 => "0010001001011000",
28661 => "0010001001100000",
28662 => "0010001001100000",
28663 => "0010001001100000",
28664 => "0010001001100000",
28665 => "0010001001100000",
28666 => "0010001001100000",
28667 => "0010001001101000",
28668 => "0010001001101000",
28669 => "0010001001101000",
28670 => "0010001001101000",
28671 => "0010001001101000",
28672 => "0010001001110000",
28673 => "0010001001110000",
28674 => "0010001001110000",
28675 => "0010001001110000",
28676 => "0010001001110000",
28677 => "0010001001111000",
28678 => "0010001001111000",
28679 => "0010001001111000",
28680 => "0010001001111000",
28681 => "0010001001111000",
28682 => "0010001010000000",
28683 => "0010001010000000",
28684 => "0010001010000000",
28685 => "0010001010000000",
28686 => "0010001010000000",
28687 => "0010001010001000",
28688 => "0010001010001000",
28689 => "0010001010001000",
28690 => "0010001010001000",
28691 => "0010001010001000",
28692 => "0010001010010000",
28693 => "0010001010010000",
28694 => "0010001010010000",
28695 => "0010001010010000",
28696 => "0010001010010000",
28697 => "0010001010011000",
28698 => "0010001010011000",
28699 => "0010001010011000",
28700 => "0010001010011000",
28701 => "0010001010011000",
28702 => "0010001010100000",
28703 => "0010001010100000",
28704 => "0010001010100000",
28705 => "0010001010100000",
28706 => "0010001010100000",
28707 => "0010001010101000",
28708 => "0010001010101000",
28709 => "0010001010101000",
28710 => "0010001010101000",
28711 => "0010001010101000",
28712 => "0010001010110000",
28713 => "0010001010110000",
28714 => "0010001010110000",
28715 => "0010001010110000",
28716 => "0010001010110000",
28717 => "0010001010111000",
28718 => "0010001010111000",
28719 => "0010001010111000",
28720 => "0010001010111000",
28721 => "0010001010111000",
28722 => "0010001011000000",
28723 => "0010001011000000",
28724 => "0010001011000000",
28725 => "0010001011000000",
28726 => "0010001011000000",
28727 => "0010001011001000",
28728 => "0010001011001000",
28729 => "0010001011001000",
28730 => "0010001011001000",
28731 => "0010001011001000",
28732 => "0010001011010000",
28733 => "0010001011010000",
28734 => "0010001011010000",
28735 => "0010001011010000",
28736 => "0010001011010000",
28737 => "0010001011010000",
28738 => "0010001011011000",
28739 => "0010001011011000",
28740 => "0010001011011000",
28741 => "0010001011011000",
28742 => "0010001011011000",
28743 => "0010001011100000",
28744 => "0010001011100000",
28745 => "0010001011100000",
28746 => "0010001011100000",
28747 => "0010001011100000",
28748 => "0010001011101000",
28749 => "0010001011101000",
28750 => "0010001011101000",
28751 => "0010001011101000",
28752 => "0010001011101000",
28753 => "0010001011110000",
28754 => "0010001011110000",
28755 => "0010001011110000",
28756 => "0010001011110000",
28757 => "0010001011110000",
28758 => "0010001011111000",
28759 => "0010001011111000",
28760 => "0010001011111000",
28761 => "0010001011111000",
28762 => "0010001011111000",
28763 => "0010001100000000",
28764 => "0010001100000000",
28765 => "0010001100000000",
28766 => "0010001100000000",
28767 => "0010001100000000",
28768 => "0010001100001000",
28769 => "0010001100001000",
28770 => "0010001100001000",
28771 => "0010001100001000",
28772 => "0010001100001000",
28773 => "0010001100010000",
28774 => "0010001100010000",
28775 => "0010001100010000",
28776 => "0010001100010000",
28777 => "0010001100010000",
28778 => "0010001100011000",
28779 => "0010001100011000",
28780 => "0010001100011000",
28781 => "0010001100011000",
28782 => "0010001100011000",
28783 => "0010001100100000",
28784 => "0010001100100000",
28785 => "0010001100100000",
28786 => "0010001100100000",
28787 => "0010001100100000",
28788 => "0010001100101000",
28789 => "0010001100101000",
28790 => "0010001100101000",
28791 => "0010001100101000",
28792 => "0010001100101000",
28793 => "0010001100110000",
28794 => "0010001100110000",
28795 => "0010001100110000",
28796 => "0010001100110000",
28797 => "0010001100110000",
28798 => "0010001100111000",
28799 => "0010001100111000",
28800 => "0010001100111000",
28801 => "0010001100111000",
28802 => "0010001100111000",
28803 => "0010001101000000",
28804 => "0010001101000000",
28805 => "0010001101000000",
28806 => "0010001101000000",
28807 => "0010001101000000",
28808 => "0010001101001000",
28809 => "0010001101001000",
28810 => "0010001101001000",
28811 => "0010001101001000",
28812 => "0010001101001000",
28813 => "0010001101010000",
28814 => "0010001101010000",
28815 => "0010001101010000",
28816 => "0010001101010000",
28817 => "0010001101010000",
28818 => "0010001101011000",
28819 => "0010001101011000",
28820 => "0010001101011000",
28821 => "0010001101011000",
28822 => "0010001101011000",
28823 => "0010001101100000",
28824 => "0010001101100000",
28825 => "0010001101100000",
28826 => "0010001101100000",
28827 => "0010001101100000",
28828 => "0010001101101000",
28829 => "0010001101101000",
28830 => "0010001101101000",
28831 => "0010001101101000",
28832 => "0010001101101000",
28833 => "0010001101110000",
28834 => "0010001101110000",
28835 => "0010001101110000",
28836 => "0010001101110000",
28837 => "0010001101110000",
28838 => "0010001101111000",
28839 => "0010001101111000",
28840 => "0010001101111000",
28841 => "0010001101111000",
28842 => "0010001101111000",
28843 => "0010001110000000",
28844 => "0010001110000000",
28845 => "0010001110000000",
28846 => "0010001110000000",
28847 => "0010001110000000",
28848 => "0010001110001000",
28849 => "0010001110001000",
28850 => "0010001110001000",
28851 => "0010001110001000",
28852 => "0010001110001000",
28853 => "0010001110010000",
28854 => "0010001110010000",
28855 => "0010001110010000",
28856 => "0010001110010000",
28857 => "0010001110010000",
28858 => "0010001110011000",
28859 => "0010001110011000",
28860 => "0010001110011000",
28861 => "0010001110011000",
28862 => "0010001110011000",
28863 => "0010001110100000",
28864 => "0010001110100000",
28865 => "0010001110100000",
28866 => "0010001110100000",
28867 => "0010001110100000",
28868 => "0010001110101000",
28869 => "0010001110101000",
28870 => "0010001110101000",
28871 => "0010001110101000",
28872 => "0010001110101000",
28873 => "0010001110110000",
28874 => "0010001110110000",
28875 => "0010001110110000",
28876 => "0010001110110000",
28877 => "0010001110110000",
28878 => "0010001110111000",
28879 => "0010001110111000",
28880 => "0010001110111000",
28881 => "0010001110111000",
28882 => "0010001110111000",
28883 => "0010001111000000",
28884 => "0010001111000000",
28885 => "0010001111000000",
28886 => "0010001111000000",
28887 => "0010001111000000",
28888 => "0010001111001000",
28889 => "0010001111001000",
28890 => "0010001111001000",
28891 => "0010001111001000",
28892 => "0010001111001000",
28893 => "0010001111010000",
28894 => "0010001111010000",
28895 => "0010001111010000",
28896 => "0010001111010000",
28897 => "0010001111010000",
28898 => "0010001111011000",
28899 => "0010001111011000",
28900 => "0010001111011000",
28901 => "0010001111011000",
28902 => "0010001111011000",
28903 => "0010001111100000",
28904 => "0010001111100000",
28905 => "0010001111100000",
28906 => "0010001111100000",
28907 => "0010001111100000",
28908 => "0010001111101000",
28909 => "0010001111101000",
28910 => "0010001111101000",
28911 => "0010001111101000",
28912 => "0010001111101000",
28913 => "0010001111110000",
28914 => "0010001111110000",
28915 => "0010001111110000",
28916 => "0010001111110000",
28917 => "0010001111111000",
28918 => "0010001111111000",
28919 => "0010001111111000",
28920 => "0010001111111000",
28921 => "0010001111111000",
28922 => "0010010000000000",
28923 => "0010010000000000",
28924 => "0010010000000000",
28925 => "0010010000000000",
28926 => "0010010000000000",
28927 => "0010010000001000",
28928 => "0010010000001000",
28929 => "0010010000001000",
28930 => "0010010000001000",
28931 => "0010010000001000",
28932 => "0010010000010000",
28933 => "0010010000010000",
28934 => "0010010000010000",
28935 => "0010010000010000",
28936 => "0010010000010000",
28937 => "0010010000011000",
28938 => "0010010000011000",
28939 => "0010010000011000",
28940 => "0010010000011000",
28941 => "0010010000011000",
28942 => "0010010000100000",
28943 => "0010010000100000",
28944 => "0010010000100000",
28945 => "0010010000100000",
28946 => "0010010000100000",
28947 => "0010010000101000",
28948 => "0010010000101000",
28949 => "0010010000101000",
28950 => "0010010000101000",
28951 => "0010010000101000",
28952 => "0010010000110000",
28953 => "0010010000110000",
28954 => "0010010000110000",
28955 => "0010010000110000",
28956 => "0010010000110000",
28957 => "0010010000111000",
28958 => "0010010000111000",
28959 => "0010010000111000",
28960 => "0010010000111000",
28961 => "0010010000111000",
28962 => "0010010001000000",
28963 => "0010010001000000",
28964 => "0010010001000000",
28965 => "0010010001000000",
28966 => "0010010001000000",
28967 => "0010010001001000",
28968 => "0010010001001000",
28969 => "0010010001001000",
28970 => "0010010001001000",
28971 => "0010010001001000",
28972 => "0010010001010000",
28973 => "0010010001010000",
28974 => "0010010001010000",
28975 => "0010010001010000",
28976 => "0010010001010000",
28977 => "0010010001011000",
28978 => "0010010001011000",
28979 => "0010010001011000",
28980 => "0010010001011000",
28981 => "0010010001011000",
28982 => "0010010001100000",
28983 => "0010010001100000",
28984 => "0010010001100000",
28985 => "0010010001100000",
28986 => "0010010001100000",
28987 => "0010010001101000",
28988 => "0010010001101000",
28989 => "0010010001101000",
28990 => "0010010001101000",
28991 => "0010010001110000",
28992 => "0010010001110000",
28993 => "0010010001110000",
28994 => "0010010001110000",
28995 => "0010010001110000",
28996 => "0010010001111000",
28997 => "0010010001111000",
28998 => "0010010001111000",
28999 => "0010010001111000",
29000 => "0010010001111000",
29001 => "0010010010000000",
29002 => "0010010010000000",
29003 => "0010010010000000",
29004 => "0010010010000000",
29005 => "0010010010000000",
29006 => "0010010010001000",
29007 => "0010010010001000",
29008 => "0010010010001000",
29009 => "0010010010001000",
29010 => "0010010010001000",
29011 => "0010010010010000",
29012 => "0010010010010000",
29013 => "0010010010010000",
29014 => "0010010010010000",
29015 => "0010010010010000",
29016 => "0010010010011000",
29017 => "0010010010011000",
29018 => "0010010010011000",
29019 => "0010010010011000",
29020 => "0010010010011000",
29021 => "0010010010100000",
29022 => "0010010010100000",
29023 => "0010010010100000",
29024 => "0010010010100000",
29025 => "0010010010100000",
29026 => "0010010010101000",
29027 => "0010010010101000",
29028 => "0010010010101000",
29029 => "0010010010101000",
29030 => "0010010010101000",
29031 => "0010010010110000",
29032 => "0010010010110000",
29033 => "0010010010110000",
29034 => "0010010010110000",
29035 => "0010010010110000",
29036 => "0010010010111000",
29037 => "0010010010111000",
29038 => "0010010010111000",
29039 => "0010010010111000",
29040 => "0010010011000000",
29041 => "0010010011000000",
29042 => "0010010011000000",
29043 => "0010010011000000",
29044 => "0010010011000000",
29045 => "0010010011001000",
29046 => "0010010011001000",
29047 => "0010010011001000",
29048 => "0010010011001000",
29049 => "0010010011001000",
29050 => "0010010011010000",
29051 => "0010010011010000",
29052 => "0010010011010000",
29053 => "0010010011010000",
29054 => "0010010011010000",
29055 => "0010010011011000",
29056 => "0010010011011000",
29057 => "0010010011011000",
29058 => "0010010011011000",
29059 => "0010010011011000",
29060 => "0010010011100000",
29061 => "0010010011100000",
29062 => "0010010011100000",
29063 => "0010010011100000",
29064 => "0010010011100000",
29065 => "0010010011101000",
29066 => "0010010011101000",
29067 => "0010010011101000",
29068 => "0010010011101000",
29069 => "0010010011101000",
29070 => "0010010011110000",
29071 => "0010010011110000",
29072 => "0010010011110000",
29073 => "0010010011110000",
29074 => "0010010011110000",
29075 => "0010010011111000",
29076 => "0010010011111000",
29077 => "0010010011111000",
29078 => "0010010011111000",
29079 => "0010010100000000",
29080 => "0010010100000000",
29081 => "0010010100000000",
29082 => "0010010100000000",
29083 => "0010010100000000",
29084 => "0010010100001000",
29085 => "0010010100001000",
29086 => "0010010100001000",
29087 => "0010010100001000",
29088 => "0010010100001000",
29089 => "0010010100010000",
29090 => "0010010100010000",
29091 => "0010010100010000",
29092 => "0010010100010000",
29093 => "0010010100010000",
29094 => "0010010100011000",
29095 => "0010010100011000",
29096 => "0010010100011000",
29097 => "0010010100011000",
29098 => "0010010100011000",
29099 => "0010010100100000",
29100 => "0010010100100000",
29101 => "0010010100100000",
29102 => "0010010100100000",
29103 => "0010010100100000",
29104 => "0010010100101000",
29105 => "0010010100101000",
29106 => "0010010100101000",
29107 => "0010010100101000",
29108 => "0010010100101000",
29109 => "0010010100110000",
29110 => "0010010100110000",
29111 => "0010010100110000",
29112 => "0010010100110000",
29113 => "0010010100111000",
29114 => "0010010100111000",
29115 => "0010010100111000",
29116 => "0010010100111000",
29117 => "0010010100111000",
29118 => "0010010101000000",
29119 => "0010010101000000",
29120 => "0010010101000000",
29121 => "0010010101000000",
29122 => "0010010101000000",
29123 => "0010010101001000",
29124 => "0010010101001000",
29125 => "0010010101001000",
29126 => "0010010101001000",
29127 => "0010010101001000",
29128 => "0010010101010000",
29129 => "0010010101010000",
29130 => "0010010101010000",
29131 => "0010010101010000",
29132 => "0010010101010000",
29133 => "0010010101011000",
29134 => "0010010101011000",
29135 => "0010010101011000",
29136 => "0010010101011000",
29137 => "0010010101011000",
29138 => "0010010101100000",
29139 => "0010010101100000",
29140 => "0010010101100000",
29141 => "0010010101100000",
29142 => "0010010101100000",
29143 => "0010010101101000",
29144 => "0010010101101000",
29145 => "0010010101101000",
29146 => "0010010101101000",
29147 => "0010010101110000",
29148 => "0010010101110000",
29149 => "0010010101110000",
29150 => "0010010101110000",
29151 => "0010010101110000",
29152 => "0010010101111000",
29153 => "0010010101111000",
29154 => "0010010101111000",
29155 => "0010010101111000",
29156 => "0010010101111000",
29157 => "0010010110000000",
29158 => "0010010110000000",
29159 => "0010010110000000",
29160 => "0010010110000000",
29161 => "0010010110000000",
29162 => "0010010110001000",
29163 => "0010010110001000",
29164 => "0010010110001000",
29165 => "0010010110001000",
29166 => "0010010110001000",
29167 => "0010010110010000",
29168 => "0010010110010000",
29169 => "0010010110010000",
29170 => "0010010110010000",
29171 => "0010010110010000",
29172 => "0010010110011000",
29173 => "0010010110011000",
29174 => "0010010110011000",
29175 => "0010010110011000",
29176 => "0010010110100000",
29177 => "0010010110100000",
29178 => "0010010110100000",
29179 => "0010010110100000",
29180 => "0010010110100000",
29181 => "0010010110101000",
29182 => "0010010110101000",
29183 => "0010010110101000",
29184 => "0010010110101000",
29185 => "0010010110101000",
29186 => "0010010110110000",
29187 => "0010010110110000",
29188 => "0010010110110000",
29189 => "0010010110110000",
29190 => "0010010110110000",
29191 => "0010010110111000",
29192 => "0010010110111000",
29193 => "0010010110111000",
29194 => "0010010110111000",
29195 => "0010010110111000",
29196 => "0010010111000000",
29197 => "0010010111000000",
29198 => "0010010111000000",
29199 => "0010010111000000",
29200 => "0010010111001000",
29201 => "0010010111001000",
29202 => "0010010111001000",
29203 => "0010010111001000",
29204 => "0010010111001000",
29205 => "0010010111010000",
29206 => "0010010111010000",
29207 => "0010010111010000",
29208 => "0010010111010000",
29209 => "0010010111010000",
29210 => "0010010111011000",
29211 => "0010010111011000",
29212 => "0010010111011000",
29213 => "0010010111011000",
29214 => "0010010111011000",
29215 => "0010010111100000",
29216 => "0010010111100000",
29217 => "0010010111100000",
29218 => "0010010111100000",
29219 => "0010010111100000",
29220 => "0010010111101000",
29221 => "0010010111101000",
29222 => "0010010111101000",
29223 => "0010010111101000",
29224 => "0010010111110000",
29225 => "0010010111110000",
29226 => "0010010111110000",
29227 => "0010010111110000",
29228 => "0010010111110000",
29229 => "0010010111111000",
29230 => "0010010111111000",
29231 => "0010010111111000",
29232 => "0010010111111000",
29233 => "0010010111111000",
29234 => "0010011000000000",
29235 => "0010011000000000",
29236 => "0010011000000000",
29237 => "0010011000000000",
29238 => "0010011000000000",
29239 => "0010011000001000",
29240 => "0010011000001000",
29241 => "0010011000001000",
29242 => "0010011000001000",
29243 => "0010011000001000",
29244 => "0010011000010000",
29245 => "0010011000010000",
29246 => "0010011000010000",
29247 => "0010011000010000",
29248 => "0010011000011000",
29249 => "0010011000011000",
29250 => "0010011000011000",
29251 => "0010011000011000",
29252 => "0010011000011000",
29253 => "0010011000100000",
29254 => "0010011000100000",
29255 => "0010011000100000",
29256 => "0010011000100000",
29257 => "0010011000100000",
29258 => "0010011000101000",
29259 => "0010011000101000",
29260 => "0010011000101000",
29261 => "0010011000101000",
29262 => "0010011000101000",
29263 => "0010011000110000",
29264 => "0010011000110000",
29265 => "0010011000110000",
29266 => "0010011000110000",
29267 => "0010011000111000",
29268 => "0010011000111000",
29269 => "0010011000111000",
29270 => "0010011000111000",
29271 => "0010011000111000",
29272 => "0010011001000000",
29273 => "0010011001000000",
29274 => "0010011001000000",
29275 => "0010011001000000",
29276 => "0010011001000000",
29277 => "0010011001001000",
29278 => "0010011001001000",
29279 => "0010011001001000",
29280 => "0010011001001000",
29281 => "0010011001001000",
29282 => "0010011001010000",
29283 => "0010011001010000",
29284 => "0010011001010000",
29285 => "0010011001010000",
29286 => "0010011001010000",
29287 => "0010011001011000",
29288 => "0010011001011000",
29289 => "0010011001011000",
29290 => "0010011001011000",
29291 => "0010011001100000",
29292 => "0010011001100000",
29293 => "0010011001100000",
29294 => "0010011001100000",
29295 => "0010011001100000",
29296 => "0010011001101000",
29297 => "0010011001101000",
29298 => "0010011001101000",
29299 => "0010011001101000",
29300 => "0010011001101000",
29301 => "0010011001110000",
29302 => "0010011001110000",
29303 => "0010011001110000",
29304 => "0010011001110000",
29305 => "0010011001110000",
29306 => "0010011001111000",
29307 => "0010011001111000",
29308 => "0010011001111000",
29309 => "0010011001111000",
29310 => "0010011010000000",
29311 => "0010011010000000",
29312 => "0010011010000000",
29313 => "0010011010000000",
29314 => "0010011010000000",
29315 => "0010011010001000",
29316 => "0010011010001000",
29317 => "0010011010001000",
29318 => "0010011010001000",
29319 => "0010011010001000",
29320 => "0010011010010000",
29321 => "0010011010010000",
29322 => "0010011010010000",
29323 => "0010011010010000",
29324 => "0010011010010000",
29325 => "0010011010011000",
29326 => "0010011010011000",
29327 => "0010011010011000",
29328 => "0010011010011000",
29329 => "0010011010100000",
29330 => "0010011010100000",
29331 => "0010011010100000",
29332 => "0010011010100000",
29333 => "0010011010100000",
29334 => "0010011010101000",
29335 => "0010011010101000",
29336 => "0010011010101000",
29337 => "0010011010101000",
29338 => "0010011010101000",
29339 => "0010011010110000",
29340 => "0010011010110000",
29341 => "0010011010110000",
29342 => "0010011010110000",
29343 => "0010011010110000",
29344 => "0010011010111000",
29345 => "0010011010111000",
29346 => "0010011010111000",
29347 => "0010011010111000",
29348 => "0010011011000000",
29349 => "0010011011000000",
29350 => "0010011011000000",
29351 => "0010011011000000",
29352 => "0010011011000000",
29353 => "0010011011001000",
29354 => "0010011011001000",
29355 => "0010011011001000",
29356 => "0010011011001000",
29357 => "0010011011001000",
29358 => "0010011011010000",
29359 => "0010011011010000",
29360 => "0010011011010000",
29361 => "0010011011010000",
29362 => "0010011011010000",
29363 => "0010011011011000",
29364 => "0010011011011000",
29365 => "0010011011011000",
29366 => "0010011011011000",
29367 => "0010011011100000",
29368 => "0010011011100000",
29369 => "0010011011100000",
29370 => "0010011011100000",
29371 => "0010011011100000",
29372 => "0010011011101000",
29373 => "0010011011101000",
29374 => "0010011011101000",
29375 => "0010011011101000",
29376 => "0010011011101000",
29377 => "0010011011110000",
29378 => "0010011011110000",
29379 => "0010011011110000",
29380 => "0010011011110000",
29381 => "0010011011111000",
29382 => "0010011011111000",
29383 => "0010011011111000",
29384 => "0010011011111000",
29385 => "0010011011111000",
29386 => "0010011100000000",
29387 => "0010011100000000",
29388 => "0010011100000000",
29389 => "0010011100000000",
29390 => "0010011100000000",
29391 => "0010011100001000",
29392 => "0010011100001000",
29393 => "0010011100001000",
29394 => "0010011100001000",
29395 => "0010011100001000",
29396 => "0010011100010000",
29397 => "0010011100010000",
29398 => "0010011100010000",
29399 => "0010011100010000",
29400 => "0010011100011000",
29401 => "0010011100011000",
29402 => "0010011100011000",
29403 => "0010011100011000",
29404 => "0010011100011000",
29405 => "0010011100100000",
29406 => "0010011100100000",
29407 => "0010011100100000",
29408 => "0010011100100000",
29409 => "0010011100100000",
29410 => "0010011100101000",
29411 => "0010011100101000",
29412 => "0010011100101000",
29413 => "0010011100101000",
29414 => "0010011100110000",
29415 => "0010011100110000",
29416 => "0010011100110000",
29417 => "0010011100110000",
29418 => "0010011100110000",
29419 => "0010011100111000",
29420 => "0010011100111000",
29421 => "0010011100111000",
29422 => "0010011100111000",
29423 => "0010011100111000",
29424 => "0010011101000000",
29425 => "0010011101000000",
29426 => "0010011101000000",
29427 => "0010011101000000",
29428 => "0010011101000000",
29429 => "0010011101001000",
29430 => "0010011101001000",
29431 => "0010011101001000",
29432 => "0010011101001000",
29433 => "0010011101010000",
29434 => "0010011101010000",
29435 => "0010011101010000",
29436 => "0010011101010000",
29437 => "0010011101010000",
29438 => "0010011101011000",
29439 => "0010011101011000",
29440 => "0010011101011000",
29441 => "0010011101011000",
29442 => "0010011101011000",
29443 => "0010011101100000",
29444 => "0010011101100000",
29445 => "0010011101100000",
29446 => "0010011101100000",
29447 => "0010011101101000",
29448 => "0010011101101000",
29449 => "0010011101101000",
29450 => "0010011101101000",
29451 => "0010011101101000",
29452 => "0010011101110000",
29453 => "0010011101110000",
29454 => "0010011101110000",
29455 => "0010011101110000",
29456 => "0010011101110000",
29457 => "0010011101111000",
29458 => "0010011101111000",
29459 => "0010011101111000",
29460 => "0010011101111000",
29461 => "0010011110000000",
29462 => "0010011110000000",
29463 => "0010011110000000",
29464 => "0010011110000000",
29465 => "0010011110000000",
29466 => "0010011110001000",
29467 => "0010011110001000",
29468 => "0010011110001000",
29469 => "0010011110001000",
29470 => "0010011110001000",
29471 => "0010011110010000",
29472 => "0010011110010000",
29473 => "0010011110010000",
29474 => "0010011110010000",
29475 => "0010011110010000",
29476 => "0010011110011000",
29477 => "0010011110011000",
29478 => "0010011110011000",
29479 => "0010011110011000",
29480 => "0010011110100000",
29481 => "0010011110100000",
29482 => "0010011110100000",
29483 => "0010011110100000",
29484 => "0010011110100000",
29485 => "0010011110101000",
29486 => "0010011110101000",
29487 => "0010011110101000",
29488 => "0010011110101000",
29489 => "0010011110101000",
29490 => "0010011110110000",
29491 => "0010011110110000",
29492 => "0010011110110000",
29493 => "0010011110110000",
29494 => "0010011110111000",
29495 => "0010011110111000",
29496 => "0010011110111000",
29497 => "0010011110111000",
29498 => "0010011110111000",
29499 => "0010011111000000",
29500 => "0010011111000000",
29501 => "0010011111000000",
29502 => "0010011111000000",
29503 => "0010011111000000",
29504 => "0010011111001000",
29505 => "0010011111001000",
29506 => "0010011111001000",
29507 => "0010011111001000",
29508 => "0010011111010000",
29509 => "0010011111010000",
29510 => "0010011111010000",
29511 => "0010011111010000",
29512 => "0010011111010000",
29513 => "0010011111011000",
29514 => "0010011111011000",
29515 => "0010011111011000",
29516 => "0010011111011000",
29517 => "0010011111011000",
29518 => "0010011111100000",
29519 => "0010011111100000",
29520 => "0010011111100000",
29521 => "0010011111100000",
29522 => "0010011111101000",
29523 => "0010011111101000",
29524 => "0010011111101000",
29525 => "0010011111101000",
29526 => "0010011111101000",
29527 => "0010011111110000",
29528 => "0010011111110000",
29529 => "0010011111110000",
29530 => "0010011111110000",
29531 => "0010011111110000",
29532 => "0010011111111000",
29533 => "0010011111111000",
29534 => "0010011111111000",
29535 => "0010011111111000",
29536 => "0010100000000000",
29537 => "0010100000000000",
29538 => "0010100000000000",
29539 => "0010100000000000",
29540 => "0010100000000000",
29541 => "0010100000001000",
29542 => "0010100000001000",
29543 => "0010100000001000",
29544 => "0010100000001000",
29545 => "0010100000001000",
29546 => "0010100000010000",
29547 => "0010100000010000",
29548 => "0010100000010000",
29549 => "0010100000010000",
29550 => "0010100000011000",
29551 => "0010100000011000",
29552 => "0010100000011000",
29553 => "0010100000011000",
29554 => "0010100000011000",
29555 => "0010100000100000",
29556 => "0010100000100000",
29557 => "0010100000100000",
29558 => "0010100000100000",
29559 => "0010100000101000",
29560 => "0010100000101000",
29561 => "0010100000101000",
29562 => "0010100000101000",
29563 => "0010100000101000",
29564 => "0010100000110000",
29565 => "0010100000110000",
29566 => "0010100000110000",
29567 => "0010100000110000",
29568 => "0010100000110000",
29569 => "0010100000111000",
29570 => "0010100000111000",
29571 => "0010100000111000",
29572 => "0010100000111000",
29573 => "0010100001000000",
29574 => "0010100001000000",
29575 => "0010100001000000",
29576 => "0010100001000000",
29577 => "0010100001000000",
29578 => "0010100001001000",
29579 => "0010100001001000",
29580 => "0010100001001000",
29581 => "0010100001001000",
29582 => "0010100001001000",
29583 => "0010100001010000",
29584 => "0010100001010000",
29585 => "0010100001010000",
29586 => "0010100001010000",
29587 => "0010100001011000",
29588 => "0010100001011000",
29589 => "0010100001011000",
29590 => "0010100001011000",
29591 => "0010100001011000",
29592 => "0010100001100000",
29593 => "0010100001100000",
29594 => "0010100001100000",
29595 => "0010100001100000",
29596 => "0010100001100000",
29597 => "0010100001101000",
29598 => "0010100001101000",
29599 => "0010100001101000",
29600 => "0010100001101000",
29601 => "0010100001110000",
29602 => "0010100001110000",
29603 => "0010100001110000",
29604 => "0010100001110000",
29605 => "0010100001110000",
29606 => "0010100001111000",
29607 => "0010100001111000",
29608 => "0010100001111000",
29609 => "0010100001111000",
29610 => "0010100010000000",
29611 => "0010100010000000",
29612 => "0010100010000000",
29613 => "0010100010000000",
29614 => "0010100010000000",
29615 => "0010100010001000",
29616 => "0010100010001000",
29617 => "0010100010001000",
29618 => "0010100010001000",
29619 => "0010100010001000",
29620 => "0010100010010000",
29621 => "0010100010010000",
29622 => "0010100010010000",
29623 => "0010100010010000",
29624 => "0010100010011000",
29625 => "0010100010011000",
29626 => "0010100010011000",
29627 => "0010100010011000",
29628 => "0010100010011000",
29629 => "0010100010100000",
29630 => "0010100010100000",
29631 => "0010100010100000",
29632 => "0010100010100000",
29633 => "0010100010100000",
29634 => "0010100010101000",
29635 => "0010100010101000",
29636 => "0010100010101000",
29637 => "0010100010101000",
29638 => "0010100010110000",
29639 => "0010100010110000",
29640 => "0010100010110000",
29641 => "0010100010110000",
29642 => "0010100010110000",
29643 => "0010100010111000",
29644 => "0010100010111000",
29645 => "0010100010111000",
29646 => "0010100010111000",
29647 => "0010100011000000",
29648 => "0010100011000000",
29649 => "0010100011000000",
29650 => "0010100011000000",
29651 => "0010100011000000",
29652 => "0010100011001000",
29653 => "0010100011001000",
29654 => "0010100011001000",
29655 => "0010100011001000",
29656 => "0010100011001000",
29657 => "0010100011010000",
29658 => "0010100011010000",
29659 => "0010100011010000",
29660 => "0010100011010000",
29661 => "0010100011011000",
29662 => "0010100011011000",
29663 => "0010100011011000",
29664 => "0010100011011000",
29665 => "0010100011011000",
29666 => "0010100011100000",
29667 => "0010100011100000",
29668 => "0010100011100000",
29669 => "0010100011100000",
29670 => "0010100011101000",
29671 => "0010100011101000",
29672 => "0010100011101000",
29673 => "0010100011101000",
29674 => "0010100011101000",
29675 => "0010100011110000",
29676 => "0010100011110000",
29677 => "0010100011110000",
29678 => "0010100011110000",
29679 => "0010100011110000",
29680 => "0010100011111000",
29681 => "0010100011111000",
29682 => "0010100011111000",
29683 => "0010100011111000",
29684 => "0010100100000000",
29685 => "0010100100000000",
29686 => "0010100100000000",
29687 => "0010100100000000",
29688 => "0010100100000000",
29689 => "0010100100001000",
29690 => "0010100100001000",
29691 => "0010100100001000",
29692 => "0010100100001000",
29693 => "0010100100010000",
29694 => "0010100100010000",
29695 => "0010100100010000",
29696 => "0010100100010000",
29697 => "0010100100010000",
29698 => "0010100100011000",
29699 => "0010100100011000",
29700 => "0010100100011000",
29701 => "0010100100011000",
29702 => "0010100100011000",
29703 => "0010100100100000",
29704 => "0010100100100000",
29705 => "0010100100100000",
29706 => "0010100100100000",
29707 => "0010100100101000",
29708 => "0010100100101000",
29709 => "0010100100101000",
29710 => "0010100100101000",
29711 => "0010100100101000",
29712 => "0010100100110000",
29713 => "0010100100110000",
29714 => "0010100100110000",
29715 => "0010100100110000",
29716 => "0010100100111000",
29717 => "0010100100111000",
29718 => "0010100100111000",
29719 => "0010100100111000",
29720 => "0010100100111000",
29721 => "0010100101000000",
29722 => "0010100101000000",
29723 => "0010100101000000",
29724 => "0010100101000000",
29725 => "0010100101001000",
29726 => "0010100101001000",
29727 => "0010100101001000",
29728 => "0010100101001000",
29729 => "0010100101001000",
29730 => "0010100101010000",
29731 => "0010100101010000",
29732 => "0010100101010000",
29733 => "0010100101010000",
29734 => "0010100101010000",
29735 => "0010100101011000",
29736 => "0010100101011000",
29737 => "0010100101011000",
29738 => "0010100101011000",
29739 => "0010100101100000",
29740 => "0010100101100000",
29741 => "0010100101100000",
29742 => "0010100101100000",
29743 => "0010100101100000",
29744 => "0010100101101000",
29745 => "0010100101101000",
29746 => "0010100101101000",
29747 => "0010100101101000",
29748 => "0010100101110000",
29749 => "0010100101110000",
29750 => "0010100101110000",
29751 => "0010100101110000",
29752 => "0010100101110000",
29753 => "0010100101111000",
29754 => "0010100101111000",
29755 => "0010100101111000",
29756 => "0010100101111000",
29757 => "0010100110000000",
29758 => "0010100110000000",
29759 => "0010100110000000",
29760 => "0010100110000000",
29761 => "0010100110000000",
29762 => "0010100110001000",
29763 => "0010100110001000",
29764 => "0010100110001000",
29765 => "0010100110001000",
29766 => "0010100110001000",
29767 => "0010100110010000",
29768 => "0010100110010000",
29769 => "0010100110010000",
29770 => "0010100110010000",
29771 => "0010100110011000",
29772 => "0010100110011000",
29773 => "0010100110011000",
29774 => "0010100110011000",
29775 => "0010100110011000",
29776 => "0010100110100000",
29777 => "0010100110100000",
29778 => "0010100110100000",
29779 => "0010100110100000",
29780 => "0010100110101000",
29781 => "0010100110101000",
29782 => "0010100110101000",
29783 => "0010100110101000",
29784 => "0010100110101000",
29785 => "0010100110110000",
29786 => "0010100110110000",
29787 => "0010100110110000",
29788 => "0010100110110000",
29789 => "0010100110111000",
29790 => "0010100110111000",
29791 => "0010100110111000",
29792 => "0010100110111000",
29793 => "0010100110111000",
29794 => "0010100111000000",
29795 => "0010100111000000",
29796 => "0010100111000000",
29797 => "0010100111000000",
29798 => "0010100111001000",
29799 => "0010100111001000",
29800 => "0010100111001000",
29801 => "0010100111001000",
29802 => "0010100111001000",
29803 => "0010100111010000",
29804 => "0010100111010000",
29805 => "0010100111010000",
29806 => "0010100111010000",
29807 => "0010100111010000",
29808 => "0010100111011000",
29809 => "0010100111011000",
29810 => "0010100111011000",
29811 => "0010100111011000",
29812 => "0010100111100000",
29813 => "0010100111100000",
29814 => "0010100111100000",
29815 => "0010100111100000",
29816 => "0010100111100000",
29817 => "0010100111101000",
29818 => "0010100111101000",
29819 => "0010100111101000",
29820 => "0010100111101000",
29821 => "0010100111110000",
29822 => "0010100111110000",
29823 => "0010100111110000",
29824 => "0010100111110000",
29825 => "0010100111110000",
29826 => "0010100111111000",
29827 => "0010100111111000",
29828 => "0010100111111000",
29829 => "0010100111111000",
29830 => "0010101000000000",
29831 => "0010101000000000",
29832 => "0010101000000000",
29833 => "0010101000000000",
29834 => "0010101000000000",
29835 => "0010101000001000",
29836 => "0010101000001000",
29837 => "0010101000001000",
29838 => "0010101000001000",
29839 => "0010101000010000",
29840 => "0010101000010000",
29841 => "0010101000010000",
29842 => "0010101000010000",
29843 => "0010101000010000",
29844 => "0010101000011000",
29845 => "0010101000011000",
29846 => "0010101000011000",
29847 => "0010101000011000",
29848 => "0010101000100000",
29849 => "0010101000100000",
29850 => "0010101000100000",
29851 => "0010101000100000",
29852 => "0010101000100000",
29853 => "0010101000101000",
29854 => "0010101000101000",
29855 => "0010101000101000",
29856 => "0010101000101000",
29857 => "0010101000110000",
29858 => "0010101000110000",
29859 => "0010101000110000",
29860 => "0010101000110000",
29861 => "0010101000110000",
29862 => "0010101000111000",
29863 => "0010101000111000",
29864 => "0010101000111000",
29865 => "0010101000111000",
29866 => "0010101000111000",
29867 => "0010101001000000",
29868 => "0010101001000000",
29869 => "0010101001000000",
29870 => "0010101001000000",
29871 => "0010101001001000",
29872 => "0010101001001000",
29873 => "0010101001001000",
29874 => "0010101001001000",
29875 => "0010101001001000",
29876 => "0010101001010000",
29877 => "0010101001010000",
29878 => "0010101001010000",
29879 => "0010101001010000",
29880 => "0010101001011000",
29881 => "0010101001011000",
29882 => "0010101001011000",
29883 => "0010101001011000",
29884 => "0010101001011000",
29885 => "0010101001100000",
29886 => "0010101001100000",
29887 => "0010101001100000",
29888 => "0010101001100000",
29889 => "0010101001101000",
29890 => "0010101001101000",
29891 => "0010101001101000",
29892 => "0010101001101000",
29893 => "0010101001101000",
29894 => "0010101001110000",
29895 => "0010101001110000",
29896 => "0010101001110000",
29897 => "0010101001110000",
29898 => "0010101001111000",
29899 => "0010101001111000",
29900 => "0010101001111000",
29901 => "0010101001111000",
29902 => "0010101001111000",
29903 => "0010101010000000",
29904 => "0010101010000000",
29905 => "0010101010000000",
29906 => "0010101010000000",
29907 => "0010101010001000",
29908 => "0010101010001000",
29909 => "0010101010001000",
29910 => "0010101010001000",
29911 => "0010101010001000",
29912 => "0010101010010000",
29913 => "0010101010010000",
29914 => "0010101010010000",
29915 => "0010101010010000",
29916 => "0010101010011000",
29917 => "0010101010011000",
29918 => "0010101010011000",
29919 => "0010101010011000",
29920 => "0010101010011000",
29921 => "0010101010100000",
29922 => "0010101010100000",
29923 => "0010101010100000",
29924 => "0010101010100000",
29925 => "0010101010101000",
29926 => "0010101010101000",
29927 => "0010101010101000",
29928 => "0010101010101000",
29929 => "0010101010101000",
29930 => "0010101010110000",
29931 => "0010101010110000",
29932 => "0010101010110000",
29933 => "0010101010110000",
29934 => "0010101010111000",
29935 => "0010101010111000",
29936 => "0010101010111000",
29937 => "0010101010111000",
29938 => "0010101010111000",
29939 => "0010101011000000",
29940 => "0010101011000000",
29941 => "0010101011000000",
29942 => "0010101011000000",
29943 => "0010101011001000",
29944 => "0010101011001000",
29945 => "0010101011001000",
29946 => "0010101011001000",
29947 => "0010101011001000",
29948 => "0010101011010000",
29949 => "0010101011010000",
29950 => "0010101011010000",
29951 => "0010101011010000",
29952 => "0010101011011000",
29953 => "0010101011011000",
29954 => "0010101011011000",
29955 => "0010101011011000",
29956 => "0010101011011000",
29957 => "0010101011100000",
29958 => "0010101011100000",
29959 => "0010101011100000",
29960 => "0010101011100000",
29961 => "0010101011101000",
29962 => "0010101011101000",
29963 => "0010101011101000",
29964 => "0010101011101000",
29965 => "0010101011101000",
29966 => "0010101011110000",
29967 => "0010101011110000",
29968 => "0010101011110000",
29969 => "0010101011110000",
29970 => "0010101011111000",
29971 => "0010101011111000",
29972 => "0010101011111000",
29973 => "0010101011111000",
29974 => "0010101011111000",
29975 => "0010101100000000",
29976 => "0010101100000000",
29977 => "0010101100000000",
29978 => "0010101100000000",
29979 => "0010101100001000",
29980 => "0010101100001000",
29981 => "0010101100001000",
29982 => "0010101100001000",
29983 => "0010101100001000",
29984 => "0010101100010000",
29985 => "0010101100010000",
29986 => "0010101100010000",
29987 => "0010101100010000",
29988 => "0010101100011000",
29989 => "0010101100011000",
29990 => "0010101100011000",
29991 => "0010101100011000",
29992 => "0010101100100000",
29993 => "0010101100100000",
29994 => "0010101100100000",
29995 => "0010101100100000",
29996 => "0010101100100000",
29997 => "0010101100101000",
29998 => "0010101100101000",
29999 => "0010101100101000",
30000 => "0010101100101000",
30001 => "0010101100110000",
30002 => "0010101100110000",
30003 => "0010101100110000",
30004 => "0010101100110000",
30005 => "0010101100110000",
30006 => "0010101100111000",
30007 => "0010101100111000",
30008 => "0010101100111000",
30009 => "0010101100111000",
30010 => "0010101101000000",
30011 => "0010101101000000",
30012 => "0010101101000000",
30013 => "0010101101000000",
30014 => "0010101101000000",
30015 => "0010101101001000",
30016 => "0010101101001000",
30017 => "0010101101001000",
30018 => "0010101101001000",
30019 => "0010101101010000",
30020 => "0010101101010000",
30021 => "0010101101010000",
30022 => "0010101101010000",
30023 => "0010101101010000",
30024 => "0010101101011000",
30025 => "0010101101011000",
30026 => "0010101101011000",
30027 => "0010101101011000",
30028 => "0010101101100000",
30029 => "0010101101100000",
30030 => "0010101101100000",
30031 => "0010101101100000",
30032 => "0010101101100000",
30033 => "0010101101101000",
30034 => "0010101101101000",
30035 => "0010101101101000",
30036 => "0010101101101000",
30037 => "0010101101110000",
30038 => "0010101101110000",
30039 => "0010101101110000",
30040 => "0010101101110000",
30041 => "0010101101110000",
30042 => "0010101101111000",
30043 => "0010101101111000",
30044 => "0010101101111000",
30045 => "0010101101111000",
30046 => "0010101110000000",
30047 => "0010101110000000",
30048 => "0010101110000000",
30049 => "0010101110000000",
30050 => "0010101110000000",
30051 => "0010101110001000",
30052 => "0010101110001000",
30053 => "0010101110001000",
30054 => "0010101110001000",
30055 => "0010101110010000",
30056 => "0010101110010000",
30057 => "0010101110010000",
30058 => "0010101110010000",
30059 => "0010101110011000",
30060 => "0010101110011000",
30061 => "0010101110011000",
30062 => "0010101110011000",
30063 => "0010101110011000",
30064 => "0010101110100000",
30065 => "0010101110100000",
30066 => "0010101110100000",
30067 => "0010101110100000",
30068 => "0010101110101000",
30069 => "0010101110101000",
30070 => "0010101110101000",
30071 => "0010101110101000",
30072 => "0010101110101000",
30073 => "0010101110110000",
30074 => "0010101110110000",
30075 => "0010101110110000",
30076 => "0010101110110000",
30077 => "0010101110111000",
30078 => "0010101110111000",
30079 => "0010101110111000",
30080 => "0010101110111000",
30081 => "0010101110111000",
30082 => "0010101111000000",
30083 => "0010101111000000",
30084 => "0010101111000000",
30085 => "0010101111000000",
30086 => "0010101111001000",
30087 => "0010101111001000",
30088 => "0010101111001000",
30089 => "0010101111001000",
30090 => "0010101111001000",
30091 => "0010101111010000",
30092 => "0010101111010000",
30093 => "0010101111010000",
30094 => "0010101111010000",
30095 => "0010101111011000",
30096 => "0010101111011000",
30097 => "0010101111011000",
30098 => "0010101111011000",
30099 => "0010101111100000",
30100 => "0010101111100000",
30101 => "0010101111100000",
30102 => "0010101111100000",
30103 => "0010101111100000",
30104 => "0010101111101000",
30105 => "0010101111101000",
30106 => "0010101111101000",
30107 => "0010101111101000",
30108 => "0010101111110000",
30109 => "0010101111110000",
30110 => "0010101111110000",
30111 => "0010101111110000",
30112 => "0010101111110000",
30113 => "0010101111111000",
30114 => "0010101111111000",
30115 => "0010101111111000",
30116 => "0010101111111000",
30117 => "0010110000000000",
30118 => "0010110000000000",
30119 => "0010110000000000",
30120 => "0010110000000000",
30121 => "0010110000000000",
30122 => "0010110000001000",
30123 => "0010110000001000",
30124 => "0010110000001000",
30125 => "0010110000001000",
30126 => "0010110000010000",
30127 => "0010110000010000",
30128 => "0010110000010000",
30129 => "0010110000010000",
30130 => "0010110000010000",
30131 => "0010110000011000",
30132 => "0010110000011000",
30133 => "0010110000011000",
30134 => "0010110000011000",
30135 => "0010110000100000",
30136 => "0010110000100000",
30137 => "0010110000100000",
30138 => "0010110000100000",
30139 => "0010110000101000",
30140 => "0010110000101000",
30141 => "0010110000101000",
30142 => "0010110000101000",
30143 => "0010110000101000",
30144 => "0010110000110000",
30145 => "0010110000110000",
30146 => "0010110000110000",
30147 => "0010110000110000",
30148 => "0010110000111000",
30149 => "0010110000111000",
30150 => "0010110000111000",
30151 => "0010110000111000",
30152 => "0010110000111000",
30153 => "0010110001000000",
30154 => "0010110001000000",
30155 => "0010110001000000",
30156 => "0010110001000000",
30157 => "0010110001001000",
30158 => "0010110001001000",
30159 => "0010110001001000",
30160 => "0010110001001000",
30161 => "0010110001001000",
30162 => "0010110001010000",
30163 => "0010110001010000",
30164 => "0010110001010000",
30165 => "0010110001010000",
30166 => "0010110001011000",
30167 => "0010110001011000",
30168 => "0010110001011000",
30169 => "0010110001011000",
30170 => "0010110001100000",
30171 => "0010110001100000",
30172 => "0010110001100000",
30173 => "0010110001100000",
30174 => "0010110001100000",
30175 => "0010110001101000",
30176 => "0010110001101000",
30177 => "0010110001101000",
30178 => "0010110001101000",
30179 => "0010110001110000",
30180 => "0010110001110000",
30181 => "0010110001110000",
30182 => "0010110001110000",
30183 => "0010110001110000",
30184 => "0010110001111000",
30185 => "0010110001111000",
30186 => "0010110001111000",
30187 => "0010110001111000",
30188 => "0010110010000000",
30189 => "0010110010000000",
30190 => "0010110010000000",
30191 => "0010110010000000",
30192 => "0010110010001000",
30193 => "0010110010001000",
30194 => "0010110010001000",
30195 => "0010110010001000",
30196 => "0010110010001000",
30197 => "0010110010010000",
30198 => "0010110010010000",
30199 => "0010110010010000",
30200 => "0010110010010000",
30201 => "0010110010011000",
30202 => "0010110010011000",
30203 => "0010110010011000",
30204 => "0010110010011000",
30205 => "0010110010011000",
30206 => "0010110010100000",
30207 => "0010110010100000",
30208 => "0010110010100000",
30209 => "0010110010100000",
30210 => "0010110010101000",
30211 => "0010110010101000",
30212 => "0010110010101000",
30213 => "0010110010101000",
30214 => "0010110010110000",
30215 => "0010110010110000",
30216 => "0010110010110000",
30217 => "0010110010110000",
30218 => "0010110010110000",
30219 => "0010110010111000",
30220 => "0010110010111000",
30221 => "0010110010111000",
30222 => "0010110010111000",
30223 => "0010110011000000",
30224 => "0010110011000000",
30225 => "0010110011000000",
30226 => "0010110011000000",
30227 => "0010110011000000",
30228 => "0010110011001000",
30229 => "0010110011001000",
30230 => "0010110011001000",
30231 => "0010110011001000",
30232 => "0010110011010000",
30233 => "0010110011010000",
30234 => "0010110011010000",
30235 => "0010110011010000",
30236 => "0010110011011000",
30237 => "0010110011011000",
30238 => "0010110011011000",
30239 => "0010110011011000",
30240 => "0010110011011000",
30241 => "0010110011100000",
30242 => "0010110011100000",
30243 => "0010110011100000",
30244 => "0010110011100000",
30245 => "0010110011101000",
30246 => "0010110011101000",
30247 => "0010110011101000",
30248 => "0010110011101000",
30249 => "0010110011101000",
30250 => "0010110011110000",
30251 => "0010110011110000",
30252 => "0010110011110000",
30253 => "0010110011110000",
30254 => "0010110011111000",
30255 => "0010110011111000",
30256 => "0010110011111000",
30257 => "0010110011111000",
30258 => "0010110100000000",
30259 => "0010110100000000",
30260 => "0010110100000000",
30261 => "0010110100000000",
30262 => "0010110100000000",
30263 => "0010110100001000",
30264 => "0010110100001000",
30265 => "0010110100001000",
30266 => "0010110100001000",
30267 => "0010110100010000",
30268 => "0010110100010000",
30269 => "0010110100010000",
30270 => "0010110100010000",
30271 => "0010110100010000",
30272 => "0010110100011000",
30273 => "0010110100011000",
30274 => "0010110100011000",
30275 => "0010110100011000",
30276 => "0010110100100000",
30277 => "0010110100100000",
30278 => "0010110100100000",
30279 => "0010110100100000",
30280 => "0010110100101000",
30281 => "0010110100101000",
30282 => "0010110100101000",
30283 => "0010110100101000",
30284 => "0010110100101000",
30285 => "0010110100110000",
30286 => "0010110100110000",
30287 => "0010110100110000",
30288 => "0010110100110000",
30289 => "0010110100111000",
30290 => "0010110100111000",
30291 => "0010110100111000",
30292 => "0010110100111000",
30293 => "0010110101000000",
30294 => "0010110101000000",
30295 => "0010110101000000",
30296 => "0010110101000000",
30297 => "0010110101000000",
30298 => "0010110101001000",
30299 => "0010110101001000",
30300 => "0010110101001000",
30301 => "0010110101001000",
30302 => "0010110101010000",
30303 => "0010110101010000",
30304 => "0010110101010000",
30305 => "0010110101010000",
30306 => "0010110101010000",
30307 => "0010110101011000",
30308 => "0010110101011000",
30309 => "0010110101011000",
30310 => "0010110101011000",
30311 => "0010110101100000",
30312 => "0010110101100000",
30313 => "0010110101100000",
30314 => "0010110101100000",
30315 => "0010110101101000",
30316 => "0010110101101000",
30317 => "0010110101101000",
30318 => "0010110101101000",
30319 => "0010110101101000",
30320 => "0010110101110000",
30321 => "0010110101110000",
30322 => "0010110101110000",
30323 => "0010110101110000",
30324 => "0010110101111000",
30325 => "0010110101111000",
30326 => "0010110101111000",
30327 => "0010110101111000",
30328 => "0010110110000000",
30329 => "0010110110000000",
30330 => "0010110110000000",
30331 => "0010110110000000",
30332 => "0010110110000000",
30333 => "0010110110001000",
30334 => "0010110110001000",
30335 => "0010110110001000",
30336 => "0010110110001000",
30337 => "0010110110010000",
30338 => "0010110110010000",
30339 => "0010110110010000",
30340 => "0010110110010000",
30341 => "0010110110011000",
30342 => "0010110110011000",
30343 => "0010110110011000",
30344 => "0010110110011000",
30345 => "0010110110011000",
30346 => "0010110110100000",
30347 => "0010110110100000",
30348 => "0010110110100000",
30349 => "0010110110100000",
30350 => "0010110110101000",
30351 => "0010110110101000",
30352 => "0010110110101000",
30353 => "0010110110101000",
30354 => "0010110110101000",
30355 => "0010110110110000",
30356 => "0010110110110000",
30357 => "0010110110110000",
30358 => "0010110110110000",
30359 => "0010110110111000",
30360 => "0010110110111000",
30361 => "0010110110111000",
30362 => "0010110110111000",
30363 => "0010110111000000",
30364 => "0010110111000000",
30365 => "0010110111000000",
30366 => "0010110111000000",
30367 => "0010110111000000",
30368 => "0010110111001000",
30369 => "0010110111001000",
30370 => "0010110111001000",
30371 => "0010110111001000",
30372 => "0010110111010000",
30373 => "0010110111010000",
30374 => "0010110111010000",
30375 => "0010110111010000",
30376 => "0010110111011000",
30377 => "0010110111011000",
30378 => "0010110111011000",
30379 => "0010110111011000",
30380 => "0010110111011000",
30381 => "0010110111100000",
30382 => "0010110111100000",
30383 => "0010110111100000",
30384 => "0010110111100000",
30385 => "0010110111101000",
30386 => "0010110111101000",
30387 => "0010110111101000",
30388 => "0010110111101000",
30389 => "0010110111110000",
30390 => "0010110111110000",
30391 => "0010110111110000",
30392 => "0010110111110000",
30393 => "0010110111110000",
30394 => "0010110111111000",
30395 => "0010110111111000",
30396 => "0010110111111000",
30397 => "0010110111111000",
30398 => "0010111000000000",
30399 => "0010111000000000",
30400 => "0010111000000000",
30401 => "0010111000000000",
30402 => "0010111000001000",
30403 => "0010111000001000",
30404 => "0010111000001000",
30405 => "0010111000001000",
30406 => "0010111000001000",
30407 => "0010111000010000",
30408 => "0010111000010000",
30409 => "0010111000010000",
30410 => "0010111000010000",
30411 => "0010111000011000",
30412 => "0010111000011000",
30413 => "0010111000011000",
30414 => "0010111000011000",
30415 => "0010111000100000",
30416 => "0010111000100000",
30417 => "0010111000100000",
30418 => "0010111000100000",
30419 => "0010111000100000",
30420 => "0010111000101000",
30421 => "0010111000101000",
30422 => "0010111000101000",
30423 => "0010111000101000",
30424 => "0010111000110000",
30425 => "0010111000110000",
30426 => "0010111000110000",
30427 => "0010111000110000",
30428 => "0010111000111000",
30429 => "0010111000111000",
30430 => "0010111000111000",
30431 => "0010111000111000",
30432 => "0010111000111000",
30433 => "0010111001000000",
30434 => "0010111001000000",
30435 => "0010111001000000",
30436 => "0010111001000000",
30437 => "0010111001001000",
30438 => "0010111001001000",
30439 => "0010111001001000",
30440 => "0010111001001000",
30441 => "0010111001010000",
30442 => "0010111001010000",
30443 => "0010111001010000",
30444 => "0010111001010000",
30445 => "0010111001010000",
30446 => "0010111001011000",
30447 => "0010111001011000",
30448 => "0010111001011000",
30449 => "0010111001011000",
30450 => "0010111001100000",
30451 => "0010111001100000",
30452 => "0010111001100000",
30453 => "0010111001100000",
30454 => "0010111001101000",
30455 => "0010111001101000",
30456 => "0010111001101000",
30457 => "0010111001101000",
30458 => "0010111001101000",
30459 => "0010111001110000",
30460 => "0010111001110000",
30461 => "0010111001110000",
30462 => "0010111001110000",
30463 => "0010111001111000",
30464 => "0010111001111000",
30465 => "0010111001111000",
30466 => "0010111001111000",
30467 => "0010111010000000",
30468 => "0010111010000000",
30469 => "0010111010000000",
30470 => "0010111010000000",
30471 => "0010111010000000",
30472 => "0010111010001000",
30473 => "0010111010001000",
30474 => "0010111010001000",
30475 => "0010111010001000",
30476 => "0010111010010000",
30477 => "0010111010010000",
30478 => "0010111010010000",
30479 => "0010111010010000",
30480 => "0010111010011000",
30481 => "0010111010011000",
30482 => "0010111010011000",
30483 => "0010111010011000",
30484 => "0010111010011000",
30485 => "0010111010100000",
30486 => "0010111010100000",
30487 => "0010111010100000",
30488 => "0010111010100000",
30489 => "0010111010101000",
30490 => "0010111010101000",
30491 => "0010111010101000",
30492 => "0010111010101000",
30493 => "0010111010110000",
30494 => "0010111010110000",
30495 => "0010111010110000",
30496 => "0010111010110000",
30497 => "0010111010110000",
30498 => "0010111010111000",
30499 => "0010111010111000",
30500 => "0010111010111000",
30501 => "0010111010111000",
30502 => "0010111011000000",
30503 => "0010111011000000",
30504 => "0010111011000000",
30505 => "0010111011000000",
30506 => "0010111011001000",
30507 => "0010111011001000",
30508 => "0010111011001000",
30509 => "0010111011001000",
30510 => "0010111011001000",
30511 => "0010111011010000",
30512 => "0010111011010000",
30513 => "0010111011010000",
30514 => "0010111011010000",
30515 => "0010111011011000",
30516 => "0010111011011000",
30517 => "0010111011011000",
30518 => "0010111011011000",
30519 => "0010111011100000",
30520 => "0010111011100000",
30521 => "0010111011100000",
30522 => "0010111011100000",
30523 => "0010111011100000",
30524 => "0010111011101000",
30525 => "0010111011101000",
30526 => "0010111011101000",
30527 => "0010111011101000",
30528 => "0010111011110000",
30529 => "0010111011110000",
30530 => "0010111011110000",
30531 => "0010111011110000",
30532 => "0010111011111000",
30533 => "0010111011111000",
30534 => "0010111011111000",
30535 => "0010111011111000",
30536 => "0010111100000000",
30537 => "0010111100000000",
30538 => "0010111100000000",
30539 => "0010111100000000",
30540 => "0010111100000000",
30541 => "0010111100001000",
30542 => "0010111100001000",
30543 => "0010111100001000",
30544 => "0010111100001000",
30545 => "0010111100010000",
30546 => "0010111100010000",
30547 => "0010111100010000",
30548 => "0010111100010000",
30549 => "0010111100011000",
30550 => "0010111100011000",
30551 => "0010111100011000",
30552 => "0010111100011000",
30553 => "0010111100011000",
30554 => "0010111100100000",
30555 => "0010111100100000",
30556 => "0010111100100000",
30557 => "0010111100100000",
30558 => "0010111100101000",
30559 => "0010111100101000",
30560 => "0010111100101000",
30561 => "0010111100101000",
30562 => "0010111100110000",
30563 => "0010111100110000",
30564 => "0010111100110000",
30565 => "0010111100110000",
30566 => "0010111100110000",
30567 => "0010111100111000",
30568 => "0010111100111000",
30569 => "0010111100111000",
30570 => "0010111100111000",
30571 => "0010111101000000",
30572 => "0010111101000000",
30573 => "0010111101000000",
30574 => "0010111101000000",
30575 => "0010111101001000",
30576 => "0010111101001000",
30577 => "0010111101001000",
30578 => "0010111101001000",
30579 => "0010111101010000",
30580 => "0010111101010000",
30581 => "0010111101010000",
30582 => "0010111101010000",
30583 => "0010111101010000",
30584 => "0010111101011000",
30585 => "0010111101011000",
30586 => "0010111101011000",
30587 => "0010111101011000",
30588 => "0010111101100000",
30589 => "0010111101100000",
30590 => "0010111101100000",
30591 => "0010111101100000",
30592 => "0010111101101000",
30593 => "0010111101101000",
30594 => "0010111101101000",
30595 => "0010111101101000",
30596 => "0010111101101000",
30597 => "0010111101110000",
30598 => "0010111101110000",
30599 => "0010111101110000",
30600 => "0010111101110000",
30601 => "0010111101111000",
30602 => "0010111101111000",
30603 => "0010111101111000",
30604 => "0010111101111000",
30605 => "0010111110000000",
30606 => "0010111110000000",
30607 => "0010111110000000",
30608 => "0010111110000000",
30609 => "0010111110001000",
30610 => "0010111110001000",
30611 => "0010111110001000",
30612 => "0010111110001000",
30613 => "0010111110001000",
30614 => "0010111110010000",
30615 => "0010111110010000",
30616 => "0010111110010000",
30617 => "0010111110010000",
30618 => "0010111110011000",
30619 => "0010111110011000",
30620 => "0010111110011000",
30621 => "0010111110011000",
30622 => "0010111110100000",
30623 => "0010111110100000",
30624 => "0010111110100000",
30625 => "0010111110100000",
30626 => "0010111110100000",
30627 => "0010111110101000",
30628 => "0010111110101000",
30629 => "0010111110101000",
30630 => "0010111110101000",
30631 => "0010111110110000",
30632 => "0010111110110000",
30633 => "0010111110110000",
30634 => "0010111110110000",
30635 => "0010111110111000",
30636 => "0010111110111000",
30637 => "0010111110111000",
30638 => "0010111110111000",
30639 => "0010111111000000",
30640 => "0010111111000000",
30641 => "0010111111000000",
30642 => "0010111111000000",
30643 => "0010111111000000",
30644 => "0010111111001000",
30645 => "0010111111001000",
30646 => "0010111111001000",
30647 => "0010111111001000",
30648 => "0010111111010000",
30649 => "0010111111010000",
30650 => "0010111111010000",
30651 => "0010111111010000",
30652 => "0010111111011000",
30653 => "0010111111011000",
30654 => "0010111111011000",
30655 => "0010111111011000",
30656 => "0010111111100000",
30657 => "0010111111100000",
30658 => "0010111111100000",
30659 => "0010111111100000",
30660 => "0010111111100000",
30661 => "0010111111101000",
30662 => "0010111111101000",
30663 => "0010111111101000",
30664 => "0010111111101000",
30665 => "0010111111110000",
30666 => "0010111111110000",
30667 => "0010111111110000",
30668 => "0010111111110000",
30669 => "0010111111111000",
30670 => "0010111111111000",
30671 => "0010111111111000",
30672 => "0010111111111000",
30673 => "0010111111111000",
30674 => "0011000000000000",
30675 => "0011000000000000",
30676 => "0011000000000000",
30677 => "0011000000000000",
30678 => "0011000000001000",
30679 => "0011000000001000",
30680 => "0011000000001000",
30681 => "0011000000001000",
30682 => "0011000000010000",
30683 => "0011000000010000",
30684 => "0011000000010000",
30685 => "0011000000010000",
30686 => "0011000000011000",
30687 => "0011000000011000",
30688 => "0011000000011000",
30689 => "0011000000011000",
30690 => "0011000000011000",
30691 => "0011000000100000",
30692 => "0011000000100000",
30693 => "0011000000100000",
30694 => "0011000000100000",
30695 => "0011000000101000",
30696 => "0011000000101000",
30697 => "0011000000101000",
30698 => "0011000000101000",
30699 => "0011000000110000",
30700 => "0011000000110000",
30701 => "0011000000110000",
30702 => "0011000000110000",
30703 => "0011000000111000",
30704 => "0011000000111000",
30705 => "0011000000111000",
30706 => "0011000000111000",
30707 => "0011000000111000",
30708 => "0011000001000000",
30709 => "0011000001000000",
30710 => "0011000001000000",
30711 => "0011000001000000",
30712 => "0011000001001000",
30713 => "0011000001001000",
30714 => "0011000001001000",
30715 => "0011000001001000",
30716 => "0011000001010000",
30717 => "0011000001010000",
30718 => "0011000001010000",
30719 => "0011000001010000",
30720 => "0011000001011000",
30721 => "0011000001011000",
30722 => "0011000001011000",
30723 => "0011000001011000",
30724 => "0011000001011000",
30725 => "0011000001100000",
30726 => "0011000001100000",
30727 => "0011000001100000",
30728 => "0011000001100000",
30729 => "0011000001101000",
30730 => "0011000001101000",
30731 => "0011000001101000",
30732 => "0011000001101000",
30733 => "0011000001110000",
30734 => "0011000001110000",
30735 => "0011000001110000",
30736 => "0011000001110000",
30737 => "0011000001111000",
30738 => "0011000001111000",
30739 => "0011000001111000",
30740 => "0011000001111000",
30741 => "0011000001111000",
30742 => "0011000010000000",
30743 => "0011000010000000",
30744 => "0011000010000000",
30745 => "0011000010000000",
30746 => "0011000010001000",
30747 => "0011000010001000",
30748 => "0011000010001000",
30749 => "0011000010001000",
30750 => "0011000010010000",
30751 => "0011000010010000",
30752 => "0011000010010000",
30753 => "0011000010010000",
30754 => "0011000010011000",
30755 => "0011000010011000",
30756 => "0011000010011000",
30757 => "0011000010011000",
30758 => "0011000010011000",
30759 => "0011000010100000",
30760 => "0011000010100000",
30761 => "0011000010100000",
30762 => "0011000010100000",
30763 => "0011000010101000",
30764 => "0011000010101000",
30765 => "0011000010101000",
30766 => "0011000010101000",
30767 => "0011000010110000",
30768 => "0011000010110000",
30769 => "0011000010110000",
30770 => "0011000010110000",
30771 => "0011000010111000",
30772 => "0011000010111000",
30773 => "0011000010111000",
30774 => "0011000010111000",
30775 => "0011000010111000",
30776 => "0011000011000000",
30777 => "0011000011000000",
30778 => "0011000011000000",
30779 => "0011000011000000",
30780 => "0011000011001000",
30781 => "0011000011001000",
30782 => "0011000011001000",
30783 => "0011000011001000",
30784 => "0011000011010000",
30785 => "0011000011010000",
30786 => "0011000011010000",
30787 => "0011000011010000",
30788 => "0011000011011000",
30789 => "0011000011011000",
30790 => "0011000011011000",
30791 => "0011000011011000",
30792 => "0011000011011000",
30793 => "0011000011100000",
30794 => "0011000011100000",
30795 => "0011000011100000",
30796 => "0011000011100000",
30797 => "0011000011101000",
30798 => "0011000011101000",
30799 => "0011000011101000",
30800 => "0011000011101000",
30801 => "0011000011110000",
30802 => "0011000011110000",
30803 => "0011000011110000",
30804 => "0011000011110000",
30805 => "0011000011111000",
30806 => "0011000011111000",
30807 => "0011000011111000",
30808 => "0011000011111000",
30809 => "0011000011111000",
30810 => "0011000100000000",
30811 => "0011000100000000",
30812 => "0011000100000000",
30813 => "0011000100000000",
30814 => "0011000100001000",
30815 => "0011000100001000",
30816 => "0011000100001000",
30817 => "0011000100001000",
30818 => "0011000100010000",
30819 => "0011000100010000",
30820 => "0011000100010000",
30821 => "0011000100010000",
30822 => "0011000100011000",
30823 => "0011000100011000",
30824 => "0011000100011000",
30825 => "0011000100011000",
30826 => "0011000100100000",
30827 => "0011000100100000",
30828 => "0011000100100000",
30829 => "0011000100100000",
30830 => "0011000100100000",
30831 => "0011000100101000",
30832 => "0011000100101000",
30833 => "0011000100101000",
30834 => "0011000100101000",
30835 => "0011000100110000",
30836 => "0011000100110000",
30837 => "0011000100110000",
30838 => "0011000100110000",
30839 => "0011000100111000",
30840 => "0011000100111000",
30841 => "0011000100111000",
30842 => "0011000100111000",
30843 => "0011000101000000",
30844 => "0011000101000000",
30845 => "0011000101000000",
30846 => "0011000101000000",
30847 => "0011000101000000",
30848 => "0011000101001000",
30849 => "0011000101001000",
30850 => "0011000101001000",
30851 => "0011000101001000",
30852 => "0011000101010000",
30853 => "0011000101010000",
30854 => "0011000101010000",
30855 => "0011000101010000",
30856 => "0011000101011000",
30857 => "0011000101011000",
30858 => "0011000101011000",
30859 => "0011000101011000",
30860 => "0011000101100000",
30861 => "0011000101100000",
30862 => "0011000101100000",
30863 => "0011000101100000",
30864 => "0011000101101000",
30865 => "0011000101101000",
30866 => "0011000101101000",
30867 => "0011000101101000",
30868 => "0011000101101000",
30869 => "0011000101110000",
30870 => "0011000101110000",
30871 => "0011000101110000",
30872 => "0011000101110000",
30873 => "0011000101111000",
30874 => "0011000101111000",
30875 => "0011000101111000",
30876 => "0011000101111000",
30877 => "0011000110000000",
30878 => "0011000110000000",
30879 => "0011000110000000",
30880 => "0011000110000000",
30881 => "0011000110001000",
30882 => "0011000110001000",
30883 => "0011000110001000",
30884 => "0011000110001000",
30885 => "0011000110001000",
30886 => "0011000110010000",
30887 => "0011000110010000",
30888 => "0011000110010000",
30889 => "0011000110010000",
30890 => "0011000110011000",
30891 => "0011000110011000",
30892 => "0011000110011000",
30893 => "0011000110011000",
30894 => "0011000110100000",
30895 => "0011000110100000",
30896 => "0011000110100000",
30897 => "0011000110100000",
30898 => "0011000110101000",
30899 => "0011000110101000",
30900 => "0011000110101000",
30901 => "0011000110101000",
30902 => "0011000110110000",
30903 => "0011000110110000",
30904 => "0011000110110000",
30905 => "0011000110110000",
30906 => "0011000110110000",
30907 => "0011000110111000",
30908 => "0011000110111000",
30909 => "0011000110111000",
30910 => "0011000110111000",
30911 => "0011000111000000",
30912 => "0011000111000000",
30913 => "0011000111000000",
30914 => "0011000111000000",
30915 => "0011000111001000",
30916 => "0011000111001000",
30917 => "0011000111001000",
30918 => "0011000111001000",
30919 => "0011000111010000",
30920 => "0011000111010000",
30921 => "0011000111010000",
30922 => "0011000111010000",
30923 => "0011000111011000",
30924 => "0011000111011000",
30925 => "0011000111011000",
30926 => "0011000111011000",
30927 => "0011000111011000",
30928 => "0011000111100000",
30929 => "0011000111100000",
30930 => "0011000111100000",
30931 => "0011000111100000",
30932 => "0011000111101000",
30933 => "0011000111101000",
30934 => "0011000111101000",
30935 => "0011000111101000",
30936 => "0011000111110000",
30937 => "0011000111110000",
30938 => "0011000111110000",
30939 => "0011000111110000",
30940 => "0011000111111000",
30941 => "0011000111111000",
30942 => "0011000111111000",
30943 => "0011000111111000",
30944 => "0011001000000000",
30945 => "0011001000000000",
30946 => "0011001000000000",
30947 => "0011001000000000",
30948 => "0011001000000000",
30949 => "0011001000001000",
30950 => "0011001000001000",
30951 => "0011001000001000",
30952 => "0011001000001000",
30953 => "0011001000010000",
30954 => "0011001000010000",
30955 => "0011001000010000",
30956 => "0011001000010000",
30957 => "0011001000011000",
30958 => "0011001000011000",
30959 => "0011001000011000",
30960 => "0011001000011000",
30961 => "0011001000100000",
30962 => "0011001000100000",
30963 => "0011001000100000",
30964 => "0011001000100000",
30965 => "0011001000101000",
30966 => "0011001000101000",
30967 => "0011001000101000",
30968 => "0011001000101000",
30969 => "0011001000101000",
30970 => "0011001000110000",
30971 => "0011001000110000",
30972 => "0011001000110000",
30973 => "0011001000110000",
30974 => "0011001000111000",
30975 => "0011001000111000",
30976 => "0011001000111000",
30977 => "0011001000111000",
30978 => "0011001001000000",
30979 => "0011001001000000",
30980 => "0011001001000000",
30981 => "0011001001000000",
30982 => "0011001001001000",
30983 => "0011001001001000",
30984 => "0011001001001000",
30985 => "0011001001001000",
30986 => "0011001001010000",
30987 => "0011001001010000",
30988 => "0011001001010000",
30989 => "0011001001010000",
30990 => "0011001001010000",
30991 => "0011001001011000",
30992 => "0011001001011000",
30993 => "0011001001011000",
30994 => "0011001001011000",
30995 => "0011001001100000",
30996 => "0011001001100000",
30997 => "0011001001100000",
30998 => "0011001001100000",
30999 => "0011001001101000",
31000 => "0011001001101000",
31001 => "0011001001101000",
31002 => "0011001001101000",
31003 => "0011001001110000",
31004 => "0011001001110000",
31005 => "0011001001110000",
31006 => "0011001001110000",
31007 => "0011001001111000",
31008 => "0011001001111000",
31009 => "0011001001111000",
31010 => "0011001001111000",
31011 => "0011001001111000",
31012 => "0011001010000000",
31013 => "0011001010000000",
31014 => "0011001010000000",
31015 => "0011001010000000",
31016 => "0011001010001000",
31017 => "0011001010001000",
31018 => "0011001010001000",
31019 => "0011001010001000",
31020 => "0011001010010000",
31021 => "0011001010010000",
31022 => "0011001010010000",
31023 => "0011001010010000",
31024 => "0011001010011000",
31025 => "0011001010011000",
31026 => "0011001010011000",
31027 => "0011001010011000",
31028 => "0011001010100000",
31029 => "0011001010100000",
31030 => "0011001010100000",
31031 => "0011001010100000",
31032 => "0011001010100000",
31033 => "0011001010101000",
31034 => "0011001010101000",
31035 => "0011001010101000",
31036 => "0011001010101000",
31037 => "0011001010110000",
31038 => "0011001010110000",
31039 => "0011001010110000",
31040 => "0011001010110000",
31041 => "0011001010111000",
31042 => "0011001010111000",
31043 => "0011001010111000",
31044 => "0011001010111000",
31045 => "0011001011000000",
31046 => "0011001011000000",
31047 => "0011001011000000",
31048 => "0011001011000000",
31049 => "0011001011001000",
31050 => "0011001011001000",
31051 => "0011001011001000",
31052 => "0011001011001000",
31053 => "0011001011010000",
31054 => "0011001011010000",
31055 => "0011001011010000",
31056 => "0011001011010000",
31057 => "0011001011010000",
31058 => "0011001011011000",
31059 => "0011001011011000",
31060 => "0011001011011000",
31061 => "0011001011011000",
31062 => "0011001011100000",
31063 => "0011001011100000",
31064 => "0011001011100000",
31065 => "0011001011100000",
31066 => "0011001011101000",
31067 => "0011001011101000",
31068 => "0011001011101000",
31069 => "0011001011101000",
31070 => "0011001011110000",
31071 => "0011001011110000",
31072 => "0011001011110000",
31073 => "0011001011110000",
31074 => "0011001011111000",
31075 => "0011001011111000",
31076 => "0011001011111000",
31077 => "0011001011111000",
31078 => "0011001100000000",
31079 => "0011001100000000",
31080 => "0011001100000000",
31081 => "0011001100000000",
31082 => "0011001100000000",
31083 => "0011001100001000",
31084 => "0011001100001000",
31085 => "0011001100001000",
31086 => "0011001100001000",
31087 => "0011001100010000",
31088 => "0011001100010000",
31089 => "0011001100010000",
31090 => "0011001100010000",
31091 => "0011001100011000",
31092 => "0011001100011000",
31093 => "0011001100011000",
31094 => "0011001100011000",
31095 => "0011001100100000",
31096 => "0011001100100000",
31097 => "0011001100100000",
31098 => "0011001100100000",
31099 => "0011001100101000",
31100 => "0011001100101000",
31101 => "0011001100101000",
31102 => "0011001100101000",
31103 => "0011001100110000",
31104 => "0011001100110000",
31105 => "0011001100110000",
31106 => "0011001100110000",
31107 => "0011001100110000",
31108 => "0011001100111000",
31109 => "0011001100111000",
31110 => "0011001100111000",
31111 => "0011001100111000",
31112 => "0011001101000000",
31113 => "0011001101000000",
31114 => "0011001101000000",
31115 => "0011001101000000",
31116 => "0011001101001000",
31117 => "0011001101001000",
31118 => "0011001101001000",
31119 => "0011001101001000",
31120 => "0011001101010000",
31121 => "0011001101010000",
31122 => "0011001101010000",
31123 => "0011001101010000",
31124 => "0011001101011000",
31125 => "0011001101011000",
31126 => "0011001101011000",
31127 => "0011001101011000",
31128 => "0011001101100000",
31129 => "0011001101100000",
31130 => "0011001101100000",
31131 => "0011001101100000",
31132 => "0011001101100000",
31133 => "0011001101101000",
31134 => "0011001101101000",
31135 => "0011001101101000",
31136 => "0011001101101000",
31137 => "0011001101110000",
31138 => "0011001101110000",
31139 => "0011001101110000",
31140 => "0011001101110000",
31141 => "0011001101111000",
31142 => "0011001101111000",
31143 => "0011001101111000",
31144 => "0011001101111000",
31145 => "0011001110000000",
31146 => "0011001110000000",
31147 => "0011001110000000",
31148 => "0011001110000000",
31149 => "0011001110001000",
31150 => "0011001110001000",
31151 => "0011001110001000",
31152 => "0011001110001000",
31153 => "0011001110010000",
31154 => "0011001110010000",
31155 => "0011001110010000",
31156 => "0011001110010000",
31157 => "0011001110010000",
31158 => "0011001110011000",
31159 => "0011001110011000",
31160 => "0011001110011000",
31161 => "0011001110011000",
31162 => "0011001110100000",
31163 => "0011001110100000",
31164 => "0011001110100000",
31165 => "0011001110100000",
31166 => "0011001110101000",
31167 => "0011001110101000",
31168 => "0011001110101000",
31169 => "0011001110101000",
31170 => "0011001110110000",
31171 => "0011001110110000",
31172 => "0011001110110000",
31173 => "0011001110110000",
31174 => "0011001110111000",
31175 => "0011001110111000",
31176 => "0011001110111000",
31177 => "0011001110111000",
31178 => "0011001111000000",
31179 => "0011001111000000",
31180 => "0011001111000000",
31181 => "0011001111000000",
31182 => "0011001111000000",
31183 => "0011001111001000",
31184 => "0011001111001000",
31185 => "0011001111001000",
31186 => "0011001111001000",
31187 => "0011001111010000",
31188 => "0011001111010000",
31189 => "0011001111010000",
31190 => "0011001111010000",
31191 => "0011001111011000",
31192 => "0011001111011000",
31193 => "0011001111011000",
31194 => "0011001111011000",
31195 => "0011001111100000",
31196 => "0011001111100000",
31197 => "0011001111100000",
31198 => "0011001111100000",
31199 => "0011001111101000",
31200 => "0011001111101000",
31201 => "0011001111101000",
31202 => "0011001111101000",
31203 => "0011001111110000",
31204 => "0011001111110000",
31205 => "0011001111110000",
31206 => "0011001111110000",
31207 => "0011001111111000",
31208 => "0011001111111000",
31209 => "0011001111111000",
31210 => "0011001111111000",
31211 => "0011001111111000",
31212 => "0011010000000000",
31213 => "0011010000000000",
31214 => "0011010000000000",
31215 => "0011010000000000",
31216 => "0011010000001000",
31217 => "0011010000001000",
31218 => "0011010000001000",
31219 => "0011010000001000",
31220 => "0011010000010000",
31221 => "0011010000010000",
31222 => "0011010000010000",
31223 => "0011010000010000",
31224 => "0011010000011000",
31225 => "0011010000011000",
31226 => "0011010000011000",
31227 => "0011010000011000",
31228 => "0011010000100000",
31229 => "0011010000100000",
31230 => "0011010000100000",
31231 => "0011010000100000",
31232 => "0011010000101000",
31233 => "0011010000101000",
31234 => "0011010000101000",
31235 => "0011010000101000",
31236 => "0011010000110000",
31237 => "0011010000110000",
31238 => "0011010000110000",
31239 => "0011010000110000",
31240 => "0011010000110000",
31241 => "0011010000111000",
31242 => "0011010000111000",
31243 => "0011010000111000",
31244 => "0011010000111000",
31245 => "0011010001000000",
31246 => "0011010001000000",
31247 => "0011010001000000",
31248 => "0011010001000000",
31249 => "0011010001001000",
31250 => "0011010001001000",
31251 => "0011010001001000",
31252 => "0011010001001000",
31253 => "0011010001010000",
31254 => "0011010001010000",
31255 => "0011010001010000",
31256 => "0011010001010000",
31257 => "0011010001011000",
31258 => "0011010001011000",
31259 => "0011010001011000",
31260 => "0011010001011000",
31261 => "0011010001100000",
31262 => "0011010001100000",
31263 => "0011010001100000",
31264 => "0011010001100000",
31265 => "0011010001101000",
31266 => "0011010001101000",
31267 => "0011010001101000",
31268 => "0011010001101000",
31269 => "0011010001101000",
31270 => "0011010001110000",
31271 => "0011010001110000",
31272 => "0011010001110000",
31273 => "0011010001110000",
31274 => "0011010001111000",
31275 => "0011010001111000",
31276 => "0011010001111000",
31277 => "0011010001111000",
31278 => "0011010010000000",
31279 => "0011010010000000",
31280 => "0011010010000000",
31281 => "0011010010000000",
31282 => "0011010010001000",
31283 => "0011010010001000",
31284 => "0011010010001000",
31285 => "0011010010001000",
31286 => "0011010010010000",
31287 => "0011010010010000",
31288 => "0011010010010000",
31289 => "0011010010010000",
31290 => "0011010010011000",
31291 => "0011010010011000",
31292 => "0011010010011000",
31293 => "0011010010011000",
31294 => "0011010010100000",
31295 => "0011010010100000",
31296 => "0011010010100000",
31297 => "0011010010100000",
31298 => "0011010010101000",
31299 => "0011010010101000",
31300 => "0011010010101000",
31301 => "0011010010101000",
31302 => "0011010010101000",
31303 => "0011010010110000",
31304 => "0011010010110000",
31305 => "0011010010110000",
31306 => "0011010010110000",
31307 => "0011010010111000",
31308 => "0011010010111000",
31309 => "0011010010111000",
31310 => "0011010010111000",
31311 => "0011010011000000",
31312 => "0011010011000000",
31313 => "0011010011000000",
31314 => "0011010011000000",
31315 => "0011010011001000",
31316 => "0011010011001000",
31317 => "0011010011001000",
31318 => "0011010011001000",
31319 => "0011010011010000",
31320 => "0011010011010000",
31321 => "0011010011010000",
31322 => "0011010011010000",
31323 => "0011010011011000",
31324 => "0011010011011000",
31325 => "0011010011011000",
31326 => "0011010011011000",
31327 => "0011010011100000",
31328 => "0011010011100000",
31329 => "0011010011100000",
31330 => "0011010011100000",
31331 => "0011010011101000",
31332 => "0011010011101000",
31333 => "0011010011101000",
31334 => "0011010011101000",
31335 => "0011010011101000",
31336 => "0011010011110000",
31337 => "0011010011110000",
31338 => "0011010011110000",
31339 => "0011010011110000",
31340 => "0011010011111000",
31341 => "0011010011111000",
31342 => "0011010011111000",
31343 => "0011010011111000",
31344 => "0011010100000000",
31345 => "0011010100000000",
31346 => "0011010100000000",
31347 => "0011010100000000",
31348 => "0011010100001000",
31349 => "0011010100001000",
31350 => "0011010100001000",
31351 => "0011010100001000",
31352 => "0011010100010000",
31353 => "0011010100010000",
31354 => "0011010100010000",
31355 => "0011010100010000",
31356 => "0011010100011000",
31357 => "0011010100011000",
31358 => "0011010100011000",
31359 => "0011010100011000",
31360 => "0011010100100000",
31361 => "0011010100100000",
31362 => "0011010100100000",
31363 => "0011010100100000",
31364 => "0011010100101000",
31365 => "0011010100101000",
31366 => "0011010100101000",
31367 => "0011010100101000",
31368 => "0011010100101000",
31369 => "0011010100110000",
31370 => "0011010100110000",
31371 => "0011010100110000",
31372 => "0011010100110000",
31373 => "0011010100111000",
31374 => "0011010100111000",
31375 => "0011010100111000",
31376 => "0011010100111000",
31377 => "0011010101000000",
31378 => "0011010101000000",
31379 => "0011010101000000",
31380 => "0011010101000000",
31381 => "0011010101001000",
31382 => "0011010101001000",
31383 => "0011010101001000",
31384 => "0011010101001000",
31385 => "0011010101010000",
31386 => "0011010101010000",
31387 => "0011010101010000",
31388 => "0011010101010000",
31389 => "0011010101011000",
31390 => "0011010101011000",
31391 => "0011010101011000",
31392 => "0011010101011000",
31393 => "0011010101100000",
31394 => "0011010101100000",
31395 => "0011010101100000",
31396 => "0011010101100000",
31397 => "0011010101101000",
31398 => "0011010101101000",
31399 => "0011010101101000",
31400 => "0011010101101000",
31401 => "0011010101110000",
31402 => "0011010101110000",
31403 => "0011010101110000",
31404 => "0011010101110000",
31405 => "0011010101110000",
31406 => "0011010101111000",
31407 => "0011010101111000",
31408 => "0011010101111000",
31409 => "0011010101111000",
31410 => "0011010110000000",
31411 => "0011010110000000",
31412 => "0011010110000000",
31413 => "0011010110000000",
31414 => "0011010110001000",
31415 => "0011010110001000",
31416 => "0011010110001000",
31417 => "0011010110001000",
31418 => "0011010110010000",
31419 => "0011010110010000",
31420 => "0011010110010000",
31421 => "0011010110010000",
31422 => "0011010110011000",
31423 => "0011010110011000",
31424 => "0011010110011000",
31425 => "0011010110011000",
31426 => "0011010110100000",
31427 => "0011010110100000",
31428 => "0011010110100000",
31429 => "0011010110100000",
31430 => "0011010110101000",
31431 => "0011010110101000",
31432 => "0011010110101000",
31433 => "0011010110101000",
31434 => "0011010110110000",
31435 => "0011010110110000",
31436 => "0011010110110000",
31437 => "0011010110110000",
31438 => "0011010110111000",
31439 => "0011010110111000",
31440 => "0011010110111000",
31441 => "0011010110111000",
31442 => "0011010110111000",
31443 => "0011010111000000",
31444 => "0011010111000000",
31445 => "0011010111000000",
31446 => "0011010111000000",
31447 => "0011010111001000",
31448 => "0011010111001000",
31449 => "0011010111001000",
31450 => "0011010111001000",
31451 => "0011010111010000",
31452 => "0011010111010000",
31453 => "0011010111010000",
31454 => "0011010111010000",
31455 => "0011010111011000",
31456 => "0011010111011000",
31457 => "0011010111011000",
31458 => "0011010111011000",
31459 => "0011010111100000",
31460 => "0011010111100000",
31461 => "0011010111100000",
31462 => "0011010111100000",
31463 => "0011010111101000",
31464 => "0011010111101000",
31465 => "0011010111101000",
31466 => "0011010111101000",
31467 => "0011010111110000",
31468 => "0011010111110000",
31469 => "0011010111110000",
31470 => "0011010111110000",
31471 => "0011010111111000",
31472 => "0011010111111000",
31473 => "0011010111111000",
31474 => "0011010111111000",
31475 => "0011011000000000",
31476 => "0011011000000000",
31477 => "0011011000000000",
31478 => "0011011000000000",
31479 => "0011011000001000",
31480 => "0011011000001000",
31481 => "0011011000001000",
31482 => "0011011000001000",
31483 => "0011011000001000",
31484 => "0011011000010000",
31485 => "0011011000010000",
31486 => "0011011000010000",
31487 => "0011011000010000",
31488 => "0011011000011000",
31489 => "0011011000011000",
31490 => "0011011000011000",
31491 => "0011011000011000",
31492 => "0011011000100000",
31493 => "0011011000100000",
31494 => "0011011000100000",
31495 => "0011011000100000",
31496 => "0011011000101000",
31497 => "0011011000101000",
31498 => "0011011000101000",
31499 => "0011011000101000",
31500 => "0011011000110000",
31501 => "0011011000110000",
31502 => "0011011000110000",
31503 => "0011011000110000",
31504 => "0011011000111000",
31505 => "0011011000111000",
31506 => "0011011000111000",
31507 => "0011011000111000",
31508 => "0011011001000000",
31509 => "0011011001000000",
31510 => "0011011001000000",
31511 => "0011011001000000",
31512 => "0011011001001000",
31513 => "0011011001001000",
31514 => "0011011001001000",
31515 => "0011011001001000",
31516 => "0011011001010000",
31517 => "0011011001010000",
31518 => "0011011001010000",
31519 => "0011011001010000",
31520 => "0011011001011000",
31521 => "0011011001011000",
31522 => "0011011001011000",
31523 => "0011011001011000",
31524 => "0011011001011000",
31525 => "0011011001100000",
31526 => "0011011001100000",
31527 => "0011011001100000",
31528 => "0011011001100000",
31529 => "0011011001101000",
31530 => "0011011001101000",
31531 => "0011011001101000",
31532 => "0011011001101000",
31533 => "0011011001110000",
31534 => "0011011001110000",
31535 => "0011011001110000",
31536 => "0011011001110000",
31537 => "0011011001111000",
31538 => "0011011001111000",
31539 => "0011011001111000",
31540 => "0011011001111000",
31541 => "0011011010000000",
31542 => "0011011010000000",
31543 => "0011011010000000",
31544 => "0011011010000000",
31545 => "0011011010001000",
31546 => "0011011010001000",
31547 => "0011011010001000",
31548 => "0011011010001000",
31549 => "0011011010010000",
31550 => "0011011010010000",
31551 => "0011011010010000",
31552 => "0011011010010000",
31553 => "0011011010011000",
31554 => "0011011010011000",
31555 => "0011011010011000",
31556 => "0011011010011000",
31557 => "0011011010100000",
31558 => "0011011010100000",
31559 => "0011011010100000",
31560 => "0011011010100000",
31561 => "0011011010101000",
31562 => "0011011010101000",
31563 => "0011011010101000",
31564 => "0011011010101000",
31565 => "0011011010110000",
31566 => "0011011010110000",
31567 => "0011011010110000",
31568 => "0011011010110000",
31569 => "0011011010110000",
31570 => "0011011010111000",
31571 => "0011011010111000",
31572 => "0011011010111000",
31573 => "0011011010111000",
31574 => "0011011011000000",
31575 => "0011011011000000",
31576 => "0011011011000000",
31577 => "0011011011000000",
31578 => "0011011011001000",
31579 => "0011011011001000",
31580 => "0011011011001000",
31581 => "0011011011001000",
31582 => "0011011011010000",
31583 => "0011011011010000",
31584 => "0011011011010000",
31585 => "0011011011010000",
31586 => "0011011011011000",
31587 => "0011011011011000",
31588 => "0011011011011000",
31589 => "0011011011011000",
31590 => "0011011011100000",
31591 => "0011011011100000",
31592 => "0011011011100000",
31593 => "0011011011100000",
31594 => "0011011011101000",
31595 => "0011011011101000",
31596 => "0011011011101000",
31597 => "0011011011101000",
31598 => "0011011011110000",
31599 => "0011011011110000",
31600 => "0011011011110000",
31601 => "0011011011110000",
31602 => "0011011011111000",
31603 => "0011011011111000",
31604 => "0011011011111000",
31605 => "0011011011111000",
31606 => "0011011100000000",
31607 => "0011011100000000",
31608 => "0011011100000000",
31609 => "0011011100000000",
31610 => "0011011100001000",
31611 => "0011011100001000",
31612 => "0011011100001000",
31613 => "0011011100001000",
31614 => "0011011100010000",
31615 => "0011011100010000",
31616 => "0011011100010000",
31617 => "0011011100010000",
31618 => "0011011100010000",
31619 => "0011011100011000",
31620 => "0011011100011000",
31621 => "0011011100011000",
31622 => "0011011100011000",
31623 => "0011011100100000",
31624 => "0011011100100000",
31625 => "0011011100100000",
31626 => "0011011100100000",
31627 => "0011011100101000",
31628 => "0011011100101000",
31629 => "0011011100101000",
31630 => "0011011100101000",
31631 => "0011011100110000",
31632 => "0011011100110000",
31633 => "0011011100110000",
31634 => "0011011100110000",
31635 => "0011011100111000",
31636 => "0011011100111000",
31637 => "0011011100111000",
31638 => "0011011100111000",
31639 => "0011011101000000",
31640 => "0011011101000000",
31641 => "0011011101000000",
31642 => "0011011101000000",
31643 => "0011011101001000",
31644 => "0011011101001000",
31645 => "0011011101001000",
31646 => "0011011101001000",
31647 => "0011011101010000",
31648 => "0011011101010000",
31649 => "0011011101010000",
31650 => "0011011101010000",
31651 => "0011011101011000",
31652 => "0011011101011000",
31653 => "0011011101011000",
31654 => "0011011101011000",
31655 => "0011011101100000",
31656 => "0011011101100000",
31657 => "0011011101100000",
31658 => "0011011101100000",
31659 => "0011011101101000",
31660 => "0011011101101000",
31661 => "0011011101101000",
31662 => "0011011101101000",
31663 => "0011011101110000",
31664 => "0011011101110000",
31665 => "0011011101110000",
31666 => "0011011101110000",
31667 => "0011011101111000",
31668 => "0011011101111000",
31669 => "0011011101111000",
31670 => "0011011101111000",
31671 => "0011011101111000",
31672 => "0011011110000000",
31673 => "0011011110000000",
31674 => "0011011110000000",
31675 => "0011011110000000",
31676 => "0011011110001000",
31677 => "0011011110001000",
31678 => "0011011110001000",
31679 => "0011011110001000",
31680 => "0011011110010000",
31681 => "0011011110010000",
31682 => "0011011110010000",
31683 => "0011011110010000",
31684 => "0011011110011000",
31685 => "0011011110011000",
31686 => "0011011110011000",
31687 => "0011011110011000",
31688 => "0011011110100000",
31689 => "0011011110100000",
31690 => "0011011110100000",
31691 => "0011011110100000",
31692 => "0011011110101000",
31693 => "0011011110101000",
31694 => "0011011110101000",
31695 => "0011011110101000",
31696 => "0011011110110000",
31697 => "0011011110110000",
31698 => "0011011110110000",
31699 => "0011011110110000",
31700 => "0011011110111000",
31701 => "0011011110111000",
31702 => "0011011110111000",
31703 => "0011011110111000",
31704 => "0011011111000000",
31705 => "0011011111000000",
31706 => "0011011111000000",
31707 => "0011011111000000",
31708 => "0011011111001000",
31709 => "0011011111001000",
31710 => "0011011111001000",
31711 => "0011011111001000",
31712 => "0011011111010000",
31713 => "0011011111010000",
31714 => "0011011111010000",
31715 => "0011011111010000",
31716 => "0011011111011000",
31717 => "0011011111011000",
31718 => "0011011111011000",
31719 => "0011011111011000",
31720 => "0011011111100000",
31721 => "0011011111100000",
31722 => "0011011111100000",
31723 => "0011011111100000",
31724 => "0011011111101000",
31725 => "0011011111101000",
31726 => "0011011111101000",
31727 => "0011011111101000",
31728 => "0011011111110000",
31729 => "0011011111110000",
31730 => "0011011111110000",
31731 => "0011011111110000",
31732 => "0011011111110000",
31733 => "0011011111111000",
31734 => "0011011111111000",
31735 => "0011011111111000",
31736 => "0011011111111000",
31737 => "0011100000000000",
31738 => "0011100000000000",
31739 => "0011100000000000",
31740 => "0011100000000000",
31741 => "0011100000001000",
31742 => "0011100000001000",
31743 => "0011100000001000",
31744 => "0011100000001000",
31745 => "0011100000010000",
31746 => "0011100000010000",
31747 => "0011100000010000",
31748 => "0011100000010000",
31749 => "0011100000011000",
31750 => "0011100000011000",
31751 => "0011100000011000",
31752 => "0011100000011000",
31753 => "0011100000100000",
31754 => "0011100000100000",
31755 => "0011100000100000",
31756 => "0011100000100000",
31757 => "0011100000101000",
31758 => "0011100000101000",
31759 => "0011100000101000",
31760 => "0011100000101000",
31761 => "0011100000110000",
31762 => "0011100000110000",
31763 => "0011100000110000",
31764 => "0011100000110000",
31765 => "0011100000111000",
31766 => "0011100000111000",
31767 => "0011100000111000",
31768 => "0011100000111000",
31769 => "0011100001000000",
31770 => "0011100001000000",
31771 => "0011100001000000",
31772 => "0011100001000000",
31773 => "0011100001001000",
31774 => "0011100001001000",
31775 => "0011100001001000",
31776 => "0011100001001000",
31777 => "0011100001010000",
31778 => "0011100001010000",
31779 => "0011100001010000",
31780 => "0011100001010000",
31781 => "0011100001011000",
31782 => "0011100001011000",
31783 => "0011100001011000",
31784 => "0011100001011000",
31785 => "0011100001100000",
31786 => "0011100001100000",
31787 => "0011100001100000",
31788 => "0011100001100000",
31789 => "0011100001101000",
31790 => "0011100001101000",
31791 => "0011100001101000",
31792 => "0011100001101000",
31793 => "0011100001110000",
31794 => "0011100001110000",
31795 => "0011100001110000",
31796 => "0011100001110000",
31797 => "0011100001111000",
31798 => "0011100001111000",
31799 => "0011100001111000",
31800 => "0011100001111000",
31801 => "0011100001111000",
31802 => "0011100010000000",
31803 => "0011100010000000",
31804 => "0011100010000000",
31805 => "0011100010000000",
31806 => "0011100010001000",
31807 => "0011100010001000",
31808 => "0011100010001000",
31809 => "0011100010001000",
31810 => "0011100010010000",
31811 => "0011100010010000",
31812 => "0011100010010000",
31813 => "0011100010010000",
31814 => "0011100010011000",
31815 => "0011100010011000",
31816 => "0011100010011000",
31817 => "0011100010011000",
31818 => "0011100010100000",
31819 => "0011100010100000",
31820 => "0011100010100000",
31821 => "0011100010100000",
31822 => "0011100010101000",
31823 => "0011100010101000",
31824 => "0011100010101000",
31825 => "0011100010101000",
31826 => "0011100010110000",
31827 => "0011100010110000",
31828 => "0011100010110000",
31829 => "0011100010110000",
31830 => "0011100010111000",
31831 => "0011100010111000",
31832 => "0011100010111000",
31833 => "0011100010111000",
31834 => "0011100011000000",
31835 => "0011100011000000",
31836 => "0011100011000000",
31837 => "0011100011000000",
31838 => "0011100011001000",
31839 => "0011100011001000",
31840 => "0011100011001000",
31841 => "0011100011001000",
31842 => "0011100011010000",
31843 => "0011100011010000",
31844 => "0011100011010000",
31845 => "0011100011010000",
31846 => "0011100011011000",
31847 => "0011100011011000",
31848 => "0011100011011000",
31849 => "0011100011011000",
31850 => "0011100011100000",
31851 => "0011100011100000",
31852 => "0011100011100000",
31853 => "0011100011100000",
31854 => "0011100011101000",
31855 => "0011100011101000",
31856 => "0011100011101000",
31857 => "0011100011101000",
31858 => "0011100011110000",
31859 => "0011100011110000",
31860 => "0011100011110000",
31861 => "0011100011110000",
31862 => "0011100011111000",
31863 => "0011100011111000",
31864 => "0011100011111000",
31865 => "0011100011111000",
31866 => "0011100100000000",
31867 => "0011100100000000",
31868 => "0011100100000000",
31869 => "0011100100000000",
31870 => "0011100100001000",
31871 => "0011100100001000",
31872 => "0011100100001000",
31873 => "0011100100001000",
31874 => "0011100100010000",
31875 => "0011100100010000",
31876 => "0011100100010000",
31877 => "0011100100010000",
31878 => "0011100100010000",
31879 => "0011100100011000",
31880 => "0011100100011000",
31881 => "0011100100011000",
31882 => "0011100100011000",
31883 => "0011100100100000",
31884 => "0011100100100000",
31885 => "0011100100100000",
31886 => "0011100100100000",
31887 => "0011100100101000",
31888 => "0011100100101000",
31889 => "0011100100101000",
31890 => "0011100100101000",
31891 => "0011100100110000",
31892 => "0011100100110000",
31893 => "0011100100110000",
31894 => "0011100100110000",
31895 => "0011100100111000",
31896 => "0011100100111000",
31897 => "0011100100111000",
31898 => "0011100100111000",
31899 => "0011100101000000",
31900 => "0011100101000000",
31901 => "0011100101000000",
31902 => "0011100101000000",
31903 => "0011100101001000",
31904 => "0011100101001000",
31905 => "0011100101001000",
31906 => "0011100101001000",
31907 => "0011100101010000",
31908 => "0011100101010000",
31909 => "0011100101010000",
31910 => "0011100101010000",
31911 => "0011100101011000",
31912 => "0011100101011000",
31913 => "0011100101011000",
31914 => "0011100101011000",
31915 => "0011100101100000",
31916 => "0011100101100000",
31917 => "0011100101100000",
31918 => "0011100101100000",
31919 => "0011100101101000",
31920 => "0011100101101000",
31921 => "0011100101101000",
31922 => "0011100101101000",
31923 => "0011100101110000",
31924 => "0011100101110000",
31925 => "0011100101110000",
31926 => "0011100101110000",
31927 => "0011100101111000",
31928 => "0011100101111000",
31929 => "0011100101111000",
31930 => "0011100101111000",
31931 => "0011100110000000",
31932 => "0011100110000000",
31933 => "0011100110000000",
31934 => "0011100110000000",
31935 => "0011100110001000",
31936 => "0011100110001000",
31937 => "0011100110001000",
31938 => "0011100110001000",
31939 => "0011100110010000",
31940 => "0011100110010000",
31941 => "0011100110010000",
31942 => "0011100110010000",
31943 => "0011100110011000",
31944 => "0011100110011000",
31945 => "0011100110011000",
31946 => "0011100110011000",
31947 => "0011100110100000",
31948 => "0011100110100000",
31949 => "0011100110100000",
31950 => "0011100110100000",
31951 => "0011100110101000",
31952 => "0011100110101000",
31953 => "0011100110101000",
31954 => "0011100110101000",
31955 => "0011100110110000",
31956 => "0011100110110000",
31957 => "0011100110110000",
31958 => "0011100110110000",
31959 => "0011100110111000",
31960 => "0011100110111000",
31961 => "0011100110111000",
31962 => "0011100110111000",
31963 => "0011100111000000",
31964 => "0011100111000000",
31965 => "0011100111000000",
31966 => "0011100111000000",
31967 => "0011100111001000",
31968 => "0011100111001000",
31969 => "0011100111001000",
31970 => "0011100111001000",
31971 => "0011100111001000",
31972 => "0011100111010000",
31973 => "0011100111010000",
31974 => "0011100111010000",
31975 => "0011100111010000",
31976 => "0011100111011000",
31977 => "0011100111011000",
31978 => "0011100111011000",
31979 => "0011100111011000",
31980 => "0011100111100000",
31981 => "0011100111100000",
31982 => "0011100111100000",
31983 => "0011100111100000",
31984 => "0011100111101000",
31985 => "0011100111101000",
31986 => "0011100111101000",
31987 => "0011100111101000",
31988 => "0011100111110000",
31989 => "0011100111110000",
31990 => "0011100111110000",
31991 => "0011100111110000",
31992 => "0011100111111000",
31993 => "0011100111111000",
31994 => "0011100111111000",
31995 => "0011100111111000",
31996 => "0011101000000000",
31997 => "0011101000000000",
31998 => "0011101000000000",
31999 => "0011101000000000",
32000 => "0011101000001000",
32001 => "0011101000001000",
32002 => "0011101000001000",
32003 => "0011101000001000",
32004 => "0011101000010000",
32005 => "0011101000010000",
32006 => "0011101000010000",
32007 => "0011101000010000",
32008 => "0011101000011000",
32009 => "0011101000011000",
32010 => "0011101000011000",
32011 => "0011101000011000",
32012 => "0011101000100000",
32013 => "0011101000100000",
32014 => "0011101000100000",
32015 => "0011101000100000",
32016 => "0011101000101000",
32017 => "0011101000101000",
32018 => "0011101000101000",
32019 => "0011101000101000",
32020 => "0011101000110000",
32021 => "0011101000110000",
32022 => "0011101000110000",
32023 => "0011101000110000",
32024 => "0011101000111000",
32025 => "0011101000111000",
32026 => "0011101000111000",
32027 => "0011101000111000",
32028 => "0011101001000000",
32029 => "0011101001000000",
32030 => "0011101001000000",
32031 => "0011101001000000",
32032 => "0011101001001000",
32033 => "0011101001001000",
32034 => "0011101001001000",
32035 => "0011101001001000",
32036 => "0011101001010000",
32037 => "0011101001010000",
32038 => "0011101001010000",
32039 => "0011101001010000",
32040 => "0011101001011000",
32041 => "0011101001011000",
32042 => "0011101001011000",
32043 => "0011101001011000",
32044 => "0011101001100000",
32045 => "0011101001100000",
32046 => "0011101001100000",
32047 => "0011101001100000",
32048 => "0011101001101000",
32049 => "0011101001101000",
32050 => "0011101001101000",
32051 => "0011101001101000",
32052 => "0011101001110000",
32053 => "0011101001110000",
32054 => "0011101001110000",
32055 => "0011101001110000",
32056 => "0011101001111000",
32057 => "0011101001111000",
32058 => "0011101001111000",
32059 => "0011101001111000",
32060 => "0011101010000000",
32061 => "0011101010000000",
32062 => "0011101010000000",
32063 => "0011101010000000",
32064 => "0011101010001000",
32065 => "0011101010001000",
32066 => "0011101010001000",
32067 => "0011101010001000",
32068 => "0011101010010000",
32069 => "0011101010010000",
32070 => "0011101010010000",
32071 => "0011101010010000",
32072 => "0011101010011000",
32073 => "0011101010011000",
32074 => "0011101010011000",
32075 => "0011101010011000",
32076 => "0011101010100000",
32077 => "0011101010100000",
32078 => "0011101010100000",
32079 => "0011101010100000",
32080 => "0011101010101000",
32081 => "0011101010101000",
32082 => "0011101010101000",
32083 => "0011101010101000",
32084 => "0011101010110000",
32085 => "0011101010110000",
32086 => "0011101010110000",
32087 => "0011101010110000",
32088 => "0011101010111000",
32089 => "0011101010111000",
32090 => "0011101010111000",
32091 => "0011101010111000",
32092 => "0011101011000000",
32093 => "0011101011000000",
32094 => "0011101011000000",
32095 => "0011101011000000",
32096 => "0011101011000000",
32097 => "0011101011001000",
32098 => "0011101011001000",
32099 => "0011101011001000",
32100 => "0011101011001000",
32101 => "0011101011010000",
32102 => "0011101011010000",
32103 => "0011101011010000",
32104 => "0011101011010000",
32105 => "0011101011011000",
32106 => "0011101011011000",
32107 => "0011101011011000",
32108 => "0011101011011000",
32109 => "0011101011100000",
32110 => "0011101011100000",
32111 => "0011101011100000",
32112 => "0011101011100000",
32113 => "0011101011101000",
32114 => "0011101011101000",
32115 => "0011101011101000",
32116 => "0011101011101000",
32117 => "0011101011110000",
32118 => "0011101011110000",
32119 => "0011101011110000",
32120 => "0011101011110000",
32121 => "0011101011111000",
32122 => "0011101011111000",
32123 => "0011101011111000",
32124 => "0011101011111000",
32125 => "0011101100000000",
32126 => "0011101100000000",
32127 => "0011101100000000",
32128 => "0011101100000000",
32129 => "0011101100001000",
32130 => "0011101100001000",
32131 => "0011101100001000",
32132 => "0011101100001000",
32133 => "0011101100010000",
32134 => "0011101100010000",
32135 => "0011101100010000",
32136 => "0011101100010000",
32137 => "0011101100011000",
32138 => "0011101100011000",
32139 => "0011101100011000",
32140 => "0011101100011000",
32141 => "0011101100100000",
32142 => "0011101100100000",
32143 => "0011101100100000",
32144 => "0011101100100000",
32145 => "0011101100101000",
32146 => "0011101100101000",
32147 => "0011101100101000",
32148 => "0011101100101000",
32149 => "0011101100110000",
32150 => "0011101100110000",
32151 => "0011101100110000",
32152 => "0011101100110000",
32153 => "0011101100111000",
32154 => "0011101100111000",
32155 => "0011101100111000",
32156 => "0011101100111000",
32157 => "0011101101000000",
32158 => "0011101101000000",
32159 => "0011101101000000",
32160 => "0011101101000000",
32161 => "0011101101001000",
32162 => "0011101101001000",
32163 => "0011101101001000",
32164 => "0011101101001000",
32165 => "0011101101010000",
32166 => "0011101101010000",
32167 => "0011101101010000",
32168 => "0011101101010000",
32169 => "0011101101011000",
32170 => "0011101101011000",
32171 => "0011101101011000",
32172 => "0011101101011000",
32173 => "0011101101100000",
32174 => "0011101101100000",
32175 => "0011101101100000",
32176 => "0011101101100000",
32177 => "0011101101101000",
32178 => "0011101101101000",
32179 => "0011101101101000",
32180 => "0011101101101000",
32181 => "0011101101110000",
32182 => "0011101101110000",
32183 => "0011101101110000",
32184 => "0011101101110000",
32185 => "0011101101111000",
32186 => "0011101101111000",
32187 => "0011101101111000",
32188 => "0011101101111000",
32189 => "0011101110000000",
32190 => "0011101110000000",
32191 => "0011101110000000",
32192 => "0011101110000000",
32193 => "0011101110001000",
32194 => "0011101110001000",
32195 => "0011101110001000",
32196 => "0011101110001000",
32197 => "0011101110010000",
32198 => "0011101110010000",
32199 => "0011101110010000",
32200 => "0011101110010000",
32201 => "0011101110011000",
32202 => "0011101110011000",
32203 => "0011101110011000",
32204 => "0011101110011000",
32205 => "0011101110100000",
32206 => "0011101110100000",
32207 => "0011101110100000",
32208 => "0011101110100000",
32209 => "0011101110101000",
32210 => "0011101110101000",
32211 => "0011101110101000",
32212 => "0011101110101000",
32213 => "0011101110110000",
32214 => "0011101110110000",
32215 => "0011101110110000",
32216 => "0011101110110000",
32217 => "0011101110111000",
32218 => "0011101110111000",
32219 => "0011101110111000",
32220 => "0011101110111000",
32221 => "0011101111000000",
32222 => "0011101111000000",
32223 => "0011101111000000",
32224 => "0011101111000000",
32225 => "0011101111001000",
32226 => "0011101111001000",
32227 => "0011101111001000",
32228 => "0011101111001000",
32229 => "0011101111010000",
32230 => "0011101111010000",
32231 => "0011101111010000",
32232 => "0011101111010000",
32233 => "0011101111011000",
32234 => "0011101111011000",
32235 => "0011101111011000",
32236 => "0011101111011000",
32237 => "0011101111100000",
32238 => "0011101111100000",
32239 => "0011101111100000",
32240 => "0011101111100000",
32241 => "0011101111101000",
32242 => "0011101111101000",
32243 => "0011101111101000",
32244 => "0011101111101000",
32245 => "0011101111110000",
32246 => "0011101111110000",
32247 => "0011101111110000",
32248 => "0011101111110000",
32249 => "0011101111111000",
32250 => "0011101111111000",
32251 => "0011101111111000",
32252 => "0011101111111000",
32253 => "0011110000000000",
32254 => "0011110000000000",
32255 => "0011110000000000",
32256 => "0011110000000000",
32257 => "0011110000001000",
32258 => "0011110000001000",
32259 => "0011110000001000",
32260 => "0011110000001000",
32261 => "0011110000010000",
32262 => "0011110000010000",
32263 => "0011110000010000",
32264 => "0011110000010000",
32265 => "0011110000011000",
32266 => "0011110000011000",
32267 => "0011110000011000",
32268 => "0011110000011000",
32269 => "0011110000100000",
32270 => "0011110000100000",
32271 => "0011110000100000",
32272 => "0011110000100000",
32273 => "0011110000101000",
32274 => "0011110000101000",
32275 => "0011110000101000",
32276 => "0011110000101000",
32277 => "0011110000110000",
32278 => "0011110000110000",
32279 => "0011110000110000",
32280 => "0011110000110000",
32281 => "0011110000111000",
32282 => "0011110000111000",
32283 => "0011110000111000",
32284 => "0011110000111000",
32285 => "0011110001000000",
32286 => "0011110001000000",
32287 => "0011110001000000",
32288 => "0011110001000000",
32289 => "0011110001001000",
32290 => "0011110001001000",
32291 => "0011110001001000",
32292 => "0011110001001000",
32293 => "0011110001010000",
32294 => "0011110001010000",
32295 => "0011110001010000",
32296 => "0011110001010000",
32297 => "0011110001011000",
32298 => "0011110001011000",
32299 => "0011110001011000",
32300 => "0011110001011000",
32301 => "0011110001011000",
32302 => "0011110001100000",
32303 => "0011110001100000",
32304 => "0011110001100000",
32305 => "0011110001100000",
32306 => "0011110001101000",
32307 => "0011110001101000",
32308 => "0011110001101000",
32309 => "0011110001101000",
32310 => "0011110001110000",
32311 => "0011110001110000",
32312 => "0011110001110000",
32313 => "0011110001110000",
32314 => "0011110001111000",
32315 => "0011110001111000",
32316 => "0011110001111000",
32317 => "0011110001111000",
32318 => "0011110010000000",
32319 => "0011110010000000",
32320 => "0011110010000000",
32321 => "0011110010000000",
32322 => "0011110010001000",
32323 => "0011110010001000",
32324 => "0011110010001000",
32325 => "0011110010001000",
32326 => "0011110010010000",
32327 => "0011110010010000",
32328 => "0011110010010000",
32329 => "0011110010010000",
32330 => "0011110010011000",
32331 => "0011110010011000",
32332 => "0011110010011000",
32333 => "0011110010011000",
32334 => "0011110010100000",
32335 => "0011110010100000",
32336 => "0011110010100000",
32337 => "0011110010100000",
32338 => "0011110010101000",
32339 => "0011110010101000",
32340 => "0011110010101000",
32341 => "0011110010101000",
32342 => "0011110010110000",
32343 => "0011110010110000",
32344 => "0011110010110000",
32345 => "0011110010110000",
32346 => "0011110010111000",
32347 => "0011110010111000",
32348 => "0011110010111000",
32349 => "0011110010111000",
32350 => "0011110011000000",
32351 => "0011110011000000",
32352 => "0011110011000000",
32353 => "0011110011000000",
32354 => "0011110011001000",
32355 => "0011110011001000",
32356 => "0011110011001000",
32357 => "0011110011001000",
32358 => "0011110011010000",
32359 => "0011110011010000",
32360 => "0011110011010000",
32361 => "0011110011010000",
32362 => "0011110011011000",
32363 => "0011110011011000",
32364 => "0011110011011000",
32365 => "0011110011011000",
32366 => "0011110011100000",
32367 => "0011110011100000",
32368 => "0011110011100000",
32369 => "0011110011100000",
32370 => "0011110011101000",
32371 => "0011110011101000",
32372 => "0011110011101000",
32373 => "0011110011101000",
32374 => "0011110011110000",
32375 => "0011110011110000",
32376 => "0011110011110000",
32377 => "0011110011110000",
32378 => "0011110011111000",
32379 => "0011110011111000",
32380 => "0011110011111000",
32381 => "0011110011111000",
32382 => "0011110100000000",
32383 => "0011110100000000",
32384 => "0011110100000000",
32385 => "0011110100000000",
32386 => "0011110100001000",
32387 => "0011110100001000",
32388 => "0011110100001000",
32389 => "0011110100001000",
32390 => "0011110100010000",
32391 => "0011110100010000",
32392 => "0011110100010000",
32393 => "0011110100010000",
32394 => "0011110100011000",
32395 => "0011110100011000",
32396 => "0011110100011000",
32397 => "0011110100011000",
32398 => "0011110100100000",
32399 => "0011110100100000",
32400 => "0011110100100000",
32401 => "0011110100100000",
32402 => "0011110100101000",
32403 => "0011110100101000",
32404 => "0011110100101000",
32405 => "0011110100101000",
32406 => "0011110100110000",
32407 => "0011110100110000",
32408 => "0011110100110000",
32409 => "0011110100110000",
32410 => "0011110100111000",
32411 => "0011110100111000",
32412 => "0011110100111000",
32413 => "0011110100111000",
32414 => "0011110101000000",
32415 => "0011110101000000",
32416 => "0011110101000000",
32417 => "0011110101000000",
32418 => "0011110101001000",
32419 => "0011110101001000",
32420 => "0011110101001000",
32421 => "0011110101001000",
32422 => "0011110101010000",
32423 => "0011110101010000",
32424 => "0011110101010000",
32425 => "0011110101010000",
32426 => "0011110101011000",
32427 => "0011110101011000",
32428 => "0011110101011000",
32429 => "0011110101011000",
32430 => "0011110101100000",
32431 => "0011110101100000",
32432 => "0011110101100000",
32433 => "0011110101100000",
32434 => "0011110101101000",
32435 => "0011110101101000",
32436 => "0011110101101000",
32437 => "0011110101101000",
32438 => "0011110101110000",
32439 => "0011110101110000",
32440 => "0011110101110000",
32441 => "0011110101110000",
32442 => "0011110101111000",
32443 => "0011110101111000",
32444 => "0011110101111000",
32445 => "0011110101111000",
32446 => "0011110110000000",
32447 => "0011110110000000",
32448 => "0011110110000000",
32449 => "0011110110000000",
32450 => "0011110110001000",
32451 => "0011110110001000",
32452 => "0011110110001000",
32453 => "0011110110001000",
32454 => "0011110110010000",
32455 => "0011110110010000",
32456 => "0011110110010000",
32457 => "0011110110010000",
32458 => "0011110110011000",
32459 => "0011110110011000",
32460 => "0011110110011000",
32461 => "0011110110011000",
32462 => "0011110110100000",
32463 => "0011110110100000",
32464 => "0011110110100000",
32465 => "0011110110100000",
32466 => "0011110110101000",
32467 => "0011110110101000",
32468 => "0011110110101000",
32469 => "0011110110101000",
32470 => "0011110110110000",
32471 => "0011110110110000",
32472 => "0011110110110000",
32473 => "0011110110110000",
32474 => "0011110110111000",
32475 => "0011110110111000",
32476 => "0011110110111000",
32477 => "0011110110111000",
32478 => "0011110111000000",
32479 => "0011110111000000",
32480 => "0011110111000000",
32481 => "0011110111000000",
32482 => "0011110111001000",
32483 => "0011110111001000",
32484 => "0011110111001000",
32485 => "0011110111001000",
32486 => "0011110111010000",
32487 => "0011110111010000",
32488 => "0011110111010000",
32489 => "0011110111010000",
32490 => "0011110111011000",
32491 => "0011110111011000",
32492 => "0011110111011000",
32493 => "0011110111011000",
32494 => "0011110111100000",
32495 => "0011110111100000",
32496 => "0011110111100000",
32497 => "0011110111100000",
32498 => "0011110111101000",
32499 => "0011110111101000",
32500 => "0011110111101000",
32501 => "0011110111101000",
32502 => "0011110111110000",
32503 => "0011110111110000",
32504 => "0011110111110000",
32505 => "0011110111110000",
32506 => "0011110111111000",
32507 => "0011110111111000",
32508 => "0011110111111000",
32509 => "0011110111111000",
32510 => "0011111000000000",
32511 => "0011111000000000",
32512 => "0011111000000000",
32513 => "0011111000000000",
32514 => "0011111000001000",
32515 => "0011111000001000",
32516 => "0011111000001000",
32517 => "0011111000001000",
32518 => "0011111000010000",
32519 => "0011111000010000",
32520 => "0011111000010000",
32521 => "0011111000010000",
32522 => "0011111000011000",
32523 => "0011111000011000",
32524 => "0011111000011000",
32525 => "0011111000011000",
32526 => "0011111000100000",
32527 => "0011111000100000",
32528 => "0011111000100000",
32529 => "0011111000100000",
32530 => "0011111000101000",
32531 => "0011111000101000",
32532 => "0011111000101000",
32533 => "0011111000101000",
32534 => "0011111000110000",
32535 => "0011111000110000",
32536 => "0011111000110000",
32537 => "0011111000110000",
32538 => "0011111000111000",
32539 => "0011111000111000",
32540 => "0011111000111000",
32541 => "0011111000111000",
32542 => "0011111001000000",
32543 => "0011111001000000",
32544 => "0011111001000000",
32545 => "0011111001000000",
32546 => "0011111001001000",
32547 => "0011111001001000",
32548 => "0011111001001000",
32549 => "0011111001001000",
32550 => "0011111001010000",
32551 => "0011111001010000",
32552 => "0011111001010000",
32553 => "0011111001010000",
32554 => "0011111001011000",
32555 => "0011111001011000",
32556 => "0011111001011000",
32557 => "0011111001011000",
32558 => "0011111001100000",
32559 => "0011111001100000",
32560 => "0011111001100000",
32561 => "0011111001100000",
32562 => "0011111001101000",
32563 => "0011111001101000",
32564 => "0011111001101000",
32565 => "0011111001101000",
32566 => "0011111001110000",
32567 => "0011111001110000",
32568 => "0011111001110000",
32569 => "0011111001110000",
32570 => "0011111001111000",
32571 => "0011111001111000",
32572 => "0011111001111000",
32573 => "0011111001111000",
32574 => "0011111010000000",
32575 => "0011111010000000",
32576 => "0011111010000000",
32577 => "0011111010000000",
32578 => "0011111010001000",
32579 => "0011111010001000",
32580 => "0011111010001000",
32581 => "0011111010001000",
32582 => "0011111010010000",
32583 => "0011111010010000",
32584 => "0011111010010000",
32585 => "0011111010010000",
32586 => "0011111010011000",
32587 => "0011111010011000",
32588 => "0011111010011000",
32589 => "0011111010011000",
32590 => "0011111010100000",
32591 => "0011111010100000",
32592 => "0011111010100000",
32593 => "0011111010100000",
32594 => "0011111010101000",
32595 => "0011111010101000",
32596 => "0011111010101000",
32597 => "0011111010101000",
32598 => "0011111010110000",
32599 => "0011111010110000",
32600 => "0011111010110000",
32601 => "0011111010110000",
32602 => "0011111010111000",
32603 => "0011111010111000",
32604 => "0011111010111000",
32605 => "0011111010111000",
32606 => "0011111011000000",
32607 => "0011111011000000",
32608 => "0011111011000000",
32609 => "0011111011000000",
32610 => "0011111011001000",
32611 => "0011111011001000",
32612 => "0011111011001000",
32613 => "0011111011001000",
32614 => "0011111011010000",
32615 => "0011111011010000",
32616 => "0011111011010000",
32617 => "0011111011010000",
32618 => "0011111011011000",
32619 => "0011111011011000",
32620 => "0011111011011000",
32621 => "0011111011011000",
32622 => "0011111011100000",
32623 => "0011111011100000",
32624 => "0011111011100000",
32625 => "0011111011100000",
32626 => "0011111011101000",
32627 => "0011111011101000",
32628 => "0011111011101000",
32629 => "0011111011101000",
32630 => "0011111011110000",
32631 => "0011111011110000",
32632 => "0011111011110000",
32633 => "0011111011110000",
32634 => "0011111011111000",
32635 => "0011111011111000",
32636 => "0011111011111000",
32637 => "0011111011111000",
32638 => "0011111100000000",
32639 => "0011111100000000",
32640 => "0011111100000000",
32641 => "0011111100000000",
32642 => "0011111100001000",
32643 => "0011111100001000",
32644 => "0011111100001000",
32645 => "0011111100001000",
32646 => "0011111100010000",
32647 => "0011111100010000",
32648 => "0011111100010000",
32649 => "0011111100010000",
32650 => "0011111100011000",
32651 => "0011111100011000",
32652 => "0011111100011000",
32653 => "0011111100011000",
32654 => "0011111100100000",
32655 => "0011111100100000",
32656 => "0011111100100000",
32657 => "0011111100100000",
32658 => "0011111100101000",
32659 => "0011111100101000",
32660 => "0011111100101000",
32661 => "0011111100101000",
32662 => "0011111100110000",
32663 => "0011111100110000",
32664 => "0011111100110000",
32665 => "0011111100110000",
32666 => "0011111100111000",
32667 => "0011111100111000",
32668 => "0011111100111000",
32669 => "0011111100111000",
32670 => "0011111101000000",
32671 => "0011111101000000",
32672 => "0011111101000000",
32673 => "0011111101000000",
32674 => "0011111101001000",
32675 => "0011111101001000",
32676 => "0011111101001000",
32677 => "0011111101001000",
32678 => "0011111101010000",
32679 => "0011111101010000",
32680 => "0011111101010000",
32681 => "0011111101010000",
32682 => "0011111101011000",
32683 => "0011111101011000",
32684 => "0011111101011000",
32685 => "0011111101011000",
32686 => "0011111101100000",
32687 => "0011111101100000",
32688 => "0011111101100000",
32689 => "0011111101100000",
32690 => "0011111101101000",
32691 => "0011111101101000",
32692 => "0011111101101000",
32693 => "0011111101101000",
32694 => "0011111101110000",
32695 => "0011111101110000",
32696 => "0011111101110000",
32697 => "0011111101110000",
32698 => "0011111101111000",
32699 => "0011111101111000",
32700 => "0011111101111000",
32701 => "0011111101111000",
32702 => "0011111110000000",
32703 => "0011111110000000",
32704 => "0011111110000000",
32705 => "0011111110000000",
32706 => "0011111110001000",
32707 => "0011111110001000",
32708 => "0011111110001000",
32709 => "0011111110001000",
32710 => "0011111110010000",
32711 => "0011111110010000",
32712 => "0011111110010000",
32713 => "0011111110010000",
32714 => "0011111110011000",
32715 => "0011111110011000",
32716 => "0011111110011000",
32717 => "0011111110011000",
32718 => "0011111110100000",
32719 => "0011111110100000",
32720 => "0011111110100000",
32721 => "0011111110100000",
32722 => "0011111110101000",
32723 => "0011111110101000",
32724 => "0011111110101000",
32725 => "0011111110101000",
32726 => "0011111110110000",
32727 => "0011111110110000",
32728 => "0011111110110000",
32729 => "0011111110110000",
32730 => "0011111110111000",
32731 => "0011111110111000",
32732 => "0011111110111000",
32733 => "0011111110111000",
32734 => "0011111111000000",
32735 => "0011111111000000",
32736 => "0011111111000000",
32737 => "0011111111000000",
32738 => "0011111111001000",
32739 => "0011111111001000",
32740 => "0011111111001000",
32741 => "0011111111001000",
32742 => "0011111111010000",
32743 => "0011111111010000",
32744 => "0011111111010000",
32745 => "0011111111010000",
32746 => "0011111111011000",
32747 => "0011111111011000",
32748 => "0011111111011000",
32749 => "0011111111011000",
32750 => "0011111111100000",
32751 => "0011111111100000",
32752 => "0011111111100000",
32753 => "0011111111100000",
32754 => "0011111111101000",
32755 => "0011111111101000",
32756 => "0011111111101000",
32757 => "0011111111101000",
32758 => "0011111111110000",
32759 => "0011111111110000",
32760 => "0011111111110000",
32761 => "0011111111110000",
32762 => "0011111111111000",
32763 => "0011111111111000",
32764 => "0011111111111000",
32765 => "0011111111111000",
32766 => "0100000000000000",
32767 => "0100000000000000",
32768 => "0100000000000000",
32769 => "0100000000000000",
32770 => "0100000000000000",
32771 => "0100000000000000",
32772 => "0100000000010000",
32773 => "0100000000010000",
32774 => "0100000000010000",
32775 => "0100000000010000",
32776 => "0100000000010000",
32777 => "0100000000010000",
32778 => "0100000000010000",
32779 => "0100000000010000",
32780 => "0100000000100000",
32781 => "0100000000100000",
32782 => "0100000000100000",
32783 => "0100000000100000",
32784 => "0100000000100000",
32785 => "0100000000100000",
32786 => "0100000000100000",
32787 => "0100000000100000",
32788 => "0100000000110000",
32789 => "0100000000110000",
32790 => "0100000000110000",
32791 => "0100000000110000",
32792 => "0100000000110000",
32793 => "0100000000110000",
32794 => "0100000000110000",
32795 => "0100000000110000",
32796 => "0100000001000000",
32797 => "0100000001000000",
32798 => "0100000001000000",
32799 => "0100000001000000",
32800 => "0100000001000000",
32801 => "0100000001000000",
32802 => "0100000001000000",
32803 => "0100000001000000",
32804 => "0100000001010000",
32805 => "0100000001010000",
32806 => "0100000001010000",
32807 => "0100000001010000",
32808 => "0100000001010000",
32809 => "0100000001010000",
32810 => "0100000001010000",
32811 => "0100000001010000",
32812 => "0100000001100000",
32813 => "0100000001100000",
32814 => "0100000001100000",
32815 => "0100000001100000",
32816 => "0100000001100000",
32817 => "0100000001100000",
32818 => "0100000001100000",
32819 => "0100000001100000",
32820 => "0100000001110000",
32821 => "0100000001110000",
32822 => "0100000001110000",
32823 => "0100000001110000",
32824 => "0100000001110000",
32825 => "0100000001110000",
32826 => "0100000001110000",
32827 => "0100000001110000",
32828 => "0100000010000000",
32829 => "0100000010000000",
32830 => "0100000010000000",
32831 => "0100000010000000",
32832 => "0100000010000000",
32833 => "0100000010000000",
32834 => "0100000010000000",
32835 => "0100000010000000",
32836 => "0100000010010000",
32837 => "0100000010010000",
32838 => "0100000010010000",
32839 => "0100000010010000",
32840 => "0100000010010000",
32841 => "0100000010010000",
32842 => "0100000010010000",
32843 => "0100000010010000",
32844 => "0100000010100000",
32845 => "0100000010100000",
32846 => "0100000010100000",
32847 => "0100000010100000",
32848 => "0100000010100000",
32849 => "0100000010100000",
32850 => "0100000010100000",
32851 => "0100000010100000",
32852 => "0100000010110000",
32853 => "0100000010110000",
32854 => "0100000010110000",
32855 => "0100000010110000",
32856 => "0100000010110000",
32857 => "0100000010110000",
32858 => "0100000010110000",
32859 => "0100000010110000",
32860 => "0100000011000000",
32861 => "0100000011000000",
32862 => "0100000011000000",
32863 => "0100000011000000",
32864 => "0100000011000000",
32865 => "0100000011000000",
32866 => "0100000011000000",
32867 => "0100000011000000",
32868 => "0100000011010000",
32869 => "0100000011010000",
32870 => "0100000011010000",
32871 => "0100000011010000",
32872 => "0100000011010000",
32873 => "0100000011010000",
32874 => "0100000011010000",
32875 => "0100000011010000",
32876 => "0100000011100000",
32877 => "0100000011100000",
32878 => "0100000011100000",
32879 => "0100000011100000",
32880 => "0100000011100000",
32881 => "0100000011100000",
32882 => "0100000011100000",
32883 => "0100000011100000",
32884 => "0100000011110000",
32885 => "0100000011110000",
32886 => "0100000011110000",
32887 => "0100000011110000",
32888 => "0100000011110000",
32889 => "0100000011110000",
32890 => "0100000011110000",
32891 => "0100000011110000",
32892 => "0100000100000000",
32893 => "0100000100000000",
32894 => "0100000100000000",
32895 => "0100000100000000",
32896 => "0100000100000000",
32897 => "0100000100000000",
32898 => "0100000100000000",
32899 => "0100000100000000",
32900 => "0100000100010000",
32901 => "0100000100010000",
32902 => "0100000100010000",
32903 => "0100000100010000",
32904 => "0100000100010000",
32905 => "0100000100010000",
32906 => "0100000100010000",
32907 => "0100000100010000",
32908 => "0100000100100000",
32909 => "0100000100100000",
32910 => "0100000100100000",
32911 => "0100000100100000",
32912 => "0100000100100000",
32913 => "0100000100100000",
32914 => "0100000100100000",
32915 => "0100000100100000",
32916 => "0100000100110000",
32917 => "0100000100110000",
32918 => "0100000100110000",
32919 => "0100000100110000",
32920 => "0100000100110000",
32921 => "0100000100110000",
32922 => "0100000100110000",
32923 => "0100000100110000",
32924 => "0100000101000000",
32925 => "0100000101000000",
32926 => "0100000101000000",
32927 => "0100000101000000",
32928 => "0100000101000000",
32929 => "0100000101000000",
32930 => "0100000101000000",
32931 => "0100000101000000",
32932 => "0100000101010000",
32933 => "0100000101010000",
32934 => "0100000101010000",
32935 => "0100000101010000",
32936 => "0100000101010000",
32937 => "0100000101010000",
32938 => "0100000101010000",
32939 => "0100000101010000",
32940 => "0100000101100000",
32941 => "0100000101100000",
32942 => "0100000101100000",
32943 => "0100000101100000",
32944 => "0100000101100000",
32945 => "0100000101100000",
32946 => "0100000101100000",
32947 => "0100000101100000",
32948 => "0100000101110000",
32949 => "0100000101110000",
32950 => "0100000101110000",
32951 => "0100000101110000",
32952 => "0100000101110000",
32953 => "0100000101110000",
32954 => "0100000101110000",
32955 => "0100000101110000",
32956 => "0100000110000000",
32957 => "0100000110000000",
32958 => "0100000110000000",
32959 => "0100000110000000",
32960 => "0100000110000000",
32961 => "0100000110000000",
32962 => "0100000110000000",
32963 => "0100000110000000",
32964 => "0100000110010000",
32965 => "0100000110010000",
32966 => "0100000110010000",
32967 => "0100000110010000",
32968 => "0100000110010000",
32969 => "0100000110010000",
32970 => "0100000110010000",
32971 => "0100000110010000",
32972 => "0100000110100000",
32973 => "0100000110100000",
32974 => "0100000110100000",
32975 => "0100000110100000",
32976 => "0100000110100000",
32977 => "0100000110100000",
32978 => "0100000110100000",
32979 => "0100000110100000",
32980 => "0100000110110000",
32981 => "0100000110110000",
32982 => "0100000110110000",
32983 => "0100000110110000",
32984 => "0100000110110000",
32985 => "0100000110110000",
32986 => "0100000110110000",
32987 => "0100000110110000",
32988 => "0100000111000000",
32989 => "0100000111000000",
32990 => "0100000111000000",
32991 => "0100000111000000",
32992 => "0100000111000000",
32993 => "0100000111000000",
32994 => "0100000111000000",
32995 => "0100000111000000",
32996 => "0100000111010000",
32997 => "0100000111010000",
32998 => "0100000111010000",
32999 => "0100000111010000",
33000 => "0100000111010000",
33001 => "0100000111010000",
33002 => "0100000111010000",
33003 => "0100000111010000",
33004 => "0100000111100000",
33005 => "0100000111100000",
33006 => "0100000111100000",
33007 => "0100000111100000",
33008 => "0100000111100000",
33009 => "0100000111100000",
33010 => "0100000111100000",
33011 => "0100000111100000",
33012 => "0100000111110000",
33013 => "0100000111110000",
33014 => "0100000111110000",
33015 => "0100000111110000",
33016 => "0100000111110000",
33017 => "0100000111110000",
33018 => "0100000111110000",
33019 => "0100000111110000",
33020 => "0100001000000000",
33021 => "0100001000000000",
33022 => "0100001000000000",
33023 => "0100001000000000",
33024 => "0100001000000000",
33025 => "0100001000000000",
33026 => "0100001000000000",
33027 => "0100001000000000",
33028 => "0100001000010000",
33029 => "0100001000010000",
33030 => "0100001000010000",
33031 => "0100001000010000",
33032 => "0100001000010000",
33033 => "0100001000010000",
33034 => "0100001000010000",
33035 => "0100001000010000",
33036 => "0100001000100000",
33037 => "0100001000100000",
33038 => "0100001000100000",
33039 => "0100001000100000",
33040 => "0100001000100000",
33041 => "0100001000100000",
33042 => "0100001000100000",
33043 => "0100001000100000",
33044 => "0100001000110000",
33045 => "0100001000110000",
33046 => "0100001000110000",
33047 => "0100001000110000",
33048 => "0100001000110000",
33049 => "0100001000110000",
33050 => "0100001000110000",
33051 => "0100001000110000",
33052 => "0100001001000000",
33053 => "0100001001000000",
33054 => "0100001001000000",
33055 => "0100001001000000",
33056 => "0100001001000000",
33057 => "0100001001000000",
33058 => "0100001001000000",
33059 => "0100001001000000",
33060 => "0100001001010000",
33061 => "0100001001010000",
33062 => "0100001001010000",
33063 => "0100001001010000",
33064 => "0100001001010000",
33065 => "0100001001010000",
33066 => "0100001001010000",
33067 => "0100001001010000",
33068 => "0100001001100000",
33069 => "0100001001100000",
33070 => "0100001001100000",
33071 => "0100001001100000",
33072 => "0100001001100000",
33073 => "0100001001100000",
33074 => "0100001001100000",
33075 => "0100001001100000",
33076 => "0100001001110000",
33077 => "0100001001110000",
33078 => "0100001001110000",
33079 => "0100001001110000",
33080 => "0100001001110000",
33081 => "0100001001110000",
33082 => "0100001001110000",
33083 => "0100001001110000",
33084 => "0100001010000000",
33085 => "0100001010000000",
33086 => "0100001010000000",
33087 => "0100001010000000",
33088 => "0100001010000000",
33089 => "0100001010000000",
33090 => "0100001010000000",
33091 => "0100001010000000",
33092 => "0100001010010000",
33093 => "0100001010010000",
33094 => "0100001010010000",
33095 => "0100001010010000",
33096 => "0100001010010000",
33097 => "0100001010010000",
33098 => "0100001010010000",
33099 => "0100001010010000",
33100 => "0100001010100000",
33101 => "0100001010100000",
33102 => "0100001010100000",
33103 => "0100001010100000",
33104 => "0100001010100000",
33105 => "0100001010100000",
33106 => "0100001010100000",
33107 => "0100001010100000",
33108 => "0100001010110000",
33109 => "0100001010110000",
33110 => "0100001010110000",
33111 => "0100001010110000",
33112 => "0100001010110000",
33113 => "0100001010110000",
33114 => "0100001010110000",
33115 => "0100001010110000",
33116 => "0100001011000000",
33117 => "0100001011000000",
33118 => "0100001011000000",
33119 => "0100001011000000",
33120 => "0100001011000000",
33121 => "0100001011000000",
33122 => "0100001011000000",
33123 => "0100001011000000",
33124 => "0100001011010000",
33125 => "0100001011010000",
33126 => "0100001011010000",
33127 => "0100001011010000",
33128 => "0100001011010000",
33129 => "0100001011010000",
33130 => "0100001011010000",
33131 => "0100001011010000",
33132 => "0100001011100000",
33133 => "0100001011100000",
33134 => "0100001011100000",
33135 => "0100001011100000",
33136 => "0100001011100000",
33137 => "0100001011100000",
33138 => "0100001011100000",
33139 => "0100001011100000",
33140 => "0100001011110000",
33141 => "0100001011110000",
33142 => "0100001011110000",
33143 => "0100001011110000",
33144 => "0100001011110000",
33145 => "0100001011110000",
33146 => "0100001011110000",
33147 => "0100001011110000",
33148 => "0100001100000000",
33149 => "0100001100000000",
33150 => "0100001100000000",
33151 => "0100001100000000",
33152 => "0100001100000000",
33153 => "0100001100000000",
33154 => "0100001100000000",
33155 => "0100001100000000",
33156 => "0100001100010000",
33157 => "0100001100010000",
33158 => "0100001100010000",
33159 => "0100001100010000",
33160 => "0100001100010000",
33161 => "0100001100010000",
33162 => "0100001100010000",
33163 => "0100001100010000",
33164 => "0100001100100000",
33165 => "0100001100100000",
33166 => "0100001100100000",
33167 => "0100001100100000",
33168 => "0100001100100000",
33169 => "0100001100100000",
33170 => "0100001100100000",
33171 => "0100001100100000",
33172 => "0100001100110000",
33173 => "0100001100110000",
33174 => "0100001100110000",
33175 => "0100001100110000",
33176 => "0100001100110000",
33177 => "0100001100110000",
33178 => "0100001100110000",
33179 => "0100001100110000",
33180 => "0100001101000000",
33181 => "0100001101000000",
33182 => "0100001101000000",
33183 => "0100001101000000",
33184 => "0100001101000000",
33185 => "0100001101000000",
33186 => "0100001101000000",
33187 => "0100001101000000",
33188 => "0100001101010000",
33189 => "0100001101010000",
33190 => "0100001101010000",
33191 => "0100001101010000",
33192 => "0100001101010000",
33193 => "0100001101010000",
33194 => "0100001101010000",
33195 => "0100001101010000",
33196 => "0100001101100000",
33197 => "0100001101100000",
33198 => "0100001101100000",
33199 => "0100001101100000",
33200 => "0100001101100000",
33201 => "0100001101100000",
33202 => "0100001101100000",
33203 => "0100001101100000",
33204 => "0100001101110000",
33205 => "0100001101110000",
33206 => "0100001101110000",
33207 => "0100001101110000",
33208 => "0100001101110000",
33209 => "0100001101110000",
33210 => "0100001101110000",
33211 => "0100001101110000",
33212 => "0100001110000000",
33213 => "0100001110000000",
33214 => "0100001110000000",
33215 => "0100001110000000",
33216 => "0100001110000000",
33217 => "0100001110000000",
33218 => "0100001110000000",
33219 => "0100001110000000",
33220 => "0100001110010000",
33221 => "0100001110010000",
33222 => "0100001110010000",
33223 => "0100001110010000",
33224 => "0100001110010000",
33225 => "0100001110010000",
33226 => "0100001110010000",
33227 => "0100001110010000",
33228 => "0100001110100000",
33229 => "0100001110100000",
33230 => "0100001110100000",
33231 => "0100001110100000",
33232 => "0100001110100000",
33233 => "0100001110100000",
33234 => "0100001110100000",
33235 => "0100001110100000",
33236 => "0100001110100000",
33237 => "0100001110110000",
33238 => "0100001110110000",
33239 => "0100001110110000",
33240 => "0100001110110000",
33241 => "0100001110110000",
33242 => "0100001110110000",
33243 => "0100001110110000",
33244 => "0100001110110000",
33245 => "0100001111000000",
33246 => "0100001111000000",
33247 => "0100001111000000",
33248 => "0100001111000000",
33249 => "0100001111000000",
33250 => "0100001111000000",
33251 => "0100001111000000",
33252 => "0100001111000000",
33253 => "0100001111010000",
33254 => "0100001111010000",
33255 => "0100001111010000",
33256 => "0100001111010000",
33257 => "0100001111010000",
33258 => "0100001111010000",
33259 => "0100001111010000",
33260 => "0100001111010000",
33261 => "0100001111100000",
33262 => "0100001111100000",
33263 => "0100001111100000",
33264 => "0100001111100000",
33265 => "0100001111100000",
33266 => "0100001111100000",
33267 => "0100001111100000",
33268 => "0100001111100000",
33269 => "0100001111110000",
33270 => "0100001111110000",
33271 => "0100001111110000",
33272 => "0100001111110000",
33273 => "0100001111110000",
33274 => "0100001111110000",
33275 => "0100001111110000",
33276 => "0100001111110000",
33277 => "0100010000000000",
33278 => "0100010000000000",
33279 => "0100010000000000",
33280 => "0100010000000000",
33281 => "0100010000000000",
33282 => "0100010000000000",
33283 => "0100010000000000",
33284 => "0100010000000000",
33285 => "0100010000010000",
33286 => "0100010000010000",
33287 => "0100010000010000",
33288 => "0100010000010000",
33289 => "0100010000010000",
33290 => "0100010000010000",
33291 => "0100010000010000",
33292 => "0100010000010000",
33293 => "0100010000100000",
33294 => "0100010000100000",
33295 => "0100010000100000",
33296 => "0100010000100000",
33297 => "0100010000100000",
33298 => "0100010000100000",
33299 => "0100010000100000",
33300 => "0100010000100000",
33301 => "0100010000110000",
33302 => "0100010000110000",
33303 => "0100010000110000",
33304 => "0100010000110000",
33305 => "0100010000110000",
33306 => "0100010000110000",
33307 => "0100010000110000",
33308 => "0100010000110000",
33309 => "0100010001000000",
33310 => "0100010001000000",
33311 => "0100010001000000",
33312 => "0100010001000000",
33313 => "0100010001000000",
33314 => "0100010001000000",
33315 => "0100010001000000",
33316 => "0100010001000000",
33317 => "0100010001010000",
33318 => "0100010001010000",
33319 => "0100010001010000",
33320 => "0100010001010000",
33321 => "0100010001010000",
33322 => "0100010001010000",
33323 => "0100010001010000",
33324 => "0100010001010000",
33325 => "0100010001100000",
33326 => "0100010001100000",
33327 => "0100010001100000",
33328 => "0100010001100000",
33329 => "0100010001100000",
33330 => "0100010001100000",
33331 => "0100010001100000",
33332 => "0100010001100000",
33333 => "0100010001110000",
33334 => "0100010001110000",
33335 => "0100010001110000",
33336 => "0100010001110000",
33337 => "0100010001110000",
33338 => "0100010001110000",
33339 => "0100010001110000",
33340 => "0100010001110000",
33341 => "0100010010000000",
33342 => "0100010010000000",
33343 => "0100010010000000",
33344 => "0100010010000000",
33345 => "0100010010000000",
33346 => "0100010010000000",
33347 => "0100010010000000",
33348 => "0100010010000000",
33349 => "0100010010010000",
33350 => "0100010010010000",
33351 => "0100010010010000",
33352 => "0100010010010000",
33353 => "0100010010010000",
33354 => "0100010010010000",
33355 => "0100010010010000",
33356 => "0100010010010000",
33357 => "0100010010100000",
33358 => "0100010010100000",
33359 => "0100010010100000",
33360 => "0100010010100000",
33361 => "0100010010100000",
33362 => "0100010010100000",
33363 => "0100010010100000",
33364 => "0100010010100000",
33365 => "0100010010110000",
33366 => "0100010010110000",
33367 => "0100010010110000",
33368 => "0100010010110000",
33369 => "0100010010110000",
33370 => "0100010010110000",
33371 => "0100010010110000",
33372 => "0100010010110000",
33373 => "0100010011000000",
33374 => "0100010011000000",
33375 => "0100010011000000",
33376 => "0100010011000000",
33377 => "0100010011000000",
33378 => "0100010011000000",
33379 => "0100010011000000",
33380 => "0100010011000000",
33381 => "0100010011010000",
33382 => "0100010011010000",
33383 => "0100010011010000",
33384 => "0100010011010000",
33385 => "0100010011010000",
33386 => "0100010011010000",
33387 => "0100010011010000",
33388 => "0100010011010000",
33389 => "0100010011100000",
33390 => "0100010011100000",
33391 => "0100010011100000",
33392 => "0100010011100000",
33393 => "0100010011100000",
33394 => "0100010011100000",
33395 => "0100010011100000",
33396 => "0100010011100000",
33397 => "0100010011110000",
33398 => "0100010011110000",
33399 => "0100010011110000",
33400 => "0100010011110000",
33401 => "0100010011110000",
33402 => "0100010011110000",
33403 => "0100010011110000",
33404 => "0100010011110000",
33405 => "0100010100000000",
33406 => "0100010100000000",
33407 => "0100010100000000",
33408 => "0100010100000000",
33409 => "0100010100000000",
33410 => "0100010100000000",
33411 => "0100010100000000",
33412 => "0100010100000000",
33413 => "0100010100010000",
33414 => "0100010100010000",
33415 => "0100010100010000",
33416 => "0100010100010000",
33417 => "0100010100010000",
33418 => "0100010100010000",
33419 => "0100010100010000",
33420 => "0100010100010000",
33421 => "0100010100100000",
33422 => "0100010100100000",
33423 => "0100010100100000",
33424 => "0100010100100000",
33425 => "0100010100100000",
33426 => "0100010100100000",
33427 => "0100010100100000",
33428 => "0100010100100000",
33429 => "0100010100110000",
33430 => "0100010100110000",
33431 => "0100010100110000",
33432 => "0100010100110000",
33433 => "0100010100110000",
33434 => "0100010100110000",
33435 => "0100010100110000",
33436 => "0100010100110000",
33437 => "0100010101000000",
33438 => "0100010101000000",
33439 => "0100010101000000",
33440 => "0100010101000000",
33441 => "0100010101000000",
33442 => "0100010101000000",
33443 => "0100010101000000",
33444 => "0100010101000000",
33445 => "0100010101000000",
33446 => "0100010101010000",
33447 => "0100010101010000",
33448 => "0100010101010000",
33449 => "0100010101010000",
33450 => "0100010101010000",
33451 => "0100010101010000",
33452 => "0100010101010000",
33453 => "0100010101010000",
33454 => "0100010101100000",
33455 => "0100010101100000",
33456 => "0100010101100000",
33457 => "0100010101100000",
33458 => "0100010101100000",
33459 => "0100010101100000",
33460 => "0100010101100000",
33461 => "0100010101100000",
33462 => "0100010101110000",
33463 => "0100010101110000",
33464 => "0100010101110000",
33465 => "0100010101110000",
33466 => "0100010101110000",
33467 => "0100010101110000",
33468 => "0100010101110000",
33469 => "0100010101110000",
33470 => "0100010110000000",
33471 => "0100010110000000",
33472 => "0100010110000000",
33473 => "0100010110000000",
33474 => "0100010110000000",
33475 => "0100010110000000",
33476 => "0100010110000000",
33477 => "0100010110000000",
33478 => "0100010110010000",
33479 => "0100010110010000",
33480 => "0100010110010000",
33481 => "0100010110010000",
33482 => "0100010110010000",
33483 => "0100010110010000",
33484 => "0100010110010000",
33485 => "0100010110010000",
33486 => "0100010110100000",
33487 => "0100010110100000",
33488 => "0100010110100000",
33489 => "0100010110100000",
33490 => "0100010110100000",
33491 => "0100010110100000",
33492 => "0100010110100000",
33493 => "0100010110100000",
33494 => "0100010110110000",
33495 => "0100010110110000",
33496 => "0100010110110000",
33497 => "0100010110110000",
33498 => "0100010110110000",
33499 => "0100010110110000",
33500 => "0100010110110000",
33501 => "0100010110110000",
33502 => "0100010111000000",
33503 => "0100010111000000",
33504 => "0100010111000000",
33505 => "0100010111000000",
33506 => "0100010111000000",
33507 => "0100010111000000",
33508 => "0100010111000000",
33509 => "0100010111000000",
33510 => "0100010111010000",
33511 => "0100010111010000",
33512 => "0100010111010000",
33513 => "0100010111010000",
33514 => "0100010111010000",
33515 => "0100010111010000",
33516 => "0100010111010000",
33517 => "0100010111010000",
33518 => "0100010111100000",
33519 => "0100010111100000",
33520 => "0100010111100000",
33521 => "0100010111100000",
33522 => "0100010111100000",
33523 => "0100010111100000",
33524 => "0100010111100000",
33525 => "0100010111100000",
33526 => "0100010111110000",
33527 => "0100010111110000",
33528 => "0100010111110000",
33529 => "0100010111110000",
33530 => "0100010111110000",
33531 => "0100010111110000",
33532 => "0100010111110000",
33533 => "0100010111110000",
33534 => "0100011000000000",
33535 => "0100011000000000",
33536 => "0100011000000000",
33537 => "0100011000000000",
33538 => "0100011000000000",
33539 => "0100011000000000",
33540 => "0100011000000000",
33541 => "0100011000000000",
33542 => "0100011000010000",
33543 => "0100011000010000",
33544 => "0100011000010000",
33545 => "0100011000010000",
33546 => "0100011000010000",
33547 => "0100011000010000",
33548 => "0100011000010000",
33549 => "0100011000010000",
33550 => "0100011000100000",
33551 => "0100011000100000",
33552 => "0100011000100000",
33553 => "0100011000100000",
33554 => "0100011000100000",
33555 => "0100011000100000",
33556 => "0100011000100000",
33557 => "0100011000100000",
33558 => "0100011000110000",
33559 => "0100011000110000",
33560 => "0100011000110000",
33561 => "0100011000110000",
33562 => "0100011000110000",
33563 => "0100011000110000",
33564 => "0100011000110000",
33565 => "0100011000110000",
33566 => "0100011000110000",
33567 => "0100011001000000",
33568 => "0100011001000000",
33569 => "0100011001000000",
33570 => "0100011001000000",
33571 => "0100011001000000",
33572 => "0100011001000000",
33573 => "0100011001000000",
33574 => "0100011001000000",
33575 => "0100011001010000",
33576 => "0100011001010000",
33577 => "0100011001010000",
33578 => "0100011001010000",
33579 => "0100011001010000",
33580 => "0100011001010000",
33581 => "0100011001010000",
33582 => "0100011001010000",
33583 => "0100011001100000",
33584 => "0100011001100000",
33585 => "0100011001100000",
33586 => "0100011001100000",
33587 => "0100011001100000",
33588 => "0100011001100000",
33589 => "0100011001100000",
33590 => "0100011001100000",
33591 => "0100011001110000",
33592 => "0100011001110000",
33593 => "0100011001110000",
33594 => "0100011001110000",
33595 => "0100011001110000",
33596 => "0100011001110000",
33597 => "0100011001110000",
33598 => "0100011001110000",
33599 => "0100011010000000",
33600 => "0100011010000000",
33601 => "0100011010000000",
33602 => "0100011010000000",
33603 => "0100011010000000",
33604 => "0100011010000000",
33605 => "0100011010000000",
33606 => "0100011010000000",
33607 => "0100011010010000",
33608 => "0100011010010000",
33609 => "0100011010010000",
33610 => "0100011010010000",
33611 => "0100011010010000",
33612 => "0100011010010000",
33613 => "0100011010010000",
33614 => "0100011010010000",
33615 => "0100011010100000",
33616 => "0100011010100000",
33617 => "0100011010100000",
33618 => "0100011010100000",
33619 => "0100011010100000",
33620 => "0100011010100000",
33621 => "0100011010100000",
33622 => "0100011010100000",
33623 => "0100011010110000",
33624 => "0100011010110000",
33625 => "0100011010110000",
33626 => "0100011010110000",
33627 => "0100011010110000",
33628 => "0100011010110000",
33629 => "0100011010110000",
33630 => "0100011010110000",
33631 => "0100011011000000",
33632 => "0100011011000000",
33633 => "0100011011000000",
33634 => "0100011011000000",
33635 => "0100011011000000",
33636 => "0100011011000000",
33637 => "0100011011000000",
33638 => "0100011011000000",
33639 => "0100011011010000",
33640 => "0100011011010000",
33641 => "0100011011010000",
33642 => "0100011011010000",
33643 => "0100011011010000",
33644 => "0100011011010000",
33645 => "0100011011010000",
33646 => "0100011011010000",
33647 => "0100011011100000",
33648 => "0100011011100000",
33649 => "0100011011100000",
33650 => "0100011011100000",
33651 => "0100011011100000",
33652 => "0100011011100000",
33653 => "0100011011100000",
33654 => "0100011011100000",
33655 => "0100011011110000",
33656 => "0100011011110000",
33657 => "0100011011110000",
33658 => "0100011011110000",
33659 => "0100011011110000",
33660 => "0100011011110000",
33661 => "0100011011110000",
33662 => "0100011011110000",
33663 => "0100011011110000",
33664 => "0100011100000000",
33665 => "0100011100000000",
33666 => "0100011100000000",
33667 => "0100011100000000",
33668 => "0100011100000000",
33669 => "0100011100000000",
33670 => "0100011100000000",
33671 => "0100011100000000",
33672 => "0100011100010000",
33673 => "0100011100010000",
33674 => "0100011100010000",
33675 => "0100011100010000",
33676 => "0100011100010000",
33677 => "0100011100010000",
33678 => "0100011100010000",
33679 => "0100011100010000",
33680 => "0100011100100000",
33681 => "0100011100100000",
33682 => "0100011100100000",
33683 => "0100011100100000",
33684 => "0100011100100000",
33685 => "0100011100100000",
33686 => "0100011100100000",
33687 => "0100011100100000",
33688 => "0100011100110000",
33689 => "0100011100110000",
33690 => "0100011100110000",
33691 => "0100011100110000",
33692 => "0100011100110000",
33693 => "0100011100110000",
33694 => "0100011100110000",
33695 => "0100011100110000",
33696 => "0100011101000000",
33697 => "0100011101000000",
33698 => "0100011101000000",
33699 => "0100011101000000",
33700 => "0100011101000000",
33701 => "0100011101000000",
33702 => "0100011101000000",
33703 => "0100011101000000",
33704 => "0100011101010000",
33705 => "0100011101010000",
33706 => "0100011101010000",
33707 => "0100011101010000",
33708 => "0100011101010000",
33709 => "0100011101010000",
33710 => "0100011101010000",
33711 => "0100011101010000",
33712 => "0100011101100000",
33713 => "0100011101100000",
33714 => "0100011101100000",
33715 => "0100011101100000",
33716 => "0100011101100000",
33717 => "0100011101100000",
33718 => "0100011101100000",
33719 => "0100011101100000",
33720 => "0100011101110000",
33721 => "0100011101110000",
33722 => "0100011101110000",
33723 => "0100011101110000",
33724 => "0100011101110000",
33725 => "0100011101110000",
33726 => "0100011101110000",
33727 => "0100011101110000",
33728 => "0100011110000000",
33729 => "0100011110000000",
33730 => "0100011110000000",
33731 => "0100011110000000",
33732 => "0100011110000000",
33733 => "0100011110000000",
33734 => "0100011110000000",
33735 => "0100011110000000",
33736 => "0100011110010000",
33737 => "0100011110010000",
33738 => "0100011110010000",
33739 => "0100011110010000",
33740 => "0100011110010000",
33741 => "0100011110010000",
33742 => "0100011110010000",
33743 => "0100011110010000",
33744 => "0100011110010000",
33745 => "0100011110100000",
33746 => "0100011110100000",
33747 => "0100011110100000",
33748 => "0100011110100000",
33749 => "0100011110100000",
33750 => "0100011110100000",
33751 => "0100011110100000",
33752 => "0100011110100000",
33753 => "0100011110110000",
33754 => "0100011110110000",
33755 => "0100011110110000",
33756 => "0100011110110000",
33757 => "0100011110110000",
33758 => "0100011110110000",
33759 => "0100011110110000",
33760 => "0100011110110000",
33761 => "0100011111000000",
33762 => "0100011111000000",
33763 => "0100011111000000",
33764 => "0100011111000000",
33765 => "0100011111000000",
33766 => "0100011111000000",
33767 => "0100011111000000",
33768 => "0100011111000000",
33769 => "0100011111010000",
33770 => "0100011111010000",
33771 => "0100011111010000",
33772 => "0100011111010000",
33773 => "0100011111010000",
33774 => "0100011111010000",
33775 => "0100011111010000",
33776 => "0100011111010000",
33777 => "0100011111100000",
33778 => "0100011111100000",
33779 => "0100011111100000",
33780 => "0100011111100000",
33781 => "0100011111100000",
33782 => "0100011111100000",
33783 => "0100011111100000",
33784 => "0100011111100000",
33785 => "0100011111110000",
33786 => "0100011111110000",
33787 => "0100011111110000",
33788 => "0100011111110000",
33789 => "0100011111110000",
33790 => "0100011111110000",
33791 => "0100011111110000",
33792 => "0100011111110000",
33793 => "0100100000000000",
33794 => "0100100000000000",
33795 => "0100100000000000",
33796 => "0100100000000000",
33797 => "0100100000000000",
33798 => "0100100000000000",
33799 => "0100100000000000",
33800 => "0100100000000000",
33801 => "0100100000010000",
33802 => "0100100000010000",
33803 => "0100100000010000",
33804 => "0100100000010000",
33805 => "0100100000010000",
33806 => "0100100000010000",
33807 => "0100100000010000",
33808 => "0100100000010000",
33809 => "0100100000010000",
33810 => "0100100000100000",
33811 => "0100100000100000",
33812 => "0100100000100000",
33813 => "0100100000100000",
33814 => "0100100000100000",
33815 => "0100100000100000",
33816 => "0100100000100000",
33817 => "0100100000100000",
33818 => "0100100000110000",
33819 => "0100100000110000",
33820 => "0100100000110000",
33821 => "0100100000110000",
33822 => "0100100000110000",
33823 => "0100100000110000",
33824 => "0100100000110000",
33825 => "0100100000110000",
33826 => "0100100001000000",
33827 => "0100100001000000",
33828 => "0100100001000000",
33829 => "0100100001000000",
33830 => "0100100001000000",
33831 => "0100100001000000",
33832 => "0100100001000000",
33833 => "0100100001000000",
33834 => "0100100001010000",
33835 => "0100100001010000",
33836 => "0100100001010000",
33837 => "0100100001010000",
33838 => "0100100001010000",
33839 => "0100100001010000",
33840 => "0100100001010000",
33841 => "0100100001010000",
33842 => "0100100001100000",
33843 => "0100100001100000",
33844 => "0100100001100000",
33845 => "0100100001100000",
33846 => "0100100001100000",
33847 => "0100100001100000",
33848 => "0100100001100000",
33849 => "0100100001100000",
33850 => "0100100001110000",
33851 => "0100100001110000",
33852 => "0100100001110000",
33853 => "0100100001110000",
33854 => "0100100001110000",
33855 => "0100100001110000",
33856 => "0100100001110000",
33857 => "0100100001110000",
33858 => "0100100010000000",
33859 => "0100100010000000",
33860 => "0100100010000000",
33861 => "0100100010000000",
33862 => "0100100010000000",
33863 => "0100100010000000",
33864 => "0100100010000000",
33865 => "0100100010000000",
33866 => "0100100010000000",
33867 => "0100100010010000",
33868 => "0100100010010000",
33869 => "0100100010010000",
33870 => "0100100010010000",
33871 => "0100100010010000",
33872 => "0100100010010000",
33873 => "0100100010010000",
33874 => "0100100010010000",
33875 => "0100100010100000",
33876 => "0100100010100000",
33877 => "0100100010100000",
33878 => "0100100010100000",
33879 => "0100100010100000",
33880 => "0100100010100000",
33881 => "0100100010100000",
33882 => "0100100010100000",
33883 => "0100100010110000",
33884 => "0100100010110000",
33885 => "0100100010110000",
33886 => "0100100010110000",
33887 => "0100100010110000",
33888 => "0100100010110000",
33889 => "0100100010110000",
33890 => "0100100010110000",
33891 => "0100100011000000",
33892 => "0100100011000000",
33893 => "0100100011000000",
33894 => "0100100011000000",
33895 => "0100100011000000",
33896 => "0100100011000000",
33897 => "0100100011000000",
33898 => "0100100011000000",
33899 => "0100100011010000",
33900 => "0100100011010000",
33901 => "0100100011010000",
33902 => "0100100011010000",
33903 => "0100100011010000",
33904 => "0100100011010000",
33905 => "0100100011010000",
33906 => "0100100011010000",
33907 => "0100100011100000",
33908 => "0100100011100000",
33909 => "0100100011100000",
33910 => "0100100011100000",
33911 => "0100100011100000",
33912 => "0100100011100000",
33913 => "0100100011100000",
33914 => "0100100011100000",
33915 => "0100100011110000",
33916 => "0100100011110000",
33917 => "0100100011110000",
33918 => "0100100011110000",
33919 => "0100100011110000",
33920 => "0100100011110000",
33921 => "0100100011110000",
33922 => "0100100011110000",
33923 => "0100100011110000",
33924 => "0100100100000000",
33925 => "0100100100000000",
33926 => "0100100100000000",
33927 => "0100100100000000",
33928 => "0100100100000000",
33929 => "0100100100000000",
33930 => "0100100100000000",
33931 => "0100100100000000",
33932 => "0100100100010000",
33933 => "0100100100010000",
33934 => "0100100100010000",
33935 => "0100100100010000",
33936 => "0100100100010000",
33937 => "0100100100010000",
33938 => "0100100100010000",
33939 => "0100100100010000",
33940 => "0100100100100000",
33941 => "0100100100100000",
33942 => "0100100100100000",
33943 => "0100100100100000",
33944 => "0100100100100000",
33945 => "0100100100100000",
33946 => "0100100100100000",
33947 => "0100100100100000",
33948 => "0100100100110000",
33949 => "0100100100110000",
33950 => "0100100100110000",
33951 => "0100100100110000",
33952 => "0100100100110000",
33953 => "0100100100110000",
33954 => "0100100100110000",
33955 => "0100100100110000",
33956 => "0100100101000000",
33957 => "0100100101000000",
33958 => "0100100101000000",
33959 => "0100100101000000",
33960 => "0100100101000000",
33961 => "0100100101000000",
33962 => "0100100101000000",
33963 => "0100100101000000",
33964 => "0100100101010000",
33965 => "0100100101010000",
33966 => "0100100101010000",
33967 => "0100100101010000",
33968 => "0100100101010000",
33969 => "0100100101010000",
33970 => "0100100101010000",
33971 => "0100100101010000",
33972 => "0100100101010000",
33973 => "0100100101100000",
33974 => "0100100101100000",
33975 => "0100100101100000",
33976 => "0100100101100000",
33977 => "0100100101100000",
33978 => "0100100101100000",
33979 => "0100100101100000",
33980 => "0100100101100000",
33981 => "0100100101110000",
33982 => "0100100101110000",
33983 => "0100100101110000",
33984 => "0100100101110000",
33985 => "0100100101110000",
33986 => "0100100101110000",
33987 => "0100100101110000",
33988 => "0100100101110000",
33989 => "0100100110000000",
33990 => "0100100110000000",
33991 => "0100100110000000",
33992 => "0100100110000000",
33993 => "0100100110000000",
33994 => "0100100110000000",
33995 => "0100100110000000",
33996 => "0100100110000000",
33997 => "0100100110010000",
33998 => "0100100110010000",
33999 => "0100100110010000",
34000 => "0100100110010000",
34001 => "0100100110010000",
34002 => "0100100110010000",
34003 => "0100100110010000",
34004 => "0100100110010000",
34005 => "0100100110100000",
34006 => "0100100110100000",
34007 => "0100100110100000",
34008 => "0100100110100000",
34009 => "0100100110100000",
34010 => "0100100110100000",
34011 => "0100100110100000",
34012 => "0100100110100000",
34013 => "0100100110110000",
34014 => "0100100110110000",
34015 => "0100100110110000",
34016 => "0100100110110000",
34017 => "0100100110110000",
34018 => "0100100110110000",
34019 => "0100100110110000",
34020 => "0100100110110000",
34021 => "0100100110110000",
34022 => "0100100111000000",
34023 => "0100100111000000",
34024 => "0100100111000000",
34025 => "0100100111000000",
34026 => "0100100111000000",
34027 => "0100100111000000",
34028 => "0100100111000000",
34029 => "0100100111000000",
34030 => "0100100111010000",
34031 => "0100100111010000",
34032 => "0100100111010000",
34033 => "0100100111010000",
34034 => "0100100111010000",
34035 => "0100100111010000",
34036 => "0100100111010000",
34037 => "0100100111010000",
34038 => "0100100111100000",
34039 => "0100100111100000",
34040 => "0100100111100000",
34041 => "0100100111100000",
34042 => "0100100111100000",
34043 => "0100100111100000",
34044 => "0100100111100000",
34045 => "0100100111100000",
34046 => "0100100111110000",
34047 => "0100100111110000",
34048 => "0100100111110000",
34049 => "0100100111110000",
34050 => "0100100111110000",
34051 => "0100100111110000",
34052 => "0100100111110000",
34053 => "0100100111110000",
34054 => "0100101000000000",
34055 => "0100101000000000",
34056 => "0100101000000000",
34057 => "0100101000000000",
34058 => "0100101000000000",
34059 => "0100101000000000",
34060 => "0100101000000000",
34061 => "0100101000000000",
34062 => "0100101000000000",
34063 => "0100101000010000",
34064 => "0100101000010000",
34065 => "0100101000010000",
34066 => "0100101000010000",
34067 => "0100101000010000",
34068 => "0100101000010000",
34069 => "0100101000010000",
34070 => "0100101000010000",
34071 => "0100101000100000",
34072 => "0100101000100000",
34073 => "0100101000100000",
34074 => "0100101000100000",
34075 => "0100101000100000",
34076 => "0100101000100000",
34077 => "0100101000100000",
34078 => "0100101000100000",
34079 => "0100101000110000",
34080 => "0100101000110000",
34081 => "0100101000110000",
34082 => "0100101000110000",
34083 => "0100101000110000",
34084 => "0100101000110000",
34085 => "0100101000110000",
34086 => "0100101000110000",
34087 => "0100101001000000",
34088 => "0100101001000000",
34089 => "0100101001000000",
34090 => "0100101001000000",
34091 => "0100101001000000",
34092 => "0100101001000000",
34093 => "0100101001000000",
34094 => "0100101001000000",
34095 => "0100101001010000",
34096 => "0100101001010000",
34097 => "0100101001010000",
34098 => "0100101001010000",
34099 => "0100101001010000",
34100 => "0100101001010000",
34101 => "0100101001010000",
34102 => "0100101001010000",
34103 => "0100101001010000",
34104 => "0100101001100000",
34105 => "0100101001100000",
34106 => "0100101001100000",
34107 => "0100101001100000",
34108 => "0100101001100000",
34109 => "0100101001100000",
34110 => "0100101001100000",
34111 => "0100101001100000",
34112 => "0100101001110000",
34113 => "0100101001110000",
34114 => "0100101001110000",
34115 => "0100101001110000",
34116 => "0100101001110000",
34117 => "0100101001110000",
34118 => "0100101001110000",
34119 => "0100101001110000",
34120 => "0100101010000000",
34121 => "0100101010000000",
34122 => "0100101010000000",
34123 => "0100101010000000",
34124 => "0100101010000000",
34125 => "0100101010000000",
34126 => "0100101010000000",
34127 => "0100101010000000",
34128 => "0100101010010000",
34129 => "0100101010010000",
34130 => "0100101010010000",
34131 => "0100101010010000",
34132 => "0100101010010000",
34133 => "0100101010010000",
34134 => "0100101010010000",
34135 => "0100101010010000",
34136 => "0100101010010000",
34137 => "0100101010100000",
34138 => "0100101010100000",
34139 => "0100101010100000",
34140 => "0100101010100000",
34141 => "0100101010100000",
34142 => "0100101010100000",
34143 => "0100101010100000",
34144 => "0100101010100000",
34145 => "0100101010110000",
34146 => "0100101010110000",
34147 => "0100101010110000",
34148 => "0100101010110000",
34149 => "0100101010110000",
34150 => "0100101010110000",
34151 => "0100101010110000",
34152 => "0100101010110000",
34153 => "0100101011000000",
34154 => "0100101011000000",
34155 => "0100101011000000",
34156 => "0100101011000000",
34157 => "0100101011000000",
34158 => "0100101011000000",
34159 => "0100101011000000",
34160 => "0100101011000000",
34161 => "0100101011010000",
34162 => "0100101011010000",
34163 => "0100101011010000",
34164 => "0100101011010000",
34165 => "0100101011010000",
34166 => "0100101011010000",
34167 => "0100101011010000",
34168 => "0100101011010000",
34169 => "0100101011100000",
34170 => "0100101011100000",
34171 => "0100101011100000",
34172 => "0100101011100000",
34173 => "0100101011100000",
34174 => "0100101011100000",
34175 => "0100101011100000",
34176 => "0100101011100000",
34177 => "0100101011100000",
34178 => "0100101011110000",
34179 => "0100101011110000",
34180 => "0100101011110000",
34181 => "0100101011110000",
34182 => "0100101011110000",
34183 => "0100101011110000",
34184 => "0100101011110000",
34185 => "0100101011110000",
34186 => "0100101100000000",
34187 => "0100101100000000",
34188 => "0100101100000000",
34189 => "0100101100000000",
34190 => "0100101100000000",
34191 => "0100101100000000",
34192 => "0100101100000000",
34193 => "0100101100000000",
34194 => "0100101100010000",
34195 => "0100101100010000",
34196 => "0100101100010000",
34197 => "0100101100010000",
34198 => "0100101100010000",
34199 => "0100101100010000",
34200 => "0100101100010000",
34201 => "0100101100010000",
34202 => "0100101100100000",
34203 => "0100101100100000",
34204 => "0100101100100000",
34205 => "0100101100100000",
34206 => "0100101100100000",
34207 => "0100101100100000",
34208 => "0100101100100000",
34209 => "0100101100100000",
34210 => "0100101100100000",
34211 => "0100101100110000",
34212 => "0100101100110000",
34213 => "0100101100110000",
34214 => "0100101100110000",
34215 => "0100101100110000",
34216 => "0100101100110000",
34217 => "0100101100110000",
34218 => "0100101100110000",
34219 => "0100101101000000",
34220 => "0100101101000000",
34221 => "0100101101000000",
34222 => "0100101101000000",
34223 => "0100101101000000",
34224 => "0100101101000000",
34225 => "0100101101000000",
34226 => "0100101101000000",
34227 => "0100101101010000",
34228 => "0100101101010000",
34229 => "0100101101010000",
34230 => "0100101101010000",
34231 => "0100101101010000",
34232 => "0100101101010000",
34233 => "0100101101010000",
34234 => "0100101101010000",
34235 => "0100101101100000",
34236 => "0100101101100000",
34237 => "0100101101100000",
34238 => "0100101101100000",
34239 => "0100101101100000",
34240 => "0100101101100000",
34241 => "0100101101100000",
34242 => "0100101101100000",
34243 => "0100101101100000",
34244 => "0100101101110000",
34245 => "0100101101110000",
34246 => "0100101101110000",
34247 => "0100101101110000",
34248 => "0100101101110000",
34249 => "0100101101110000",
34250 => "0100101101110000",
34251 => "0100101101110000",
34252 => "0100101110000000",
34253 => "0100101110000000",
34254 => "0100101110000000",
34255 => "0100101110000000",
34256 => "0100101110000000",
34257 => "0100101110000000",
34258 => "0100101110000000",
34259 => "0100101110000000",
34260 => "0100101110010000",
34261 => "0100101110010000",
34262 => "0100101110010000",
34263 => "0100101110010000",
34264 => "0100101110010000",
34265 => "0100101110010000",
34266 => "0100101110010000",
34267 => "0100101110010000",
34268 => "0100101110010000",
34269 => "0100101110100000",
34270 => "0100101110100000",
34271 => "0100101110100000",
34272 => "0100101110100000",
34273 => "0100101110100000",
34274 => "0100101110100000",
34275 => "0100101110100000",
34276 => "0100101110100000",
34277 => "0100101110110000",
34278 => "0100101110110000",
34279 => "0100101110110000",
34280 => "0100101110110000",
34281 => "0100101110110000",
34282 => "0100101110110000",
34283 => "0100101110110000",
34284 => "0100101110110000",
34285 => "0100101111000000",
34286 => "0100101111000000",
34287 => "0100101111000000",
34288 => "0100101111000000",
34289 => "0100101111000000",
34290 => "0100101111000000",
34291 => "0100101111000000",
34292 => "0100101111000000",
34293 => "0100101111010000",
34294 => "0100101111010000",
34295 => "0100101111010000",
34296 => "0100101111010000",
34297 => "0100101111010000",
34298 => "0100101111010000",
34299 => "0100101111010000",
34300 => "0100101111010000",
34301 => "0100101111010000",
34302 => "0100101111100000",
34303 => "0100101111100000",
34304 => "0100101111100000",
34305 => "0100101111100000",
34306 => "0100101111100000",
34307 => "0100101111100000",
34308 => "0100101111100000",
34309 => "0100101111100000",
34310 => "0100101111110000",
34311 => "0100101111110000",
34312 => "0100101111110000",
34313 => "0100101111110000",
34314 => "0100101111110000",
34315 => "0100101111110000",
34316 => "0100101111110000",
34317 => "0100101111110000",
34318 => "0100110000000000",
34319 => "0100110000000000",
34320 => "0100110000000000",
34321 => "0100110000000000",
34322 => "0100110000000000",
34323 => "0100110000000000",
34324 => "0100110000000000",
34325 => "0100110000000000",
34326 => "0100110000000000",
34327 => "0100110000010000",
34328 => "0100110000010000",
34329 => "0100110000010000",
34330 => "0100110000010000",
34331 => "0100110000010000",
34332 => "0100110000010000",
34333 => "0100110000010000",
34334 => "0100110000010000",
34335 => "0100110000100000",
34336 => "0100110000100000",
34337 => "0100110000100000",
34338 => "0100110000100000",
34339 => "0100110000100000",
34340 => "0100110000100000",
34341 => "0100110000100000",
34342 => "0100110000100000",
34343 => "0100110000110000",
34344 => "0100110000110000",
34345 => "0100110000110000",
34346 => "0100110000110000",
34347 => "0100110000110000",
34348 => "0100110000110000",
34349 => "0100110000110000",
34350 => "0100110000110000",
34351 => "0100110001000000",
34352 => "0100110001000000",
34353 => "0100110001000000",
34354 => "0100110001000000",
34355 => "0100110001000000",
34356 => "0100110001000000",
34357 => "0100110001000000",
34358 => "0100110001000000",
34359 => "0100110001000000",
34360 => "0100110001010000",
34361 => "0100110001010000",
34362 => "0100110001010000",
34363 => "0100110001010000",
34364 => "0100110001010000",
34365 => "0100110001010000",
34366 => "0100110001010000",
34367 => "0100110001010000",
34368 => "0100110001100000",
34369 => "0100110001100000",
34370 => "0100110001100000",
34371 => "0100110001100000",
34372 => "0100110001100000",
34373 => "0100110001100000",
34374 => "0100110001100000",
34375 => "0100110001100000",
34376 => "0100110001110000",
34377 => "0100110001110000",
34378 => "0100110001110000",
34379 => "0100110001110000",
34380 => "0100110001110000",
34381 => "0100110001110000",
34382 => "0100110001110000",
34383 => "0100110001110000",
34384 => "0100110001110000",
34385 => "0100110010000000",
34386 => "0100110010000000",
34387 => "0100110010000000",
34388 => "0100110010000000",
34389 => "0100110010000000",
34390 => "0100110010000000",
34391 => "0100110010000000",
34392 => "0100110010000000",
34393 => "0100110010010000",
34394 => "0100110010010000",
34395 => "0100110010010000",
34396 => "0100110010010000",
34397 => "0100110010010000",
34398 => "0100110010010000",
34399 => "0100110010010000",
34400 => "0100110010010000",
34401 => "0100110010100000",
34402 => "0100110010100000",
34403 => "0100110010100000",
34404 => "0100110010100000",
34405 => "0100110010100000",
34406 => "0100110010100000",
34407 => "0100110010100000",
34408 => "0100110010100000",
34409 => "0100110010100000",
34410 => "0100110010110000",
34411 => "0100110010110000",
34412 => "0100110010110000",
34413 => "0100110010110000",
34414 => "0100110010110000",
34415 => "0100110010110000",
34416 => "0100110010110000",
34417 => "0100110010110000",
34418 => "0100110011000000",
34419 => "0100110011000000",
34420 => "0100110011000000",
34421 => "0100110011000000",
34422 => "0100110011000000",
34423 => "0100110011000000",
34424 => "0100110011000000",
34425 => "0100110011000000",
34426 => "0100110011010000",
34427 => "0100110011010000",
34428 => "0100110011010000",
34429 => "0100110011010000",
34430 => "0100110011010000",
34431 => "0100110011010000",
34432 => "0100110011010000",
34433 => "0100110011010000",
34434 => "0100110011010000",
34435 => "0100110011100000",
34436 => "0100110011100000",
34437 => "0100110011100000",
34438 => "0100110011100000",
34439 => "0100110011100000",
34440 => "0100110011100000",
34441 => "0100110011100000",
34442 => "0100110011100000",
34443 => "0100110011110000",
34444 => "0100110011110000",
34445 => "0100110011110000",
34446 => "0100110011110000",
34447 => "0100110011110000",
34448 => "0100110011110000",
34449 => "0100110011110000",
34450 => "0100110011110000",
34451 => "0100110100000000",
34452 => "0100110100000000",
34453 => "0100110100000000",
34454 => "0100110100000000",
34455 => "0100110100000000",
34456 => "0100110100000000",
34457 => "0100110100000000",
34458 => "0100110100000000",
34459 => "0100110100000000",
34460 => "0100110100010000",
34461 => "0100110100010000",
34462 => "0100110100010000",
34463 => "0100110100010000",
34464 => "0100110100010000",
34465 => "0100110100010000",
34466 => "0100110100010000",
34467 => "0100110100010000",
34468 => "0100110100100000",
34469 => "0100110100100000",
34470 => "0100110100100000",
34471 => "0100110100100000",
34472 => "0100110100100000",
34473 => "0100110100100000",
34474 => "0100110100100000",
34475 => "0100110100100000",
34476 => "0100110100110000",
34477 => "0100110100110000",
34478 => "0100110100110000",
34479 => "0100110100110000",
34480 => "0100110100110000",
34481 => "0100110100110000",
34482 => "0100110100110000",
34483 => "0100110100110000",
34484 => "0100110100110000",
34485 => "0100110101000000",
34486 => "0100110101000000",
34487 => "0100110101000000",
34488 => "0100110101000000",
34489 => "0100110101000000",
34490 => "0100110101000000",
34491 => "0100110101000000",
34492 => "0100110101000000",
34493 => "0100110101010000",
34494 => "0100110101010000",
34495 => "0100110101010000",
34496 => "0100110101010000",
34497 => "0100110101010000",
34498 => "0100110101010000",
34499 => "0100110101010000",
34500 => "0100110101010000",
34501 => "0100110101100000",
34502 => "0100110101100000",
34503 => "0100110101100000",
34504 => "0100110101100000",
34505 => "0100110101100000",
34506 => "0100110101100000",
34507 => "0100110101100000",
34508 => "0100110101100000",
34509 => "0100110101100000",
34510 => "0100110101110000",
34511 => "0100110101110000",
34512 => "0100110101110000",
34513 => "0100110101110000",
34514 => "0100110101110000",
34515 => "0100110101110000",
34516 => "0100110101110000",
34517 => "0100110101110000",
34518 => "0100110110000000",
34519 => "0100110110000000",
34520 => "0100110110000000",
34521 => "0100110110000000",
34522 => "0100110110000000",
34523 => "0100110110000000",
34524 => "0100110110000000",
34525 => "0100110110000000",
34526 => "0100110110010000",
34527 => "0100110110010000",
34528 => "0100110110010000",
34529 => "0100110110010000",
34530 => "0100110110010000",
34531 => "0100110110010000",
34532 => "0100110110010000",
34533 => "0100110110010000",
34534 => "0100110110010000",
34535 => "0100110110100000",
34536 => "0100110110100000",
34537 => "0100110110100000",
34538 => "0100110110100000",
34539 => "0100110110100000",
34540 => "0100110110100000",
34541 => "0100110110100000",
34542 => "0100110110100000",
34543 => "0100110110110000",
34544 => "0100110110110000",
34545 => "0100110110110000",
34546 => "0100110110110000",
34547 => "0100110110110000",
34548 => "0100110110110000",
34549 => "0100110110110000",
34550 => "0100110110110000",
34551 => "0100110110110000",
34552 => "0100110111000000",
34553 => "0100110111000000",
34554 => "0100110111000000",
34555 => "0100110111000000",
34556 => "0100110111000000",
34557 => "0100110111000000",
34558 => "0100110111000000",
34559 => "0100110111000000",
34560 => "0100110111010000",
34561 => "0100110111010000",
34562 => "0100110111010000",
34563 => "0100110111010000",
34564 => "0100110111010000",
34565 => "0100110111010000",
34566 => "0100110111010000",
34567 => "0100110111010000",
34568 => "0100110111100000",
34569 => "0100110111100000",
34570 => "0100110111100000",
34571 => "0100110111100000",
34572 => "0100110111100000",
34573 => "0100110111100000",
34574 => "0100110111100000",
34575 => "0100110111100000",
34576 => "0100110111100000",
34577 => "0100110111110000",
34578 => "0100110111110000",
34579 => "0100110111110000",
34580 => "0100110111110000",
34581 => "0100110111110000",
34582 => "0100110111110000",
34583 => "0100110111110000",
34584 => "0100110111110000",
34585 => "0100111000000000",
34586 => "0100111000000000",
34587 => "0100111000000000",
34588 => "0100111000000000",
34589 => "0100111000000000",
34590 => "0100111000000000",
34591 => "0100111000000000",
34592 => "0100111000000000",
34593 => "0100111000000000",
34594 => "0100111000010000",
34595 => "0100111000010000",
34596 => "0100111000010000",
34597 => "0100111000010000",
34598 => "0100111000010000",
34599 => "0100111000010000",
34600 => "0100111000010000",
34601 => "0100111000010000",
34602 => "0100111000100000",
34603 => "0100111000100000",
34604 => "0100111000100000",
34605 => "0100111000100000",
34606 => "0100111000100000",
34607 => "0100111000100000",
34608 => "0100111000100000",
34609 => "0100111000100000",
34610 => "0100111000110000",
34611 => "0100111000110000",
34612 => "0100111000110000",
34613 => "0100111000110000",
34614 => "0100111000110000",
34615 => "0100111000110000",
34616 => "0100111000110000",
34617 => "0100111000110000",
34618 => "0100111000110000",
34619 => "0100111001000000",
34620 => "0100111001000000",
34621 => "0100111001000000",
34622 => "0100111001000000",
34623 => "0100111001000000",
34624 => "0100111001000000",
34625 => "0100111001000000",
34626 => "0100111001000000",
34627 => "0100111001010000",
34628 => "0100111001010000",
34629 => "0100111001010000",
34630 => "0100111001010000",
34631 => "0100111001010000",
34632 => "0100111001010000",
34633 => "0100111001010000",
34634 => "0100111001010000",
34635 => "0100111001010000",
34636 => "0100111001100000",
34637 => "0100111001100000",
34638 => "0100111001100000",
34639 => "0100111001100000",
34640 => "0100111001100000",
34641 => "0100111001100000",
34642 => "0100111001100000",
34643 => "0100111001100000",
34644 => "0100111001110000",
34645 => "0100111001110000",
34646 => "0100111001110000",
34647 => "0100111001110000",
34648 => "0100111001110000",
34649 => "0100111001110000",
34650 => "0100111001110000",
34651 => "0100111001110000",
34652 => "0100111001110000",
34653 => "0100111010000000",
34654 => "0100111010000000",
34655 => "0100111010000000",
34656 => "0100111010000000",
34657 => "0100111010000000",
34658 => "0100111010000000",
34659 => "0100111010000000",
34660 => "0100111010000000",
34661 => "0100111010010000",
34662 => "0100111010010000",
34663 => "0100111010010000",
34664 => "0100111010010000",
34665 => "0100111010010000",
34666 => "0100111010010000",
34667 => "0100111010010000",
34668 => "0100111010010000",
34669 => "0100111010100000",
34670 => "0100111010100000",
34671 => "0100111010100000",
34672 => "0100111010100000",
34673 => "0100111010100000",
34674 => "0100111010100000",
34675 => "0100111010100000",
34676 => "0100111010100000",
34677 => "0100111010100000",
34678 => "0100111010110000",
34679 => "0100111010110000",
34680 => "0100111010110000",
34681 => "0100111010110000",
34682 => "0100111010110000",
34683 => "0100111010110000",
34684 => "0100111010110000",
34685 => "0100111010110000",
34686 => "0100111011000000",
34687 => "0100111011000000",
34688 => "0100111011000000",
34689 => "0100111011000000",
34690 => "0100111011000000",
34691 => "0100111011000000",
34692 => "0100111011000000",
34693 => "0100111011000000",
34694 => "0100111011000000",
34695 => "0100111011010000",
34696 => "0100111011010000",
34697 => "0100111011010000",
34698 => "0100111011010000",
34699 => "0100111011010000",
34700 => "0100111011010000",
34701 => "0100111011010000",
34702 => "0100111011010000",
34703 => "0100111011100000",
34704 => "0100111011100000",
34705 => "0100111011100000",
34706 => "0100111011100000",
34707 => "0100111011100000",
34708 => "0100111011100000",
34709 => "0100111011100000",
34710 => "0100111011100000",
34711 => "0100111011100000",
34712 => "0100111011110000",
34713 => "0100111011110000",
34714 => "0100111011110000",
34715 => "0100111011110000",
34716 => "0100111011110000",
34717 => "0100111011110000",
34718 => "0100111011110000",
34719 => "0100111011110000",
34720 => "0100111100000000",
34721 => "0100111100000000",
34722 => "0100111100000000",
34723 => "0100111100000000",
34724 => "0100111100000000",
34725 => "0100111100000000",
34726 => "0100111100000000",
34727 => "0100111100000000",
34728 => "0100111100000000",
34729 => "0100111100010000",
34730 => "0100111100010000",
34731 => "0100111100010000",
34732 => "0100111100010000",
34733 => "0100111100010000",
34734 => "0100111100010000",
34735 => "0100111100010000",
34736 => "0100111100010000",
34737 => "0100111100100000",
34738 => "0100111100100000",
34739 => "0100111100100000",
34740 => "0100111100100000",
34741 => "0100111100100000",
34742 => "0100111100100000",
34743 => "0100111100100000",
34744 => "0100111100100000",
34745 => "0100111100100000",
34746 => "0100111100110000",
34747 => "0100111100110000",
34748 => "0100111100110000",
34749 => "0100111100110000",
34750 => "0100111100110000",
34751 => "0100111100110000",
34752 => "0100111100110000",
34753 => "0100111100110000",
34754 => "0100111101000000",
34755 => "0100111101000000",
34756 => "0100111101000000",
34757 => "0100111101000000",
34758 => "0100111101000000",
34759 => "0100111101000000",
34760 => "0100111101000000",
34761 => "0100111101000000",
34762 => "0100111101010000",
34763 => "0100111101010000",
34764 => "0100111101010000",
34765 => "0100111101010000",
34766 => "0100111101010000",
34767 => "0100111101010000",
34768 => "0100111101010000",
34769 => "0100111101010000",
34770 => "0100111101010000",
34771 => "0100111101100000",
34772 => "0100111101100000",
34773 => "0100111101100000",
34774 => "0100111101100000",
34775 => "0100111101100000",
34776 => "0100111101100000",
34777 => "0100111101100000",
34778 => "0100111101100000",
34779 => "0100111101110000",
34780 => "0100111101110000",
34781 => "0100111101110000",
34782 => "0100111101110000",
34783 => "0100111101110000",
34784 => "0100111101110000",
34785 => "0100111101110000",
34786 => "0100111101110000",
34787 => "0100111101110000",
34788 => "0100111110000000",
34789 => "0100111110000000",
34790 => "0100111110000000",
34791 => "0100111110000000",
34792 => "0100111110000000",
34793 => "0100111110000000",
34794 => "0100111110000000",
34795 => "0100111110000000",
34796 => "0100111110010000",
34797 => "0100111110010000",
34798 => "0100111110010000",
34799 => "0100111110010000",
34800 => "0100111110010000",
34801 => "0100111110010000",
34802 => "0100111110010000",
34803 => "0100111110010000",
34804 => "0100111110010000",
34805 => "0100111110100000",
34806 => "0100111110100000",
34807 => "0100111110100000",
34808 => "0100111110100000",
34809 => "0100111110100000",
34810 => "0100111110100000",
34811 => "0100111110100000",
34812 => "0100111110100000",
34813 => "0100111110110000",
34814 => "0100111110110000",
34815 => "0100111110110000",
34816 => "0100111110110000",
34817 => "0100111110110000",
34818 => "0100111110110000",
34819 => "0100111110110000",
34820 => "0100111110110000",
34821 => "0100111110110000",
34822 => "0100111111000000",
34823 => "0100111111000000",
34824 => "0100111111000000",
34825 => "0100111111000000",
34826 => "0100111111000000",
34827 => "0100111111000000",
34828 => "0100111111000000",
34829 => "0100111111000000",
34830 => "0100111111010000",
34831 => "0100111111010000",
34832 => "0100111111010000",
34833 => "0100111111010000",
34834 => "0100111111010000",
34835 => "0100111111010000",
34836 => "0100111111010000",
34837 => "0100111111010000",
34838 => "0100111111010000",
34839 => "0100111111100000",
34840 => "0100111111100000",
34841 => "0100111111100000",
34842 => "0100111111100000",
34843 => "0100111111100000",
34844 => "0100111111100000",
34845 => "0100111111100000",
34846 => "0100111111100000",
34847 => "0100111111100000",
34848 => "0100111111110000",
34849 => "0100111111110000",
34850 => "0100111111110000",
34851 => "0100111111110000",
34852 => "0100111111110000",
34853 => "0100111111110000",
34854 => "0100111111110000",
34855 => "0100111111110000",
34856 => "0101000000000000",
34857 => "0101000000000000",
34858 => "0101000000000000",
34859 => "0101000000000000",
34860 => "0101000000000000",
34861 => "0101000000000000",
34862 => "0101000000000000",
34863 => "0101000000000000",
34864 => "0101000000000000",
34865 => "0101000000010000",
34866 => "0101000000010000",
34867 => "0101000000010000",
34868 => "0101000000010000",
34869 => "0101000000010000",
34870 => "0101000000010000",
34871 => "0101000000010000",
34872 => "0101000000010000",
34873 => "0101000000100000",
34874 => "0101000000100000",
34875 => "0101000000100000",
34876 => "0101000000100000",
34877 => "0101000000100000",
34878 => "0101000000100000",
34879 => "0101000000100000",
34880 => "0101000000100000",
34881 => "0101000000100000",
34882 => "0101000000110000",
34883 => "0101000000110000",
34884 => "0101000000110000",
34885 => "0101000000110000",
34886 => "0101000000110000",
34887 => "0101000000110000",
34888 => "0101000000110000",
34889 => "0101000000110000",
34890 => "0101000001000000",
34891 => "0101000001000000",
34892 => "0101000001000000",
34893 => "0101000001000000",
34894 => "0101000001000000",
34895 => "0101000001000000",
34896 => "0101000001000000",
34897 => "0101000001000000",
34898 => "0101000001000000",
34899 => "0101000001010000",
34900 => "0101000001010000",
34901 => "0101000001010000",
34902 => "0101000001010000",
34903 => "0101000001010000",
34904 => "0101000001010000",
34905 => "0101000001010000",
34906 => "0101000001010000",
34907 => "0101000001100000",
34908 => "0101000001100000",
34909 => "0101000001100000",
34910 => "0101000001100000",
34911 => "0101000001100000",
34912 => "0101000001100000",
34913 => "0101000001100000",
34914 => "0101000001100000",
34915 => "0101000001100000",
34916 => "0101000001110000",
34917 => "0101000001110000",
34918 => "0101000001110000",
34919 => "0101000001110000",
34920 => "0101000001110000",
34921 => "0101000001110000",
34922 => "0101000001110000",
34923 => "0101000001110000",
34924 => "0101000010000000",
34925 => "0101000010000000",
34926 => "0101000010000000",
34927 => "0101000010000000",
34928 => "0101000010000000",
34929 => "0101000010000000",
34930 => "0101000010000000",
34931 => "0101000010000000",
34932 => "0101000010000000",
34933 => "0101000010010000",
34934 => "0101000010010000",
34935 => "0101000010010000",
34936 => "0101000010010000",
34937 => "0101000010010000",
34938 => "0101000010010000",
34939 => "0101000010010000",
34940 => "0101000010010000",
34941 => "0101000010010000",
34942 => "0101000010100000",
34943 => "0101000010100000",
34944 => "0101000010100000",
34945 => "0101000010100000",
34946 => "0101000010100000",
34947 => "0101000010100000",
34948 => "0101000010100000",
34949 => "0101000010100000",
34950 => "0101000010110000",
34951 => "0101000010110000",
34952 => "0101000010110000",
34953 => "0101000010110000",
34954 => "0101000010110000",
34955 => "0101000010110000",
34956 => "0101000010110000",
34957 => "0101000010110000",
34958 => "0101000010110000",
34959 => "0101000011000000",
34960 => "0101000011000000",
34961 => "0101000011000000",
34962 => "0101000011000000",
34963 => "0101000011000000",
34964 => "0101000011000000",
34965 => "0101000011000000",
34966 => "0101000011000000",
34967 => "0101000011010000",
34968 => "0101000011010000",
34969 => "0101000011010000",
34970 => "0101000011010000",
34971 => "0101000011010000",
34972 => "0101000011010000",
34973 => "0101000011010000",
34974 => "0101000011010000",
34975 => "0101000011010000",
34976 => "0101000011100000",
34977 => "0101000011100000",
34978 => "0101000011100000",
34979 => "0101000011100000",
34980 => "0101000011100000",
34981 => "0101000011100000",
34982 => "0101000011100000",
34983 => "0101000011100000",
34984 => "0101000011100000",
34985 => "0101000011110000",
34986 => "0101000011110000",
34987 => "0101000011110000",
34988 => "0101000011110000",
34989 => "0101000011110000",
34990 => "0101000011110000",
34991 => "0101000011110000",
34992 => "0101000011110000",
34993 => "0101000100000000",
34994 => "0101000100000000",
34995 => "0101000100000000",
34996 => "0101000100000000",
34997 => "0101000100000000",
34998 => "0101000100000000",
34999 => "0101000100000000",
35000 => "0101000100000000",
35001 => "0101000100000000",
35002 => "0101000100010000",
35003 => "0101000100010000",
35004 => "0101000100010000",
35005 => "0101000100010000",
35006 => "0101000100010000",
35007 => "0101000100010000",
35008 => "0101000100010000",
35009 => "0101000100010000",
35010 => "0101000100100000",
35011 => "0101000100100000",
35012 => "0101000100100000",
35013 => "0101000100100000",
35014 => "0101000100100000",
35015 => "0101000100100000",
35016 => "0101000100100000",
35017 => "0101000100100000",
35018 => "0101000100100000",
35019 => "0101000100110000",
35020 => "0101000100110000",
35021 => "0101000100110000",
35022 => "0101000100110000",
35023 => "0101000100110000",
35024 => "0101000100110000",
35025 => "0101000100110000",
35026 => "0101000100110000",
35027 => "0101000100110000",
35028 => "0101000101000000",
35029 => "0101000101000000",
35030 => "0101000101000000",
35031 => "0101000101000000",
35032 => "0101000101000000",
35033 => "0101000101000000",
35034 => "0101000101000000",
35035 => "0101000101000000",
35036 => "0101000101010000",
35037 => "0101000101010000",
35038 => "0101000101010000",
35039 => "0101000101010000",
35040 => "0101000101010000",
35041 => "0101000101010000",
35042 => "0101000101010000",
35043 => "0101000101010000",
35044 => "0101000101010000",
35045 => "0101000101100000",
35046 => "0101000101100000",
35047 => "0101000101100000",
35048 => "0101000101100000",
35049 => "0101000101100000",
35050 => "0101000101100000",
35051 => "0101000101100000",
35052 => "0101000101100000",
35053 => "0101000101110000",
35054 => "0101000101110000",
35055 => "0101000101110000",
35056 => "0101000101110000",
35057 => "0101000101110000",
35058 => "0101000101110000",
35059 => "0101000101110000",
35060 => "0101000101110000",
35061 => "0101000101110000",
35062 => "0101000110000000",
35063 => "0101000110000000",
35064 => "0101000110000000",
35065 => "0101000110000000",
35066 => "0101000110000000",
35067 => "0101000110000000",
35068 => "0101000110000000",
35069 => "0101000110000000",
35070 => "0101000110000000",
35071 => "0101000110010000",
35072 => "0101000110010000",
35073 => "0101000110010000",
35074 => "0101000110010000",
35075 => "0101000110010000",
35076 => "0101000110010000",
35077 => "0101000110010000",
35078 => "0101000110010000",
35079 => "0101000110100000",
35080 => "0101000110100000",
35081 => "0101000110100000",
35082 => "0101000110100000",
35083 => "0101000110100000",
35084 => "0101000110100000",
35085 => "0101000110100000",
35086 => "0101000110100000",
35087 => "0101000110100000",
35088 => "0101000110110000",
35089 => "0101000110110000",
35090 => "0101000110110000",
35091 => "0101000110110000",
35092 => "0101000110110000",
35093 => "0101000110110000",
35094 => "0101000110110000",
35095 => "0101000110110000",
35096 => "0101000110110000",
35097 => "0101000111000000",
35098 => "0101000111000000",
35099 => "0101000111000000",
35100 => "0101000111000000",
35101 => "0101000111000000",
35102 => "0101000111000000",
35103 => "0101000111000000",
35104 => "0101000111000000",
35105 => "0101000111010000",
35106 => "0101000111010000",
35107 => "0101000111010000",
35108 => "0101000111010000",
35109 => "0101000111010000",
35110 => "0101000111010000",
35111 => "0101000111010000",
35112 => "0101000111010000",
35113 => "0101000111010000",
35114 => "0101000111100000",
35115 => "0101000111100000",
35116 => "0101000111100000",
35117 => "0101000111100000",
35118 => "0101000111100000",
35119 => "0101000111100000",
35120 => "0101000111100000",
35121 => "0101000111100000",
35122 => "0101000111100000",
35123 => "0101000111110000",
35124 => "0101000111110000",
35125 => "0101000111110000",
35126 => "0101000111110000",
35127 => "0101000111110000",
35128 => "0101000111110000",
35129 => "0101000111110000",
35130 => "0101000111110000",
35131 => "0101001000000000",
35132 => "0101001000000000",
35133 => "0101001000000000",
35134 => "0101001000000000",
35135 => "0101001000000000",
35136 => "0101001000000000",
35137 => "0101001000000000",
35138 => "0101001000000000",
35139 => "0101001000000000",
35140 => "0101001000010000",
35141 => "0101001000010000",
35142 => "0101001000010000",
35143 => "0101001000010000",
35144 => "0101001000010000",
35145 => "0101001000010000",
35146 => "0101001000010000",
35147 => "0101001000010000",
35148 => "0101001000010000",
35149 => "0101001000100000",
35150 => "0101001000100000",
35151 => "0101001000100000",
35152 => "0101001000100000",
35153 => "0101001000100000",
35154 => "0101001000100000",
35155 => "0101001000100000",
35156 => "0101001000100000",
35157 => "0101001000100000",
35158 => "0101001000110000",
35159 => "0101001000110000",
35160 => "0101001000110000",
35161 => "0101001000110000",
35162 => "0101001000110000",
35163 => "0101001000110000",
35164 => "0101001000110000",
35165 => "0101001000110000",
35166 => "0101001001000000",
35167 => "0101001001000000",
35168 => "0101001001000000",
35169 => "0101001001000000",
35170 => "0101001001000000",
35171 => "0101001001000000",
35172 => "0101001001000000",
35173 => "0101001001000000",
35174 => "0101001001000000",
35175 => "0101001001010000",
35176 => "0101001001010000",
35177 => "0101001001010000",
35178 => "0101001001010000",
35179 => "0101001001010000",
35180 => "0101001001010000",
35181 => "0101001001010000",
35182 => "0101001001010000",
35183 => "0101001001010000",
35184 => "0101001001100000",
35185 => "0101001001100000",
35186 => "0101001001100000",
35187 => "0101001001100000",
35188 => "0101001001100000",
35189 => "0101001001100000",
35190 => "0101001001100000",
35191 => "0101001001100000",
35192 => "0101001001110000",
35193 => "0101001001110000",
35194 => "0101001001110000",
35195 => "0101001001110000",
35196 => "0101001001110000",
35197 => "0101001001110000",
35198 => "0101001001110000",
35199 => "0101001001110000",
35200 => "0101001001110000",
35201 => "0101001010000000",
35202 => "0101001010000000",
35203 => "0101001010000000",
35204 => "0101001010000000",
35205 => "0101001010000000",
35206 => "0101001010000000",
35207 => "0101001010000000",
35208 => "0101001010000000",
35209 => "0101001010000000",
35210 => "0101001010010000",
35211 => "0101001010010000",
35212 => "0101001010010000",
35213 => "0101001010010000",
35214 => "0101001010010000",
35215 => "0101001010010000",
35216 => "0101001010010000",
35217 => "0101001010010000",
35218 => "0101001010010000",
35219 => "0101001010100000",
35220 => "0101001010100000",
35221 => "0101001010100000",
35222 => "0101001010100000",
35223 => "0101001010100000",
35224 => "0101001010100000",
35225 => "0101001010100000",
35226 => "0101001010100000",
35227 => "0101001010110000",
35228 => "0101001010110000",
35229 => "0101001010110000",
35230 => "0101001010110000",
35231 => "0101001010110000",
35232 => "0101001010110000",
35233 => "0101001010110000",
35234 => "0101001010110000",
35235 => "0101001010110000",
35236 => "0101001011000000",
35237 => "0101001011000000",
35238 => "0101001011000000",
35239 => "0101001011000000",
35240 => "0101001011000000",
35241 => "0101001011000000",
35242 => "0101001011000000",
35243 => "0101001011000000",
35244 => "0101001011000000",
35245 => "0101001011010000",
35246 => "0101001011010000",
35247 => "0101001011010000",
35248 => "0101001011010000",
35249 => "0101001011010000",
35250 => "0101001011010000",
35251 => "0101001011010000",
35252 => "0101001011010000",
35253 => "0101001011010000",
35254 => "0101001011100000",
35255 => "0101001011100000",
35256 => "0101001011100000",
35257 => "0101001011100000",
35258 => "0101001011100000",
35259 => "0101001011100000",
35260 => "0101001011100000",
35261 => "0101001011100000",
35262 => "0101001011110000",
35263 => "0101001011110000",
35264 => "0101001011110000",
35265 => "0101001011110000",
35266 => "0101001011110000",
35267 => "0101001011110000",
35268 => "0101001011110000",
35269 => "0101001011110000",
35270 => "0101001011110000",
35271 => "0101001100000000",
35272 => "0101001100000000",
35273 => "0101001100000000",
35274 => "0101001100000000",
35275 => "0101001100000000",
35276 => "0101001100000000",
35277 => "0101001100000000",
35278 => "0101001100000000",
35279 => "0101001100000000",
35280 => "0101001100010000",
35281 => "0101001100010000",
35282 => "0101001100010000",
35283 => "0101001100010000",
35284 => "0101001100010000",
35285 => "0101001100010000",
35286 => "0101001100010000",
35287 => "0101001100010000",
35288 => "0101001100010000",
35289 => "0101001100100000",
35290 => "0101001100100000",
35291 => "0101001100100000",
35292 => "0101001100100000",
35293 => "0101001100100000",
35294 => "0101001100100000",
35295 => "0101001100100000",
35296 => "0101001100100000",
35297 => "0101001100110000",
35298 => "0101001100110000",
35299 => "0101001100110000",
35300 => "0101001100110000",
35301 => "0101001100110000",
35302 => "0101001100110000",
35303 => "0101001100110000",
35304 => "0101001100110000",
35305 => "0101001100110000",
35306 => "0101001101000000",
35307 => "0101001101000000",
35308 => "0101001101000000",
35309 => "0101001101000000",
35310 => "0101001101000000",
35311 => "0101001101000000",
35312 => "0101001101000000",
35313 => "0101001101000000",
35314 => "0101001101000000",
35315 => "0101001101010000",
35316 => "0101001101010000",
35317 => "0101001101010000",
35318 => "0101001101010000",
35319 => "0101001101010000",
35320 => "0101001101010000",
35321 => "0101001101010000",
35322 => "0101001101010000",
35323 => "0101001101010000",
35324 => "0101001101100000",
35325 => "0101001101100000",
35326 => "0101001101100000",
35327 => "0101001101100000",
35328 => "0101001101100000",
35329 => "0101001101100000",
35330 => "0101001101100000",
35331 => "0101001101100000",
35332 => "0101001101100000",
35333 => "0101001101110000",
35334 => "0101001101110000",
35335 => "0101001101110000",
35336 => "0101001101110000",
35337 => "0101001101110000",
35338 => "0101001101110000",
35339 => "0101001101110000",
35340 => "0101001101110000",
35341 => "0101001110000000",
35342 => "0101001110000000",
35343 => "0101001110000000",
35344 => "0101001110000000",
35345 => "0101001110000000",
35346 => "0101001110000000",
35347 => "0101001110000000",
35348 => "0101001110000000",
35349 => "0101001110000000",
35350 => "0101001110010000",
35351 => "0101001110010000",
35352 => "0101001110010000",
35353 => "0101001110010000",
35354 => "0101001110010000",
35355 => "0101001110010000",
35356 => "0101001110010000",
35357 => "0101001110010000",
35358 => "0101001110010000",
35359 => "0101001110100000",
35360 => "0101001110100000",
35361 => "0101001110100000",
35362 => "0101001110100000",
35363 => "0101001110100000",
35364 => "0101001110100000",
35365 => "0101001110100000",
35366 => "0101001110100000",
35367 => "0101001110100000",
35368 => "0101001110110000",
35369 => "0101001110110000",
35370 => "0101001110110000",
35371 => "0101001110110000",
35372 => "0101001110110000",
35373 => "0101001110110000",
35374 => "0101001110110000",
35375 => "0101001110110000",
35376 => "0101001110110000",
35377 => "0101001111000000",
35378 => "0101001111000000",
35379 => "0101001111000000",
35380 => "0101001111000000",
35381 => "0101001111000000",
35382 => "0101001111000000",
35383 => "0101001111000000",
35384 => "0101001111000000",
35385 => "0101001111000000",
35386 => "0101001111010000",
35387 => "0101001111010000",
35388 => "0101001111010000",
35389 => "0101001111010000",
35390 => "0101001111010000",
35391 => "0101001111010000",
35392 => "0101001111010000",
35393 => "0101001111010000",
35394 => "0101001111100000",
35395 => "0101001111100000",
35396 => "0101001111100000",
35397 => "0101001111100000",
35398 => "0101001111100000",
35399 => "0101001111100000",
35400 => "0101001111100000",
35401 => "0101001111100000",
35402 => "0101001111100000",
35403 => "0101001111110000",
35404 => "0101001111110000",
35405 => "0101001111110000",
35406 => "0101001111110000",
35407 => "0101001111110000",
35408 => "0101001111110000",
35409 => "0101001111110000",
35410 => "0101001111110000",
35411 => "0101001111110000",
35412 => "0101010000000000",
35413 => "0101010000000000",
35414 => "0101010000000000",
35415 => "0101010000000000",
35416 => "0101010000000000",
35417 => "0101010000000000",
35418 => "0101010000000000",
35419 => "0101010000000000",
35420 => "0101010000000000",
35421 => "0101010000010000",
35422 => "0101010000010000",
35423 => "0101010000010000",
35424 => "0101010000010000",
35425 => "0101010000010000",
35426 => "0101010000010000",
35427 => "0101010000010000",
35428 => "0101010000010000",
35429 => "0101010000010000",
35430 => "0101010000100000",
35431 => "0101010000100000",
35432 => "0101010000100000",
35433 => "0101010000100000",
35434 => "0101010000100000",
35435 => "0101010000100000",
35436 => "0101010000100000",
35437 => "0101010000100000",
35438 => "0101010000100000",
35439 => "0101010000110000",
35440 => "0101010000110000",
35441 => "0101010000110000",
35442 => "0101010000110000",
35443 => "0101010000110000",
35444 => "0101010000110000",
35445 => "0101010000110000",
35446 => "0101010000110000",
35447 => "0101010000110000",
35448 => "0101010001000000",
35449 => "0101010001000000",
35450 => "0101010001000000",
35451 => "0101010001000000",
35452 => "0101010001000000",
35453 => "0101010001000000",
35454 => "0101010001000000",
35455 => "0101010001000000",
35456 => "0101010001000000",
35457 => "0101010001010000",
35458 => "0101010001010000",
35459 => "0101010001010000",
35460 => "0101010001010000",
35461 => "0101010001010000",
35462 => "0101010001010000",
35463 => "0101010001010000",
35464 => "0101010001010000",
35465 => "0101010001100000",
35466 => "0101010001100000",
35467 => "0101010001100000",
35468 => "0101010001100000",
35469 => "0101010001100000",
35470 => "0101010001100000",
35471 => "0101010001100000",
35472 => "0101010001100000",
35473 => "0101010001100000",
35474 => "0101010001110000",
35475 => "0101010001110000",
35476 => "0101010001110000",
35477 => "0101010001110000",
35478 => "0101010001110000",
35479 => "0101010001110000",
35480 => "0101010001110000",
35481 => "0101010001110000",
35482 => "0101010001110000",
35483 => "0101010010000000",
35484 => "0101010010000000",
35485 => "0101010010000000",
35486 => "0101010010000000",
35487 => "0101010010000000",
35488 => "0101010010000000",
35489 => "0101010010000000",
35490 => "0101010010000000",
35491 => "0101010010000000",
35492 => "0101010010010000",
35493 => "0101010010010000",
35494 => "0101010010010000",
35495 => "0101010010010000",
35496 => "0101010010010000",
35497 => "0101010010010000",
35498 => "0101010010010000",
35499 => "0101010010010000",
35500 => "0101010010010000",
35501 => "0101010010100000",
35502 => "0101010010100000",
35503 => "0101010010100000",
35504 => "0101010010100000",
35505 => "0101010010100000",
35506 => "0101010010100000",
35507 => "0101010010100000",
35508 => "0101010010100000",
35509 => "0101010010100000",
35510 => "0101010010110000",
35511 => "0101010010110000",
35512 => "0101010010110000",
35513 => "0101010010110000",
35514 => "0101010010110000",
35515 => "0101010010110000",
35516 => "0101010010110000",
35517 => "0101010010110000",
35518 => "0101010010110000",
35519 => "0101010011000000",
35520 => "0101010011000000",
35521 => "0101010011000000",
35522 => "0101010011000000",
35523 => "0101010011000000",
35524 => "0101010011000000",
35525 => "0101010011000000",
35526 => "0101010011000000",
35527 => "0101010011000000",
35528 => "0101010011010000",
35529 => "0101010011010000",
35530 => "0101010011010000",
35531 => "0101010011010000",
35532 => "0101010011010000",
35533 => "0101010011010000",
35534 => "0101010011010000",
35535 => "0101010011010000",
35536 => "0101010011010000",
35537 => "0101010011100000",
35538 => "0101010011100000",
35539 => "0101010011100000",
35540 => "0101010011100000",
35541 => "0101010011100000",
35542 => "0101010011100000",
35543 => "0101010011100000",
35544 => "0101010011100000",
35545 => "0101010011100000",
35546 => "0101010011110000",
35547 => "0101010011110000",
35548 => "0101010011110000",
35549 => "0101010011110000",
35550 => "0101010011110000",
35551 => "0101010011110000",
35552 => "0101010011110000",
35553 => "0101010011110000",
35554 => "0101010011110000",
35555 => "0101010100000000",
35556 => "0101010100000000",
35557 => "0101010100000000",
35558 => "0101010100000000",
35559 => "0101010100000000",
35560 => "0101010100000000",
35561 => "0101010100000000",
35562 => "0101010100000000",
35563 => "0101010100000000",
35564 => "0101010100010000",
35565 => "0101010100010000",
35566 => "0101010100010000",
35567 => "0101010100010000",
35568 => "0101010100010000",
35569 => "0101010100010000",
35570 => "0101010100010000",
35571 => "0101010100010000",
35572 => "0101010100010000",
35573 => "0101010100100000",
35574 => "0101010100100000",
35575 => "0101010100100000",
35576 => "0101010100100000",
35577 => "0101010100100000",
35578 => "0101010100100000",
35579 => "0101010100100000",
35580 => "0101010100100000",
35581 => "0101010100100000",
35582 => "0101010100110000",
35583 => "0101010100110000",
35584 => "0101010100110000",
35585 => "0101010100110000",
35586 => "0101010100110000",
35587 => "0101010100110000",
35588 => "0101010100110000",
35589 => "0101010100110000",
35590 => "0101010100110000",
35591 => "0101010101000000",
35592 => "0101010101000000",
35593 => "0101010101000000",
35594 => "0101010101000000",
35595 => "0101010101000000",
35596 => "0101010101000000",
35597 => "0101010101000000",
35598 => "0101010101000000",
35599 => "0101010101000000",
35600 => "0101010101010000",
35601 => "0101010101010000",
35602 => "0101010101010000",
35603 => "0101010101010000",
35604 => "0101010101010000",
35605 => "0101010101010000",
35606 => "0101010101010000",
35607 => "0101010101010000",
35608 => "0101010101010000",
35609 => "0101010101100000",
35610 => "0101010101100000",
35611 => "0101010101100000",
35612 => "0101010101100000",
35613 => "0101010101100000",
35614 => "0101010101100000",
35615 => "0101010101100000",
35616 => "0101010101100000",
35617 => "0101010101100000",
35618 => "0101010101110000",
35619 => "0101010101110000",
35620 => "0101010101110000",
35621 => "0101010101110000",
35622 => "0101010101110000",
35623 => "0101010101110000",
35624 => "0101010101110000",
35625 => "0101010101110000",
35626 => "0101010101110000",
35627 => "0101010110000000",
35628 => "0101010110000000",
35629 => "0101010110000000",
35630 => "0101010110000000",
35631 => "0101010110000000",
35632 => "0101010110000000",
35633 => "0101010110000000",
35634 => "0101010110000000",
35635 => "0101010110000000",
35636 => "0101010110010000",
35637 => "0101010110010000",
35638 => "0101010110010000",
35639 => "0101010110010000",
35640 => "0101010110010000",
35641 => "0101010110010000",
35642 => "0101010110010000",
35643 => "0101010110010000",
35644 => "0101010110010000",
35645 => "0101010110100000",
35646 => "0101010110100000",
35647 => "0101010110100000",
35648 => "0101010110100000",
35649 => "0101010110100000",
35650 => "0101010110100000",
35651 => "0101010110100000",
35652 => "0101010110100000",
35653 => "0101010110100000",
35654 => "0101010110110000",
35655 => "0101010110110000",
35656 => "0101010110110000",
35657 => "0101010110110000",
35658 => "0101010110110000",
35659 => "0101010110110000",
35660 => "0101010110110000",
35661 => "0101010110110000",
35662 => "0101010110110000",
35663 => "0101010111000000",
35664 => "0101010111000000",
35665 => "0101010111000000",
35666 => "0101010111000000",
35667 => "0101010111000000",
35668 => "0101010111000000",
35669 => "0101010111000000",
35670 => "0101010111000000",
35671 => "0101010111000000",
35672 => "0101010111010000",
35673 => "0101010111010000",
35674 => "0101010111010000",
35675 => "0101010111010000",
35676 => "0101010111010000",
35677 => "0101010111010000",
35678 => "0101010111010000",
35679 => "0101010111010000",
35680 => "0101010111010000",
35681 => "0101010111100000",
35682 => "0101010111100000",
35683 => "0101010111100000",
35684 => "0101010111100000",
35685 => "0101010111100000",
35686 => "0101010111100000",
35687 => "0101010111100000",
35688 => "0101010111100000",
35689 => "0101010111100000",
35690 => "0101010111110000",
35691 => "0101010111110000",
35692 => "0101010111110000",
35693 => "0101010111110000",
35694 => "0101010111110000",
35695 => "0101010111110000",
35696 => "0101010111110000",
35697 => "0101010111110000",
35698 => "0101010111110000",
35699 => "0101011000000000",
35700 => "0101011000000000",
35701 => "0101011000000000",
35702 => "0101011000000000",
35703 => "0101011000000000",
35704 => "0101011000000000",
35705 => "0101011000000000",
35706 => "0101011000000000",
35707 => "0101011000000000",
35708 => "0101011000010000",
35709 => "0101011000010000",
35710 => "0101011000010000",
35711 => "0101011000010000",
35712 => "0101011000010000",
35713 => "0101011000010000",
35714 => "0101011000010000",
35715 => "0101011000010000",
35716 => "0101011000010000",
35717 => "0101011000100000",
35718 => "0101011000100000",
35719 => "0101011000100000",
35720 => "0101011000100000",
35721 => "0101011000100000",
35722 => "0101011000100000",
35723 => "0101011000100000",
35724 => "0101011000100000",
35725 => "0101011000100000",
35726 => "0101011000110000",
35727 => "0101011000110000",
35728 => "0101011000110000",
35729 => "0101011000110000",
35730 => "0101011000110000",
35731 => "0101011000110000",
35732 => "0101011000110000",
35733 => "0101011000110000",
35734 => "0101011000110000",
35735 => "0101011001000000",
35736 => "0101011001000000",
35737 => "0101011001000000",
35738 => "0101011001000000",
35739 => "0101011001000000",
35740 => "0101011001000000",
35741 => "0101011001000000",
35742 => "0101011001000000",
35743 => "0101011001000000",
35744 => "0101011001010000",
35745 => "0101011001010000",
35746 => "0101011001010000",
35747 => "0101011001010000",
35748 => "0101011001010000",
35749 => "0101011001010000",
35750 => "0101011001010000",
35751 => "0101011001010000",
35752 => "0101011001010000",
35753 => "0101011001100000",
35754 => "0101011001100000",
35755 => "0101011001100000",
35756 => "0101011001100000",
35757 => "0101011001100000",
35758 => "0101011001100000",
35759 => "0101011001100000",
35760 => "0101011001100000",
35761 => "0101011001100000",
35762 => "0101011001100000",
35763 => "0101011001110000",
35764 => "0101011001110000",
35765 => "0101011001110000",
35766 => "0101011001110000",
35767 => "0101011001110000",
35768 => "0101011001110000",
35769 => "0101011001110000",
35770 => "0101011001110000",
35771 => "0101011001110000",
35772 => "0101011010000000",
35773 => "0101011010000000",
35774 => "0101011010000000",
35775 => "0101011010000000",
35776 => "0101011010000000",
35777 => "0101011010000000",
35778 => "0101011010000000",
35779 => "0101011010000000",
35780 => "0101011010000000",
35781 => "0101011010010000",
35782 => "0101011010010000",
35783 => "0101011010010000",
35784 => "0101011010010000",
35785 => "0101011010010000",
35786 => "0101011010010000",
35787 => "0101011010010000",
35788 => "0101011010010000",
35789 => "0101011010010000",
35790 => "0101011010100000",
35791 => "0101011010100000",
35792 => "0101011010100000",
35793 => "0101011010100000",
35794 => "0101011010100000",
35795 => "0101011010100000",
35796 => "0101011010100000",
35797 => "0101011010100000",
35798 => "0101011010100000",
35799 => "0101011010110000",
35800 => "0101011010110000",
35801 => "0101011010110000",
35802 => "0101011010110000",
35803 => "0101011010110000",
35804 => "0101011010110000",
35805 => "0101011010110000",
35806 => "0101011010110000",
35807 => "0101011010110000",
35808 => "0101011011000000",
35809 => "0101011011000000",
35810 => "0101011011000000",
35811 => "0101011011000000",
35812 => "0101011011000000",
35813 => "0101011011000000",
35814 => "0101011011000000",
35815 => "0101011011000000",
35816 => "0101011011000000",
35817 => "0101011011010000",
35818 => "0101011011010000",
35819 => "0101011011010000",
35820 => "0101011011010000",
35821 => "0101011011010000",
35822 => "0101011011010000",
35823 => "0101011011010000",
35824 => "0101011011010000",
35825 => "0101011011010000",
35826 => "0101011011010000",
35827 => "0101011011100000",
35828 => "0101011011100000",
35829 => "0101011011100000",
35830 => "0101011011100000",
35831 => "0101011011100000",
35832 => "0101011011100000",
35833 => "0101011011100000",
35834 => "0101011011100000",
35835 => "0101011011100000",
35836 => "0101011011110000",
35837 => "0101011011110000",
35838 => "0101011011110000",
35839 => "0101011011110000",
35840 => "0101011011110000",
35841 => "0101011011110000",
35842 => "0101011011110000",
35843 => "0101011011110000",
35844 => "0101011011110000",
35845 => "0101011100000000",
35846 => "0101011100000000",
35847 => "0101011100000000",
35848 => "0101011100000000",
35849 => "0101011100000000",
35850 => "0101011100000000",
35851 => "0101011100000000",
35852 => "0101011100000000",
35853 => "0101011100000000",
35854 => "0101011100010000",
35855 => "0101011100010000",
35856 => "0101011100010000",
35857 => "0101011100010000",
35858 => "0101011100010000",
35859 => "0101011100010000",
35860 => "0101011100010000",
35861 => "0101011100010000",
35862 => "0101011100010000",
35863 => "0101011100100000",
35864 => "0101011100100000",
35865 => "0101011100100000",
35866 => "0101011100100000",
35867 => "0101011100100000",
35868 => "0101011100100000",
35869 => "0101011100100000",
35870 => "0101011100100000",
35871 => "0101011100100000",
35872 => "0101011100100000",
35873 => "0101011100110000",
35874 => "0101011100110000",
35875 => "0101011100110000",
35876 => "0101011100110000",
35877 => "0101011100110000",
35878 => "0101011100110000",
35879 => "0101011100110000",
35880 => "0101011100110000",
35881 => "0101011100110000",
35882 => "0101011101000000",
35883 => "0101011101000000",
35884 => "0101011101000000",
35885 => "0101011101000000",
35886 => "0101011101000000",
35887 => "0101011101000000",
35888 => "0101011101000000",
35889 => "0101011101000000",
35890 => "0101011101000000",
35891 => "0101011101010000",
35892 => "0101011101010000",
35893 => "0101011101010000",
35894 => "0101011101010000",
35895 => "0101011101010000",
35896 => "0101011101010000",
35897 => "0101011101010000",
35898 => "0101011101010000",
35899 => "0101011101010000",
35900 => "0101011101100000",
35901 => "0101011101100000",
35902 => "0101011101100000",
35903 => "0101011101100000",
35904 => "0101011101100000",
35905 => "0101011101100000",
35906 => "0101011101100000",
35907 => "0101011101100000",
35908 => "0101011101100000",
35909 => "0101011101110000",
35910 => "0101011101110000",
35911 => "0101011101110000",
35912 => "0101011101110000",
35913 => "0101011101110000",
35914 => "0101011101110000",
35915 => "0101011101110000",
35916 => "0101011101110000",
35917 => "0101011101110000",
35918 => "0101011101110000",
35919 => "0101011110000000",
35920 => "0101011110000000",
35921 => "0101011110000000",
35922 => "0101011110000000",
35923 => "0101011110000000",
35924 => "0101011110000000",
35925 => "0101011110000000",
35926 => "0101011110000000",
35927 => "0101011110000000",
35928 => "0101011110010000",
35929 => "0101011110010000",
35930 => "0101011110010000",
35931 => "0101011110010000",
35932 => "0101011110010000",
35933 => "0101011110010000",
35934 => "0101011110010000",
35935 => "0101011110010000",
35936 => "0101011110010000",
35937 => "0101011110100000",
35938 => "0101011110100000",
35939 => "0101011110100000",
35940 => "0101011110100000",
35941 => "0101011110100000",
35942 => "0101011110100000",
35943 => "0101011110100000",
35944 => "0101011110100000",
35945 => "0101011110100000",
35946 => "0101011110110000",
35947 => "0101011110110000",
35948 => "0101011110110000",
35949 => "0101011110110000",
35950 => "0101011110110000",
35951 => "0101011110110000",
35952 => "0101011110110000",
35953 => "0101011110110000",
35954 => "0101011110110000",
35955 => "0101011110110000",
35956 => "0101011111000000",
35957 => "0101011111000000",
35958 => "0101011111000000",
35959 => "0101011111000000",
35960 => "0101011111000000",
35961 => "0101011111000000",
35962 => "0101011111000000",
35963 => "0101011111000000",
35964 => "0101011111000000",
35965 => "0101011111010000",
35966 => "0101011111010000",
35967 => "0101011111010000",
35968 => "0101011111010000",
35969 => "0101011111010000",
35970 => "0101011111010000",
35971 => "0101011111010000",
35972 => "0101011111010000",
35973 => "0101011111010000",
35974 => "0101011111100000",
35975 => "0101011111100000",
35976 => "0101011111100000",
35977 => "0101011111100000",
35978 => "0101011111100000",
35979 => "0101011111100000",
35980 => "0101011111100000",
35981 => "0101011111100000",
35982 => "0101011111100000",
35983 => "0101011111100000",
35984 => "0101011111110000",
35985 => "0101011111110000",
35986 => "0101011111110000",
35987 => "0101011111110000",
35988 => "0101011111110000",
35989 => "0101011111110000",
35990 => "0101011111110000",
35991 => "0101011111110000",
35992 => "0101011111110000",
35993 => "0101100000000000",
35994 => "0101100000000000",
35995 => "0101100000000000",
35996 => "0101100000000000",
35997 => "0101100000000000",
35998 => "0101100000000000",
35999 => "0101100000000000",
36000 => "0101100000000000",
36001 => "0101100000000000",
36002 => "0101100000010000",
36003 => "0101100000010000",
36004 => "0101100000010000",
36005 => "0101100000010000",
36006 => "0101100000010000",
36007 => "0101100000010000",
36008 => "0101100000010000",
36009 => "0101100000010000",
36010 => "0101100000010000",
36011 => "0101100000100000",
36012 => "0101100000100000",
36013 => "0101100000100000",
36014 => "0101100000100000",
36015 => "0101100000100000",
36016 => "0101100000100000",
36017 => "0101100000100000",
36018 => "0101100000100000",
36019 => "0101100000100000",
36020 => "0101100000100000",
36021 => "0101100000110000",
36022 => "0101100000110000",
36023 => "0101100000110000",
36024 => "0101100000110000",
36025 => "0101100000110000",
36026 => "0101100000110000",
36027 => "0101100000110000",
36028 => "0101100000110000",
36029 => "0101100000110000",
36030 => "0101100001000000",
36031 => "0101100001000000",
36032 => "0101100001000000",
36033 => "0101100001000000",
36034 => "0101100001000000",
36035 => "0101100001000000",
36036 => "0101100001000000",
36037 => "0101100001000000",
36038 => "0101100001000000",
36039 => "0101100001010000",
36040 => "0101100001010000",
36041 => "0101100001010000",
36042 => "0101100001010000",
36043 => "0101100001010000",
36044 => "0101100001010000",
36045 => "0101100001010000",
36046 => "0101100001010000",
36047 => "0101100001010000",
36048 => "0101100001010000",
36049 => "0101100001100000",
36050 => "0101100001100000",
36051 => "0101100001100000",
36052 => "0101100001100000",
36053 => "0101100001100000",
36054 => "0101100001100000",
36055 => "0101100001100000",
36056 => "0101100001100000",
36057 => "0101100001100000",
36058 => "0101100001110000",
36059 => "0101100001110000",
36060 => "0101100001110000",
36061 => "0101100001110000",
36062 => "0101100001110000",
36063 => "0101100001110000",
36064 => "0101100001110000",
36065 => "0101100001110000",
36066 => "0101100001110000",
36067 => "0101100001110000",
36068 => "0101100010000000",
36069 => "0101100010000000",
36070 => "0101100010000000",
36071 => "0101100010000000",
36072 => "0101100010000000",
36073 => "0101100010000000",
36074 => "0101100010000000",
36075 => "0101100010000000",
36076 => "0101100010000000",
36077 => "0101100010010000",
36078 => "0101100010010000",
36079 => "0101100010010000",
36080 => "0101100010010000",
36081 => "0101100010010000",
36082 => "0101100010010000",
36083 => "0101100010010000",
36084 => "0101100010010000",
36085 => "0101100010010000",
36086 => "0101100010100000",
36087 => "0101100010100000",
36088 => "0101100010100000",
36089 => "0101100010100000",
36090 => "0101100010100000",
36091 => "0101100010100000",
36092 => "0101100010100000",
36093 => "0101100010100000",
36094 => "0101100010100000",
36095 => "0101100010100000",
36096 => "0101100010110000",
36097 => "0101100010110000",
36098 => "0101100010110000",
36099 => "0101100010110000",
36100 => "0101100010110000",
36101 => "0101100010110000",
36102 => "0101100010110000",
36103 => "0101100010110000",
36104 => "0101100010110000",
36105 => "0101100011000000",
36106 => "0101100011000000",
36107 => "0101100011000000",
36108 => "0101100011000000",
36109 => "0101100011000000",
36110 => "0101100011000000",
36111 => "0101100011000000",
36112 => "0101100011000000",
36113 => "0101100011000000",
36114 => "0101100011010000",
36115 => "0101100011010000",
36116 => "0101100011010000",
36117 => "0101100011010000",
36118 => "0101100011010000",
36119 => "0101100011010000",
36120 => "0101100011010000",
36121 => "0101100011010000",
36122 => "0101100011010000",
36123 => "0101100011010000",
36124 => "0101100011100000",
36125 => "0101100011100000",
36126 => "0101100011100000",
36127 => "0101100011100000",
36128 => "0101100011100000",
36129 => "0101100011100000",
36130 => "0101100011100000",
36131 => "0101100011100000",
36132 => "0101100011100000",
36133 => "0101100011110000",
36134 => "0101100011110000",
36135 => "0101100011110000",
36136 => "0101100011110000",
36137 => "0101100011110000",
36138 => "0101100011110000",
36139 => "0101100011110000",
36140 => "0101100011110000",
36141 => "0101100011110000",
36142 => "0101100011110000",
36143 => "0101100100000000",
36144 => "0101100100000000",
36145 => "0101100100000000",
36146 => "0101100100000000",
36147 => "0101100100000000",
36148 => "0101100100000000",
36149 => "0101100100000000",
36150 => "0101100100000000",
36151 => "0101100100000000",
36152 => "0101100100010000",
36153 => "0101100100010000",
36154 => "0101100100010000",
36155 => "0101100100010000",
36156 => "0101100100010000",
36157 => "0101100100010000",
36158 => "0101100100010000",
36159 => "0101100100010000",
36160 => "0101100100010000",
36161 => "0101100100010000",
36162 => "0101100100100000",
36163 => "0101100100100000",
36164 => "0101100100100000",
36165 => "0101100100100000",
36166 => "0101100100100000",
36167 => "0101100100100000",
36168 => "0101100100100000",
36169 => "0101100100100000",
36170 => "0101100100100000",
36171 => "0101100100110000",
36172 => "0101100100110000",
36173 => "0101100100110000",
36174 => "0101100100110000",
36175 => "0101100100110000",
36176 => "0101100100110000",
36177 => "0101100100110000",
36178 => "0101100100110000",
36179 => "0101100100110000",
36180 => "0101100100110000",
36181 => "0101100101000000",
36182 => "0101100101000000",
36183 => "0101100101000000",
36184 => "0101100101000000",
36185 => "0101100101000000",
36186 => "0101100101000000",
36187 => "0101100101000000",
36188 => "0101100101000000",
36189 => "0101100101000000",
36190 => "0101100101010000",
36191 => "0101100101010000",
36192 => "0101100101010000",
36193 => "0101100101010000",
36194 => "0101100101010000",
36195 => "0101100101010000",
36196 => "0101100101010000",
36197 => "0101100101010000",
36198 => "0101100101010000",
36199 => "0101100101010000",
36200 => "0101100101100000",
36201 => "0101100101100000",
36202 => "0101100101100000",
36203 => "0101100101100000",
36204 => "0101100101100000",
36205 => "0101100101100000",
36206 => "0101100101100000",
36207 => "0101100101100000",
36208 => "0101100101100000",
36209 => "0101100101110000",
36210 => "0101100101110000",
36211 => "0101100101110000",
36212 => "0101100101110000",
36213 => "0101100101110000",
36214 => "0101100101110000",
36215 => "0101100101110000",
36216 => "0101100101110000",
36217 => "0101100101110000",
36218 => "0101100110000000",
36219 => "0101100110000000",
36220 => "0101100110000000",
36221 => "0101100110000000",
36222 => "0101100110000000",
36223 => "0101100110000000",
36224 => "0101100110000000",
36225 => "0101100110000000",
36226 => "0101100110000000",
36227 => "0101100110000000",
36228 => "0101100110010000",
36229 => "0101100110010000",
36230 => "0101100110010000",
36231 => "0101100110010000",
36232 => "0101100110010000",
36233 => "0101100110010000",
36234 => "0101100110010000",
36235 => "0101100110010000",
36236 => "0101100110010000",
36237 => "0101100110010000",
36238 => "0101100110100000",
36239 => "0101100110100000",
36240 => "0101100110100000",
36241 => "0101100110100000",
36242 => "0101100110100000",
36243 => "0101100110100000",
36244 => "0101100110100000",
36245 => "0101100110100000",
36246 => "0101100110100000",
36247 => "0101100110110000",
36248 => "0101100110110000",
36249 => "0101100110110000",
36250 => "0101100110110000",
36251 => "0101100110110000",
36252 => "0101100110110000",
36253 => "0101100110110000",
36254 => "0101100110110000",
36255 => "0101100110110000",
36256 => "0101100110110000",
36257 => "0101100111000000",
36258 => "0101100111000000",
36259 => "0101100111000000",
36260 => "0101100111000000",
36261 => "0101100111000000",
36262 => "0101100111000000",
36263 => "0101100111000000",
36264 => "0101100111000000",
36265 => "0101100111000000",
36266 => "0101100111010000",
36267 => "0101100111010000",
36268 => "0101100111010000",
36269 => "0101100111010000",
36270 => "0101100111010000",
36271 => "0101100111010000",
36272 => "0101100111010000",
36273 => "0101100111010000",
36274 => "0101100111010000",
36275 => "0101100111010000",
36276 => "0101100111100000",
36277 => "0101100111100000",
36278 => "0101100111100000",
36279 => "0101100111100000",
36280 => "0101100111100000",
36281 => "0101100111100000",
36282 => "0101100111100000",
36283 => "0101100111100000",
36284 => "0101100111100000",
36285 => "0101100111110000",
36286 => "0101100111110000",
36287 => "0101100111110000",
36288 => "0101100111110000",
36289 => "0101100111110000",
36290 => "0101100111110000",
36291 => "0101100111110000",
36292 => "0101100111110000",
36293 => "0101100111110000",
36294 => "0101100111110000",
36295 => "0101101000000000",
36296 => "0101101000000000",
36297 => "0101101000000000",
36298 => "0101101000000000",
36299 => "0101101000000000",
36300 => "0101101000000000",
36301 => "0101101000000000",
36302 => "0101101000000000",
36303 => "0101101000000000",
36304 => "0101101000010000",
36305 => "0101101000010000",
36306 => "0101101000010000",
36307 => "0101101000010000",
36308 => "0101101000010000",
36309 => "0101101000010000",
36310 => "0101101000010000",
36311 => "0101101000010000",
36312 => "0101101000010000",
36313 => "0101101000010000",
36314 => "0101101000100000",
36315 => "0101101000100000",
36316 => "0101101000100000",
36317 => "0101101000100000",
36318 => "0101101000100000",
36319 => "0101101000100000",
36320 => "0101101000100000",
36321 => "0101101000100000",
36322 => "0101101000100000",
36323 => "0101101000100000",
36324 => "0101101000110000",
36325 => "0101101000110000",
36326 => "0101101000110000",
36327 => "0101101000110000",
36328 => "0101101000110000",
36329 => "0101101000110000",
36330 => "0101101000110000",
36331 => "0101101000110000",
36332 => "0101101000110000",
36333 => "0101101001000000",
36334 => "0101101001000000",
36335 => "0101101001000000",
36336 => "0101101001000000",
36337 => "0101101001000000",
36338 => "0101101001000000",
36339 => "0101101001000000",
36340 => "0101101001000000",
36341 => "0101101001000000",
36342 => "0101101001000000",
36343 => "0101101001010000",
36344 => "0101101001010000",
36345 => "0101101001010000",
36346 => "0101101001010000",
36347 => "0101101001010000",
36348 => "0101101001010000",
36349 => "0101101001010000",
36350 => "0101101001010000",
36351 => "0101101001010000",
36352 => "0101101001100000",
36353 => "0101101001100000",
36354 => "0101101001100000",
36355 => "0101101001100000",
36356 => "0101101001100000",
36357 => "0101101001100000",
36358 => "0101101001100000",
36359 => "0101101001100000",
36360 => "0101101001100000",
36361 => "0101101001100000",
36362 => "0101101001110000",
36363 => "0101101001110000",
36364 => "0101101001110000",
36365 => "0101101001110000",
36366 => "0101101001110000",
36367 => "0101101001110000",
36368 => "0101101001110000",
36369 => "0101101001110000",
36370 => "0101101001110000",
36371 => "0101101001110000",
36372 => "0101101010000000",
36373 => "0101101010000000",
36374 => "0101101010000000",
36375 => "0101101010000000",
36376 => "0101101010000000",
36377 => "0101101010000000",
36378 => "0101101010000000",
36379 => "0101101010000000",
36380 => "0101101010000000",
36381 => "0101101010010000",
36382 => "0101101010010000",
36383 => "0101101010010000",
36384 => "0101101010010000",
36385 => "0101101010010000",
36386 => "0101101010010000",
36387 => "0101101010010000",
36388 => "0101101010010000",
36389 => "0101101010010000",
36390 => "0101101010010000",
36391 => "0101101010100000",
36392 => "0101101010100000",
36393 => "0101101010100000",
36394 => "0101101010100000",
36395 => "0101101010100000",
36396 => "0101101010100000",
36397 => "0101101010100000",
36398 => "0101101010100000",
36399 => "0101101010100000",
36400 => "0101101010100000",
36401 => "0101101010110000",
36402 => "0101101010110000",
36403 => "0101101010110000",
36404 => "0101101010110000",
36405 => "0101101010110000",
36406 => "0101101010110000",
36407 => "0101101010110000",
36408 => "0101101010110000",
36409 => "0101101010110000",
36410 => "0101101011000000",
36411 => "0101101011000000",
36412 => "0101101011000000",
36413 => "0101101011000000",
36414 => "0101101011000000",
36415 => "0101101011000000",
36416 => "0101101011000000",
36417 => "0101101011000000",
36418 => "0101101011000000",
36419 => "0101101011000000",
36420 => "0101101011010000",
36421 => "0101101011010000",
36422 => "0101101011010000",
36423 => "0101101011010000",
36424 => "0101101011010000",
36425 => "0101101011010000",
36426 => "0101101011010000",
36427 => "0101101011010000",
36428 => "0101101011010000",
36429 => "0101101011010000",
36430 => "0101101011100000",
36431 => "0101101011100000",
36432 => "0101101011100000",
36433 => "0101101011100000",
36434 => "0101101011100000",
36435 => "0101101011100000",
36436 => "0101101011100000",
36437 => "0101101011100000",
36438 => "0101101011100000",
36439 => "0101101011100000",
36440 => "0101101011110000",
36441 => "0101101011110000",
36442 => "0101101011110000",
36443 => "0101101011110000",
36444 => "0101101011110000",
36445 => "0101101011110000",
36446 => "0101101011110000",
36447 => "0101101011110000",
36448 => "0101101011110000",
36449 => "0101101100000000",
36450 => "0101101100000000",
36451 => "0101101100000000",
36452 => "0101101100000000",
36453 => "0101101100000000",
36454 => "0101101100000000",
36455 => "0101101100000000",
36456 => "0101101100000000",
36457 => "0101101100000000",
36458 => "0101101100000000",
36459 => "0101101100010000",
36460 => "0101101100010000",
36461 => "0101101100010000",
36462 => "0101101100010000",
36463 => "0101101100010000",
36464 => "0101101100010000",
36465 => "0101101100010000",
36466 => "0101101100010000",
36467 => "0101101100010000",
36468 => "0101101100010000",
36469 => "0101101100100000",
36470 => "0101101100100000",
36471 => "0101101100100000",
36472 => "0101101100100000",
36473 => "0101101100100000",
36474 => "0101101100100000",
36475 => "0101101100100000",
36476 => "0101101100100000",
36477 => "0101101100100000",
36478 => "0101101100110000",
36479 => "0101101100110000",
36480 => "0101101100110000",
36481 => "0101101100110000",
36482 => "0101101100110000",
36483 => "0101101100110000",
36484 => "0101101100110000",
36485 => "0101101100110000",
36486 => "0101101100110000",
36487 => "0101101100110000",
36488 => "0101101101000000",
36489 => "0101101101000000",
36490 => "0101101101000000",
36491 => "0101101101000000",
36492 => "0101101101000000",
36493 => "0101101101000000",
36494 => "0101101101000000",
36495 => "0101101101000000",
36496 => "0101101101000000",
36497 => "0101101101000000",
36498 => "0101101101010000",
36499 => "0101101101010000",
36500 => "0101101101010000",
36501 => "0101101101010000",
36502 => "0101101101010000",
36503 => "0101101101010000",
36504 => "0101101101010000",
36505 => "0101101101010000",
36506 => "0101101101010000",
36507 => "0101101101010000",
36508 => "0101101101100000",
36509 => "0101101101100000",
36510 => "0101101101100000",
36511 => "0101101101100000",
36512 => "0101101101100000",
36513 => "0101101101100000",
36514 => "0101101101100000",
36515 => "0101101101100000",
36516 => "0101101101100000",
36517 => "0101101101100000",
36518 => "0101101101110000",
36519 => "0101101101110000",
36520 => "0101101101110000",
36521 => "0101101101110000",
36522 => "0101101101110000",
36523 => "0101101101110000",
36524 => "0101101101110000",
36525 => "0101101101110000",
36526 => "0101101101110000",
36527 => "0101101110000000",
36528 => "0101101110000000",
36529 => "0101101110000000",
36530 => "0101101110000000",
36531 => "0101101110000000",
36532 => "0101101110000000",
36533 => "0101101110000000",
36534 => "0101101110000000",
36535 => "0101101110000000",
36536 => "0101101110000000",
36537 => "0101101110010000",
36538 => "0101101110010000",
36539 => "0101101110010000",
36540 => "0101101110010000",
36541 => "0101101110010000",
36542 => "0101101110010000",
36543 => "0101101110010000",
36544 => "0101101110010000",
36545 => "0101101110010000",
36546 => "0101101110010000",
36547 => "0101101110100000",
36548 => "0101101110100000",
36549 => "0101101110100000",
36550 => "0101101110100000",
36551 => "0101101110100000",
36552 => "0101101110100000",
36553 => "0101101110100000",
36554 => "0101101110100000",
36555 => "0101101110100000",
36556 => "0101101110100000",
36557 => "0101101110110000",
36558 => "0101101110110000",
36559 => "0101101110110000",
36560 => "0101101110110000",
36561 => "0101101110110000",
36562 => "0101101110110000",
36563 => "0101101110110000",
36564 => "0101101110110000",
36565 => "0101101110110000",
36566 => "0101101110110000",
36567 => "0101101111000000",
36568 => "0101101111000000",
36569 => "0101101111000000",
36570 => "0101101111000000",
36571 => "0101101111000000",
36572 => "0101101111000000",
36573 => "0101101111000000",
36574 => "0101101111000000",
36575 => "0101101111000000",
36576 => "0101101111000000",
36577 => "0101101111010000",
36578 => "0101101111010000",
36579 => "0101101111010000",
36580 => "0101101111010000",
36581 => "0101101111010000",
36582 => "0101101111010000",
36583 => "0101101111010000",
36584 => "0101101111010000",
36585 => "0101101111010000",
36586 => "0101101111100000",
36587 => "0101101111100000",
36588 => "0101101111100000",
36589 => "0101101111100000",
36590 => "0101101111100000",
36591 => "0101101111100000",
36592 => "0101101111100000",
36593 => "0101101111100000",
36594 => "0101101111100000",
36595 => "0101101111100000",
36596 => "0101101111110000",
36597 => "0101101111110000",
36598 => "0101101111110000",
36599 => "0101101111110000",
36600 => "0101101111110000",
36601 => "0101101111110000",
36602 => "0101101111110000",
36603 => "0101101111110000",
36604 => "0101101111110000",
36605 => "0101101111110000",
36606 => "0101110000000000",
36607 => "0101110000000000",
36608 => "0101110000000000",
36609 => "0101110000000000",
36610 => "0101110000000000",
36611 => "0101110000000000",
36612 => "0101110000000000",
36613 => "0101110000000000",
36614 => "0101110000000000",
36615 => "0101110000000000",
36616 => "0101110000010000",
36617 => "0101110000010000",
36618 => "0101110000010000",
36619 => "0101110000010000",
36620 => "0101110000010000",
36621 => "0101110000010000",
36622 => "0101110000010000",
36623 => "0101110000010000",
36624 => "0101110000010000",
36625 => "0101110000010000",
36626 => "0101110000100000",
36627 => "0101110000100000",
36628 => "0101110000100000",
36629 => "0101110000100000",
36630 => "0101110000100000",
36631 => "0101110000100000",
36632 => "0101110000100000",
36633 => "0101110000100000",
36634 => "0101110000100000",
36635 => "0101110000100000",
36636 => "0101110000110000",
36637 => "0101110000110000",
36638 => "0101110000110000",
36639 => "0101110000110000",
36640 => "0101110000110000",
36641 => "0101110000110000",
36642 => "0101110000110000",
36643 => "0101110000110000",
36644 => "0101110000110000",
36645 => "0101110000110000",
36646 => "0101110001000000",
36647 => "0101110001000000",
36648 => "0101110001000000",
36649 => "0101110001000000",
36650 => "0101110001000000",
36651 => "0101110001000000",
36652 => "0101110001000000",
36653 => "0101110001000000",
36654 => "0101110001000000",
36655 => "0101110001000000",
36656 => "0101110001010000",
36657 => "0101110001010000",
36658 => "0101110001010000",
36659 => "0101110001010000",
36660 => "0101110001010000",
36661 => "0101110001010000",
36662 => "0101110001010000",
36663 => "0101110001010000",
36664 => "0101110001010000",
36665 => "0101110001010000",
36666 => "0101110001100000",
36667 => "0101110001100000",
36668 => "0101110001100000",
36669 => "0101110001100000",
36670 => "0101110001100000",
36671 => "0101110001100000",
36672 => "0101110001100000",
36673 => "0101110001100000",
36674 => "0101110001100000",
36675 => "0101110001100000",
36676 => "0101110001110000",
36677 => "0101110001110000",
36678 => "0101110001110000",
36679 => "0101110001110000",
36680 => "0101110001110000",
36681 => "0101110001110000",
36682 => "0101110001110000",
36683 => "0101110001110000",
36684 => "0101110001110000",
36685 => "0101110001110000",
36686 => "0101110010000000",
36687 => "0101110010000000",
36688 => "0101110010000000",
36689 => "0101110010000000",
36690 => "0101110010000000",
36691 => "0101110010000000",
36692 => "0101110010000000",
36693 => "0101110010000000",
36694 => "0101110010000000",
36695 => "0101110010000000",
36696 => "0101110010010000",
36697 => "0101110010010000",
36698 => "0101110010010000",
36699 => "0101110010010000",
36700 => "0101110010010000",
36701 => "0101110010010000",
36702 => "0101110010010000",
36703 => "0101110010010000",
36704 => "0101110010010000",
36705 => "0101110010010000",
36706 => "0101110010100000",
36707 => "0101110010100000",
36708 => "0101110010100000",
36709 => "0101110010100000",
36710 => "0101110010100000",
36711 => "0101110010100000",
36712 => "0101110010100000",
36713 => "0101110010100000",
36714 => "0101110010100000",
36715 => "0101110010100000",
36716 => "0101110010110000",
36717 => "0101110010110000",
36718 => "0101110010110000",
36719 => "0101110010110000",
36720 => "0101110010110000",
36721 => "0101110010110000",
36722 => "0101110010110000",
36723 => "0101110010110000",
36724 => "0101110010110000",
36725 => "0101110010110000",
36726 => "0101110011000000",
36727 => "0101110011000000",
36728 => "0101110011000000",
36729 => "0101110011000000",
36730 => "0101110011000000",
36731 => "0101110011000000",
36732 => "0101110011000000",
36733 => "0101110011000000",
36734 => "0101110011000000",
36735 => "0101110011000000",
36736 => "0101110011010000",
36737 => "0101110011010000",
36738 => "0101110011010000",
36739 => "0101110011010000",
36740 => "0101110011010000",
36741 => "0101110011010000",
36742 => "0101110011010000",
36743 => "0101110011010000",
36744 => "0101110011010000",
36745 => "0101110011010000",
36746 => "0101110011100000",
36747 => "0101110011100000",
36748 => "0101110011100000",
36749 => "0101110011100000",
36750 => "0101110011100000",
36751 => "0101110011100000",
36752 => "0101110011100000",
36753 => "0101110011100000",
36754 => "0101110011100000",
36755 => "0101110011100000",
36756 => "0101110011110000",
36757 => "0101110011110000",
36758 => "0101110011110000",
36759 => "0101110011110000",
36760 => "0101110011110000",
36761 => "0101110011110000",
36762 => "0101110011110000",
36763 => "0101110011110000",
36764 => "0101110011110000",
36765 => "0101110011110000",
36766 => "0101110100000000",
36767 => "0101110100000000",
36768 => "0101110100000000",
36769 => "0101110100000000",
36770 => "0101110100000000",
36771 => "0101110100000000",
36772 => "0101110100000000",
36773 => "0101110100000000",
36774 => "0101110100000000",
36775 => "0101110100000000",
36776 => "0101110100010000",
36777 => "0101110100010000",
36778 => "0101110100010000",
36779 => "0101110100010000",
36780 => "0101110100010000",
36781 => "0101110100010000",
36782 => "0101110100010000",
36783 => "0101110100010000",
36784 => "0101110100010000",
36785 => "0101110100010000",
36786 => "0101110100100000",
36787 => "0101110100100000",
36788 => "0101110100100000",
36789 => "0101110100100000",
36790 => "0101110100100000",
36791 => "0101110100100000",
36792 => "0101110100100000",
36793 => "0101110100100000",
36794 => "0101110100100000",
36795 => "0101110100100000",
36796 => "0101110100110000",
36797 => "0101110100110000",
36798 => "0101110100110000",
36799 => "0101110100110000",
36800 => "0101110100110000",
36801 => "0101110100110000",
36802 => "0101110100110000",
36803 => "0101110100110000",
36804 => "0101110100110000",
36805 => "0101110100110000",
36806 => "0101110101000000",
36807 => "0101110101000000",
36808 => "0101110101000000",
36809 => "0101110101000000",
36810 => "0101110101000000",
36811 => "0101110101000000",
36812 => "0101110101000000",
36813 => "0101110101000000",
36814 => "0101110101000000",
36815 => "0101110101000000",
36816 => "0101110101010000",
36817 => "0101110101010000",
36818 => "0101110101010000",
36819 => "0101110101010000",
36820 => "0101110101010000",
36821 => "0101110101010000",
36822 => "0101110101010000",
36823 => "0101110101010000",
36824 => "0101110101010000",
36825 => "0101110101010000",
36826 => "0101110101100000",
36827 => "0101110101100000",
36828 => "0101110101100000",
36829 => "0101110101100000",
36830 => "0101110101100000",
36831 => "0101110101100000",
36832 => "0101110101100000",
36833 => "0101110101100000",
36834 => "0101110101100000",
36835 => "0101110101100000",
36836 => "0101110101110000",
36837 => "0101110101110000",
36838 => "0101110101110000",
36839 => "0101110101110000",
36840 => "0101110101110000",
36841 => "0101110101110000",
36842 => "0101110101110000",
36843 => "0101110101110000",
36844 => "0101110101110000",
36845 => "0101110101110000",
36846 => "0101110101110000",
36847 => "0101110110000000",
36848 => "0101110110000000",
36849 => "0101110110000000",
36850 => "0101110110000000",
36851 => "0101110110000000",
36852 => "0101110110000000",
36853 => "0101110110000000",
36854 => "0101110110000000",
36855 => "0101110110000000",
36856 => "0101110110000000",
36857 => "0101110110010000",
36858 => "0101110110010000",
36859 => "0101110110010000",
36860 => "0101110110010000",
36861 => "0101110110010000",
36862 => "0101110110010000",
36863 => "0101110110010000",
36864 => "0101110110010000",
36865 => "0101110110010000",
36866 => "0101110110010000",
36867 => "0101110110100000",
36868 => "0101110110100000",
36869 => "0101110110100000",
36870 => "0101110110100000",
36871 => "0101110110100000",
36872 => "0101110110100000",
36873 => "0101110110100000",
36874 => "0101110110100000",
36875 => "0101110110100000",
36876 => "0101110110100000",
36877 => "0101110110110000",
36878 => "0101110110110000",
36879 => "0101110110110000",
36880 => "0101110110110000",
36881 => "0101110110110000",
36882 => "0101110110110000",
36883 => "0101110110110000",
36884 => "0101110110110000",
36885 => "0101110110110000",
36886 => "0101110110110000",
36887 => "0101110111000000",
36888 => "0101110111000000",
36889 => "0101110111000000",
36890 => "0101110111000000",
36891 => "0101110111000000",
36892 => "0101110111000000",
36893 => "0101110111000000",
36894 => "0101110111000000",
36895 => "0101110111000000",
36896 => "0101110111000000",
36897 => "0101110111010000",
36898 => "0101110111010000",
36899 => "0101110111010000",
36900 => "0101110111010000",
36901 => "0101110111010000",
36902 => "0101110111010000",
36903 => "0101110111010000",
36904 => "0101110111010000",
36905 => "0101110111010000",
36906 => "0101110111010000",
36907 => "0101110111010000",
36908 => "0101110111100000",
36909 => "0101110111100000",
36910 => "0101110111100000",
36911 => "0101110111100000",
36912 => "0101110111100000",
36913 => "0101110111100000",
36914 => "0101110111100000",
36915 => "0101110111100000",
36916 => "0101110111100000",
36917 => "0101110111100000",
36918 => "0101110111110000",
36919 => "0101110111110000",
36920 => "0101110111110000",
36921 => "0101110111110000",
36922 => "0101110111110000",
36923 => "0101110111110000",
36924 => "0101110111110000",
36925 => "0101110111110000",
36926 => "0101110111110000",
36927 => "0101110111110000",
36928 => "0101111000000000",
36929 => "0101111000000000",
36930 => "0101111000000000",
36931 => "0101111000000000",
36932 => "0101111000000000",
36933 => "0101111000000000",
36934 => "0101111000000000",
36935 => "0101111000000000",
36936 => "0101111000000000",
36937 => "0101111000000000",
36938 => "0101111000010000",
36939 => "0101111000010000",
36940 => "0101111000010000",
36941 => "0101111000010000",
36942 => "0101111000010000",
36943 => "0101111000010000",
36944 => "0101111000010000",
36945 => "0101111000010000",
36946 => "0101111000010000",
36947 => "0101111000010000",
36948 => "0101111000010000",
36949 => "0101111000100000",
36950 => "0101111000100000",
36951 => "0101111000100000",
36952 => "0101111000100000",
36953 => "0101111000100000",
36954 => "0101111000100000",
36955 => "0101111000100000",
36956 => "0101111000100000",
36957 => "0101111000100000",
36958 => "0101111000100000",
36959 => "0101111000110000",
36960 => "0101111000110000",
36961 => "0101111000110000",
36962 => "0101111000110000",
36963 => "0101111000110000",
36964 => "0101111000110000",
36965 => "0101111000110000",
36966 => "0101111000110000",
36967 => "0101111000110000",
36968 => "0101111000110000",
36969 => "0101111001000000",
36970 => "0101111001000000",
36971 => "0101111001000000",
36972 => "0101111001000000",
36973 => "0101111001000000",
36974 => "0101111001000000",
36975 => "0101111001000000",
36976 => "0101111001000000",
36977 => "0101111001000000",
36978 => "0101111001000000",
36979 => "0101111001000000",
36980 => "0101111001010000",
36981 => "0101111001010000",
36982 => "0101111001010000",
36983 => "0101111001010000",
36984 => "0101111001010000",
36985 => "0101111001010000",
36986 => "0101111001010000",
36987 => "0101111001010000",
36988 => "0101111001010000",
36989 => "0101111001010000",
36990 => "0101111001100000",
36991 => "0101111001100000",
36992 => "0101111001100000",
36993 => "0101111001100000",
36994 => "0101111001100000",
36995 => "0101111001100000",
36996 => "0101111001100000",
36997 => "0101111001100000",
36998 => "0101111001100000",
36999 => "0101111001100000",
37000 => "0101111001110000",
37001 => "0101111001110000",
37002 => "0101111001110000",
37003 => "0101111001110000",
37004 => "0101111001110000",
37005 => "0101111001110000",
37006 => "0101111001110000",
37007 => "0101111001110000",
37008 => "0101111001110000",
37009 => "0101111001110000",
37010 => "0101111001110000",
37011 => "0101111010000000",
37012 => "0101111010000000",
37013 => "0101111010000000",
37014 => "0101111010000000",
37015 => "0101111010000000",
37016 => "0101111010000000",
37017 => "0101111010000000",
37018 => "0101111010000000",
37019 => "0101111010000000",
37020 => "0101111010000000",
37021 => "0101111010010000",
37022 => "0101111010010000",
37023 => "0101111010010000",
37024 => "0101111010010000",
37025 => "0101111010010000",
37026 => "0101111010010000",
37027 => "0101111010010000",
37028 => "0101111010010000",
37029 => "0101111010010000",
37030 => "0101111010010000",
37031 => "0101111010100000",
37032 => "0101111010100000",
37033 => "0101111010100000",
37034 => "0101111010100000",
37035 => "0101111010100000",
37036 => "0101111010100000",
37037 => "0101111010100000",
37038 => "0101111010100000",
37039 => "0101111010100000",
37040 => "0101111010100000",
37041 => "0101111010100000",
37042 => "0101111010110000",
37043 => "0101111010110000",
37044 => "0101111010110000",
37045 => "0101111010110000",
37046 => "0101111010110000",
37047 => "0101111010110000",
37048 => "0101111010110000",
37049 => "0101111010110000",
37050 => "0101111010110000",
37051 => "0101111010110000",
37052 => "0101111011000000",
37053 => "0101111011000000",
37054 => "0101111011000000",
37055 => "0101111011000000",
37056 => "0101111011000000",
37057 => "0101111011000000",
37058 => "0101111011000000",
37059 => "0101111011000000",
37060 => "0101111011000000",
37061 => "0101111011000000",
37062 => "0101111011010000",
37063 => "0101111011010000",
37064 => "0101111011010000",
37065 => "0101111011010000",
37066 => "0101111011010000",
37067 => "0101111011010000",
37068 => "0101111011010000",
37069 => "0101111011010000",
37070 => "0101111011010000",
37071 => "0101111011010000",
37072 => "0101111011010000",
37073 => "0101111011100000",
37074 => "0101111011100000",
37075 => "0101111011100000",
37076 => "0101111011100000",
37077 => "0101111011100000",
37078 => "0101111011100000",
37079 => "0101111011100000",
37080 => "0101111011100000",
37081 => "0101111011100000",
37082 => "0101111011100000",
37083 => "0101111011110000",
37084 => "0101111011110000",
37085 => "0101111011110000",
37086 => "0101111011110000",
37087 => "0101111011110000",
37088 => "0101111011110000",
37089 => "0101111011110000",
37090 => "0101111011110000",
37091 => "0101111011110000",
37092 => "0101111011110000",
37093 => "0101111011110000",
37094 => "0101111100000000",
37095 => "0101111100000000",
37096 => "0101111100000000",
37097 => "0101111100000000",
37098 => "0101111100000000",
37099 => "0101111100000000",
37100 => "0101111100000000",
37101 => "0101111100000000",
37102 => "0101111100000000",
37103 => "0101111100000000",
37104 => "0101111100010000",
37105 => "0101111100010000",
37106 => "0101111100010000",
37107 => "0101111100010000",
37108 => "0101111100010000",
37109 => "0101111100010000",
37110 => "0101111100010000",
37111 => "0101111100010000",
37112 => "0101111100010000",
37113 => "0101111100010000",
37114 => "0101111100010000",
37115 => "0101111100100000",
37116 => "0101111100100000",
37117 => "0101111100100000",
37118 => "0101111100100000",
37119 => "0101111100100000",
37120 => "0101111100100000",
37121 => "0101111100100000",
37122 => "0101111100100000",
37123 => "0101111100100000",
37124 => "0101111100100000",
37125 => "0101111100110000",
37126 => "0101111100110000",
37127 => "0101111100110000",
37128 => "0101111100110000",
37129 => "0101111100110000",
37130 => "0101111100110000",
37131 => "0101111100110000",
37132 => "0101111100110000",
37133 => "0101111100110000",
37134 => "0101111100110000",
37135 => "0101111100110000",
37136 => "0101111101000000",
37137 => "0101111101000000",
37138 => "0101111101000000",
37139 => "0101111101000000",
37140 => "0101111101000000",
37141 => "0101111101000000",
37142 => "0101111101000000",
37143 => "0101111101000000",
37144 => "0101111101000000",
37145 => "0101111101000000",
37146 => "0101111101010000",
37147 => "0101111101010000",
37148 => "0101111101010000",
37149 => "0101111101010000",
37150 => "0101111101010000",
37151 => "0101111101010000",
37152 => "0101111101010000",
37153 => "0101111101010000",
37154 => "0101111101010000",
37155 => "0101111101010000",
37156 => "0101111101010000",
37157 => "0101111101100000",
37158 => "0101111101100000",
37159 => "0101111101100000",
37160 => "0101111101100000",
37161 => "0101111101100000",
37162 => "0101111101100000",
37163 => "0101111101100000",
37164 => "0101111101100000",
37165 => "0101111101100000",
37166 => "0101111101100000",
37167 => "0101111101110000",
37168 => "0101111101110000",
37169 => "0101111101110000",
37170 => "0101111101110000",
37171 => "0101111101110000",
37172 => "0101111101110000",
37173 => "0101111101110000",
37174 => "0101111101110000",
37175 => "0101111101110000",
37176 => "0101111101110000",
37177 => "0101111101110000",
37178 => "0101111110000000",
37179 => "0101111110000000",
37180 => "0101111110000000",
37181 => "0101111110000000",
37182 => "0101111110000000",
37183 => "0101111110000000",
37184 => "0101111110000000",
37185 => "0101111110000000",
37186 => "0101111110000000",
37187 => "0101111110000000",
37188 => "0101111110010000",
37189 => "0101111110010000",
37190 => "0101111110010000",
37191 => "0101111110010000",
37192 => "0101111110010000",
37193 => "0101111110010000",
37194 => "0101111110010000",
37195 => "0101111110010000",
37196 => "0101111110010000",
37197 => "0101111110010000",
37198 => "0101111110010000",
37199 => "0101111110100000",
37200 => "0101111110100000",
37201 => "0101111110100000",
37202 => "0101111110100000",
37203 => "0101111110100000",
37204 => "0101111110100000",
37205 => "0101111110100000",
37206 => "0101111110100000",
37207 => "0101111110100000",
37208 => "0101111110100000",
37209 => "0101111110110000",
37210 => "0101111110110000",
37211 => "0101111110110000",
37212 => "0101111110110000",
37213 => "0101111110110000",
37214 => "0101111110110000",
37215 => "0101111110110000",
37216 => "0101111110110000",
37217 => "0101111110110000",
37218 => "0101111110110000",
37219 => "0101111110110000",
37220 => "0101111111000000",
37221 => "0101111111000000",
37222 => "0101111111000000",
37223 => "0101111111000000",
37224 => "0101111111000000",
37225 => "0101111111000000",
37226 => "0101111111000000",
37227 => "0101111111000000",
37228 => "0101111111000000",
37229 => "0101111111000000",
37230 => "0101111111000000",
37231 => "0101111111010000",
37232 => "0101111111010000",
37233 => "0101111111010000",
37234 => "0101111111010000",
37235 => "0101111111010000",
37236 => "0101111111010000",
37237 => "0101111111010000",
37238 => "0101111111010000",
37239 => "0101111111010000",
37240 => "0101111111010000",
37241 => "0101111111100000",
37242 => "0101111111100000",
37243 => "0101111111100000",
37244 => "0101111111100000",
37245 => "0101111111100000",
37246 => "0101111111100000",
37247 => "0101111111100000",
37248 => "0101111111100000",
37249 => "0101111111100000",
37250 => "0101111111100000",
37251 => "0101111111100000",
37252 => "0101111111110000",
37253 => "0101111111110000",
37254 => "0101111111110000",
37255 => "0101111111110000",
37256 => "0101111111110000",
37257 => "0101111111110000",
37258 => "0101111111110000",
37259 => "0101111111110000",
37260 => "0101111111110000",
37261 => "0101111111110000",
37262 => "0101111111110000",
37263 => "0110000000000000",
37264 => "0110000000000000",
37265 => "0110000000000000",
37266 => "0110000000000000",
37267 => "0110000000000000",
37268 => "0110000000000000",
37269 => "0110000000000000",
37270 => "0110000000000000",
37271 => "0110000000000000",
37272 => "0110000000000000",
37273 => "0110000000010000",
37274 => "0110000000010000",
37275 => "0110000000010000",
37276 => "0110000000010000",
37277 => "0110000000010000",
37278 => "0110000000010000",
37279 => "0110000000010000",
37280 => "0110000000010000",
37281 => "0110000000010000",
37282 => "0110000000010000",
37283 => "0110000000010000",
37284 => "0110000000100000",
37285 => "0110000000100000",
37286 => "0110000000100000",
37287 => "0110000000100000",
37288 => "0110000000100000",
37289 => "0110000000100000",
37290 => "0110000000100000",
37291 => "0110000000100000",
37292 => "0110000000100000",
37293 => "0110000000100000",
37294 => "0110000000100000",
37295 => "0110000000110000",
37296 => "0110000000110000",
37297 => "0110000000110000",
37298 => "0110000000110000",
37299 => "0110000000110000",
37300 => "0110000000110000",
37301 => "0110000000110000",
37302 => "0110000000110000",
37303 => "0110000000110000",
37304 => "0110000000110000",
37305 => "0110000001000000",
37306 => "0110000001000000",
37307 => "0110000001000000",
37308 => "0110000001000000",
37309 => "0110000001000000",
37310 => "0110000001000000",
37311 => "0110000001000000",
37312 => "0110000001000000",
37313 => "0110000001000000",
37314 => "0110000001000000",
37315 => "0110000001000000",
37316 => "0110000001010000",
37317 => "0110000001010000",
37318 => "0110000001010000",
37319 => "0110000001010000",
37320 => "0110000001010000",
37321 => "0110000001010000",
37322 => "0110000001010000",
37323 => "0110000001010000",
37324 => "0110000001010000",
37325 => "0110000001010000",
37326 => "0110000001010000",
37327 => "0110000001100000",
37328 => "0110000001100000",
37329 => "0110000001100000",
37330 => "0110000001100000",
37331 => "0110000001100000",
37332 => "0110000001100000",
37333 => "0110000001100000",
37334 => "0110000001100000",
37335 => "0110000001100000",
37336 => "0110000001100000",
37337 => "0110000001110000",
37338 => "0110000001110000",
37339 => "0110000001110000",
37340 => "0110000001110000",
37341 => "0110000001110000",
37342 => "0110000001110000",
37343 => "0110000001110000",
37344 => "0110000001110000",
37345 => "0110000001110000",
37346 => "0110000001110000",
37347 => "0110000001110000",
37348 => "0110000010000000",
37349 => "0110000010000000",
37350 => "0110000010000000",
37351 => "0110000010000000",
37352 => "0110000010000000",
37353 => "0110000010000000",
37354 => "0110000010000000",
37355 => "0110000010000000",
37356 => "0110000010000000",
37357 => "0110000010000000",
37358 => "0110000010000000",
37359 => "0110000010010000",
37360 => "0110000010010000",
37361 => "0110000010010000",
37362 => "0110000010010000",
37363 => "0110000010010000",
37364 => "0110000010010000",
37365 => "0110000010010000",
37366 => "0110000010010000",
37367 => "0110000010010000",
37368 => "0110000010010000",
37369 => "0110000010010000",
37370 => "0110000010100000",
37371 => "0110000010100000",
37372 => "0110000010100000",
37373 => "0110000010100000",
37374 => "0110000010100000",
37375 => "0110000010100000",
37376 => "0110000010100000",
37377 => "0110000010100000",
37378 => "0110000010100000",
37379 => "0110000010100000",
37380 => "0110000010100000",
37381 => "0110000010110000",
37382 => "0110000010110000",
37383 => "0110000010110000",
37384 => "0110000010110000",
37385 => "0110000010110000",
37386 => "0110000010110000",
37387 => "0110000010110000",
37388 => "0110000010110000",
37389 => "0110000010110000",
37390 => "0110000010110000",
37391 => "0110000011000000",
37392 => "0110000011000000",
37393 => "0110000011000000",
37394 => "0110000011000000",
37395 => "0110000011000000",
37396 => "0110000011000000",
37397 => "0110000011000000",
37398 => "0110000011000000",
37399 => "0110000011000000",
37400 => "0110000011000000",
37401 => "0110000011000000",
37402 => "0110000011010000",
37403 => "0110000011010000",
37404 => "0110000011010000",
37405 => "0110000011010000",
37406 => "0110000011010000",
37407 => "0110000011010000",
37408 => "0110000011010000",
37409 => "0110000011010000",
37410 => "0110000011010000",
37411 => "0110000011010000",
37412 => "0110000011010000",
37413 => "0110000011100000",
37414 => "0110000011100000",
37415 => "0110000011100000",
37416 => "0110000011100000",
37417 => "0110000011100000",
37418 => "0110000011100000",
37419 => "0110000011100000",
37420 => "0110000011100000",
37421 => "0110000011100000",
37422 => "0110000011100000",
37423 => "0110000011100000",
37424 => "0110000011110000",
37425 => "0110000011110000",
37426 => "0110000011110000",
37427 => "0110000011110000",
37428 => "0110000011110000",
37429 => "0110000011110000",
37430 => "0110000011110000",
37431 => "0110000011110000",
37432 => "0110000011110000",
37433 => "0110000011110000",
37434 => "0110000011110000",
37435 => "0110000100000000",
37436 => "0110000100000000",
37437 => "0110000100000000",
37438 => "0110000100000000",
37439 => "0110000100000000",
37440 => "0110000100000000",
37441 => "0110000100000000",
37442 => "0110000100000000",
37443 => "0110000100000000",
37444 => "0110000100000000",
37445 => "0110000100000000",
37446 => "0110000100010000",
37447 => "0110000100010000",
37448 => "0110000100010000",
37449 => "0110000100010000",
37450 => "0110000100010000",
37451 => "0110000100010000",
37452 => "0110000100010000",
37453 => "0110000100010000",
37454 => "0110000100010000",
37455 => "0110000100010000",
37456 => "0110000100010000",
37457 => "0110000100100000",
37458 => "0110000100100000",
37459 => "0110000100100000",
37460 => "0110000100100000",
37461 => "0110000100100000",
37462 => "0110000100100000",
37463 => "0110000100100000",
37464 => "0110000100100000",
37465 => "0110000100100000",
37466 => "0110000100100000",
37467 => "0110000100100000",
37468 => "0110000100110000",
37469 => "0110000100110000",
37470 => "0110000100110000",
37471 => "0110000100110000",
37472 => "0110000100110000",
37473 => "0110000100110000",
37474 => "0110000100110000",
37475 => "0110000100110000",
37476 => "0110000100110000",
37477 => "0110000100110000",
37478 => "0110000100110000",
37479 => "0110000101000000",
37480 => "0110000101000000",
37481 => "0110000101000000",
37482 => "0110000101000000",
37483 => "0110000101000000",
37484 => "0110000101000000",
37485 => "0110000101000000",
37486 => "0110000101000000",
37487 => "0110000101000000",
37488 => "0110000101000000",
37489 => "0110000101000000",
37490 => "0110000101010000",
37491 => "0110000101010000",
37492 => "0110000101010000",
37493 => "0110000101010000",
37494 => "0110000101010000",
37495 => "0110000101010000",
37496 => "0110000101010000",
37497 => "0110000101010000",
37498 => "0110000101010000",
37499 => "0110000101010000",
37500 => "0110000101100000",
37501 => "0110000101100000",
37502 => "0110000101100000",
37503 => "0110000101100000",
37504 => "0110000101100000",
37505 => "0110000101100000",
37506 => "0110000101100000",
37507 => "0110000101100000",
37508 => "0110000101100000",
37509 => "0110000101100000",
37510 => "0110000101100000",
37511 => "0110000101110000",
37512 => "0110000101110000",
37513 => "0110000101110000",
37514 => "0110000101110000",
37515 => "0110000101110000",
37516 => "0110000101110000",
37517 => "0110000101110000",
37518 => "0110000101110000",
37519 => "0110000101110000",
37520 => "0110000101110000",
37521 => "0110000101110000",
37522 => "0110000110000000",
37523 => "0110000110000000",
37524 => "0110000110000000",
37525 => "0110000110000000",
37526 => "0110000110000000",
37527 => "0110000110000000",
37528 => "0110000110000000",
37529 => "0110000110000000",
37530 => "0110000110000000",
37531 => "0110000110000000",
37532 => "0110000110000000",
37533 => "0110000110000000",
37534 => "0110000110010000",
37535 => "0110000110010000",
37536 => "0110000110010000",
37537 => "0110000110010000",
37538 => "0110000110010000",
37539 => "0110000110010000",
37540 => "0110000110010000",
37541 => "0110000110010000",
37542 => "0110000110010000",
37543 => "0110000110010000",
37544 => "0110000110010000",
37545 => "0110000110100000",
37546 => "0110000110100000",
37547 => "0110000110100000",
37548 => "0110000110100000",
37549 => "0110000110100000",
37550 => "0110000110100000",
37551 => "0110000110100000",
37552 => "0110000110100000",
37553 => "0110000110100000",
37554 => "0110000110100000",
37555 => "0110000110100000",
37556 => "0110000110110000",
37557 => "0110000110110000",
37558 => "0110000110110000",
37559 => "0110000110110000",
37560 => "0110000110110000",
37561 => "0110000110110000",
37562 => "0110000110110000",
37563 => "0110000110110000",
37564 => "0110000110110000",
37565 => "0110000110110000",
37566 => "0110000110110000",
37567 => "0110000111000000",
37568 => "0110000111000000",
37569 => "0110000111000000",
37570 => "0110000111000000",
37571 => "0110000111000000",
37572 => "0110000111000000",
37573 => "0110000111000000",
37574 => "0110000111000000",
37575 => "0110000111000000",
37576 => "0110000111000000",
37577 => "0110000111000000",
37578 => "0110000111010000",
37579 => "0110000111010000",
37580 => "0110000111010000",
37581 => "0110000111010000",
37582 => "0110000111010000",
37583 => "0110000111010000",
37584 => "0110000111010000",
37585 => "0110000111010000",
37586 => "0110000111010000",
37587 => "0110000111010000",
37588 => "0110000111010000",
37589 => "0110000111100000",
37590 => "0110000111100000",
37591 => "0110000111100000",
37592 => "0110000111100000",
37593 => "0110000111100000",
37594 => "0110000111100000",
37595 => "0110000111100000",
37596 => "0110000111100000",
37597 => "0110000111100000",
37598 => "0110000111100000",
37599 => "0110000111100000",
37600 => "0110000111110000",
37601 => "0110000111110000",
37602 => "0110000111110000",
37603 => "0110000111110000",
37604 => "0110000111110000",
37605 => "0110000111110000",
37606 => "0110000111110000",
37607 => "0110000111110000",
37608 => "0110000111110000",
37609 => "0110000111110000",
37610 => "0110000111110000",
37611 => "0110001000000000",
37612 => "0110001000000000",
37613 => "0110001000000000",
37614 => "0110001000000000",
37615 => "0110001000000000",
37616 => "0110001000000000",
37617 => "0110001000000000",
37618 => "0110001000000000",
37619 => "0110001000000000",
37620 => "0110001000000000",
37621 => "0110001000000000",
37622 => "0110001000010000",
37623 => "0110001000010000",
37624 => "0110001000010000",
37625 => "0110001000010000",
37626 => "0110001000010000",
37627 => "0110001000010000",
37628 => "0110001000010000",
37629 => "0110001000010000",
37630 => "0110001000010000",
37631 => "0110001000010000",
37632 => "0110001000010000",
37633 => "0110001000100000",
37634 => "0110001000100000",
37635 => "0110001000100000",
37636 => "0110001000100000",
37637 => "0110001000100000",
37638 => "0110001000100000",
37639 => "0110001000100000",
37640 => "0110001000100000",
37641 => "0110001000100000",
37642 => "0110001000100000",
37643 => "0110001000100000",
37644 => "0110001000100000",
37645 => "0110001000110000",
37646 => "0110001000110000",
37647 => "0110001000110000",
37648 => "0110001000110000",
37649 => "0110001000110000",
37650 => "0110001000110000",
37651 => "0110001000110000",
37652 => "0110001000110000",
37653 => "0110001000110000",
37654 => "0110001000110000",
37655 => "0110001000110000",
37656 => "0110001001000000",
37657 => "0110001001000000",
37658 => "0110001001000000",
37659 => "0110001001000000",
37660 => "0110001001000000",
37661 => "0110001001000000",
37662 => "0110001001000000",
37663 => "0110001001000000",
37664 => "0110001001000000",
37665 => "0110001001000000",
37666 => "0110001001000000",
37667 => "0110001001010000",
37668 => "0110001001010000",
37669 => "0110001001010000",
37670 => "0110001001010000",
37671 => "0110001001010000",
37672 => "0110001001010000",
37673 => "0110001001010000",
37674 => "0110001001010000",
37675 => "0110001001010000",
37676 => "0110001001010000",
37677 => "0110001001010000",
37678 => "0110001001100000",
37679 => "0110001001100000",
37680 => "0110001001100000",
37681 => "0110001001100000",
37682 => "0110001001100000",
37683 => "0110001001100000",
37684 => "0110001001100000",
37685 => "0110001001100000",
37686 => "0110001001100000",
37687 => "0110001001100000",
37688 => "0110001001100000",
37689 => "0110001001110000",
37690 => "0110001001110000",
37691 => "0110001001110000",
37692 => "0110001001110000",
37693 => "0110001001110000",
37694 => "0110001001110000",
37695 => "0110001001110000",
37696 => "0110001001110000",
37697 => "0110001001110000",
37698 => "0110001001110000",
37699 => "0110001001110000",
37700 => "0110001001110000",
37701 => "0110001010000000",
37702 => "0110001010000000",
37703 => "0110001010000000",
37704 => "0110001010000000",
37705 => "0110001010000000",
37706 => "0110001010000000",
37707 => "0110001010000000",
37708 => "0110001010000000",
37709 => "0110001010000000",
37710 => "0110001010000000",
37711 => "0110001010000000",
37712 => "0110001010010000",
37713 => "0110001010010000",
37714 => "0110001010010000",
37715 => "0110001010010000",
37716 => "0110001010010000",
37717 => "0110001010010000",
37718 => "0110001010010000",
37719 => "0110001010010000",
37720 => "0110001010010000",
37721 => "0110001010010000",
37722 => "0110001010010000",
37723 => "0110001010100000",
37724 => "0110001010100000",
37725 => "0110001010100000",
37726 => "0110001010100000",
37727 => "0110001010100000",
37728 => "0110001010100000",
37729 => "0110001010100000",
37730 => "0110001010100000",
37731 => "0110001010100000",
37732 => "0110001010100000",
37733 => "0110001010100000",
37734 => "0110001010100000",
37735 => "0110001010110000",
37736 => "0110001010110000",
37737 => "0110001010110000",
37738 => "0110001010110000",
37739 => "0110001010110000",
37740 => "0110001010110000",
37741 => "0110001010110000",
37742 => "0110001010110000",
37743 => "0110001010110000",
37744 => "0110001010110000",
37745 => "0110001010110000",
37746 => "0110001011000000",
37747 => "0110001011000000",
37748 => "0110001011000000",
37749 => "0110001011000000",
37750 => "0110001011000000",
37751 => "0110001011000000",
37752 => "0110001011000000",
37753 => "0110001011000000",
37754 => "0110001011000000",
37755 => "0110001011000000",
37756 => "0110001011000000",
37757 => "0110001011010000",
37758 => "0110001011010000",
37759 => "0110001011010000",
37760 => "0110001011010000",
37761 => "0110001011010000",
37762 => "0110001011010000",
37763 => "0110001011010000",
37764 => "0110001011010000",
37765 => "0110001011010000",
37766 => "0110001011010000",
37767 => "0110001011010000",
37768 => "0110001011010000",
37769 => "0110001011100000",
37770 => "0110001011100000",
37771 => "0110001011100000",
37772 => "0110001011100000",
37773 => "0110001011100000",
37774 => "0110001011100000",
37775 => "0110001011100000",
37776 => "0110001011100000",
37777 => "0110001011100000",
37778 => "0110001011100000",
37779 => "0110001011100000",
37780 => "0110001011110000",
37781 => "0110001011110000",
37782 => "0110001011110000",
37783 => "0110001011110000",
37784 => "0110001011110000",
37785 => "0110001011110000",
37786 => "0110001011110000",
37787 => "0110001011110000",
37788 => "0110001011110000",
37789 => "0110001011110000",
37790 => "0110001011110000",
37791 => "0110001100000000",
37792 => "0110001100000000",
37793 => "0110001100000000",
37794 => "0110001100000000",
37795 => "0110001100000000",
37796 => "0110001100000000",
37797 => "0110001100000000",
37798 => "0110001100000000",
37799 => "0110001100000000",
37800 => "0110001100000000",
37801 => "0110001100000000",
37802 => "0110001100000000",
37803 => "0110001100010000",
37804 => "0110001100010000",
37805 => "0110001100010000",
37806 => "0110001100010000",
37807 => "0110001100010000",
37808 => "0110001100010000",
37809 => "0110001100010000",
37810 => "0110001100010000",
37811 => "0110001100010000",
37812 => "0110001100010000",
37813 => "0110001100010000",
37814 => "0110001100100000",
37815 => "0110001100100000",
37816 => "0110001100100000",
37817 => "0110001100100000",
37818 => "0110001100100000",
37819 => "0110001100100000",
37820 => "0110001100100000",
37821 => "0110001100100000",
37822 => "0110001100100000",
37823 => "0110001100100000",
37824 => "0110001100100000",
37825 => "0110001100100000",
37826 => "0110001100110000",
37827 => "0110001100110000",
37828 => "0110001100110000",
37829 => "0110001100110000",
37830 => "0110001100110000",
37831 => "0110001100110000",
37832 => "0110001100110000",
37833 => "0110001100110000",
37834 => "0110001100110000",
37835 => "0110001100110000",
37836 => "0110001100110000",
37837 => "0110001101000000",
37838 => "0110001101000000",
37839 => "0110001101000000",
37840 => "0110001101000000",
37841 => "0110001101000000",
37842 => "0110001101000000",
37843 => "0110001101000000",
37844 => "0110001101000000",
37845 => "0110001101000000",
37846 => "0110001101000000",
37847 => "0110001101000000",
37848 => "0110001101000000",
37849 => "0110001101010000",
37850 => "0110001101010000",
37851 => "0110001101010000",
37852 => "0110001101010000",
37853 => "0110001101010000",
37854 => "0110001101010000",
37855 => "0110001101010000",
37856 => "0110001101010000",
37857 => "0110001101010000",
37858 => "0110001101010000",
37859 => "0110001101010000",
37860 => "0110001101100000",
37861 => "0110001101100000",
37862 => "0110001101100000",
37863 => "0110001101100000",
37864 => "0110001101100000",
37865 => "0110001101100000",
37866 => "0110001101100000",
37867 => "0110001101100000",
37868 => "0110001101100000",
37869 => "0110001101100000",
37870 => "0110001101100000",
37871 => "0110001101100000",
37872 => "0110001101110000",
37873 => "0110001101110000",
37874 => "0110001101110000",
37875 => "0110001101110000",
37876 => "0110001101110000",
37877 => "0110001101110000",
37878 => "0110001101110000",
37879 => "0110001101110000",
37880 => "0110001101110000",
37881 => "0110001101110000",
37882 => "0110001101110000",
37883 => "0110001110000000",
37884 => "0110001110000000",
37885 => "0110001110000000",
37886 => "0110001110000000",
37887 => "0110001110000000",
37888 => "0110001110000000",
37889 => "0110001110000000",
37890 => "0110001110000000",
37891 => "0110001110000000",
37892 => "0110001110000000",
37893 => "0110001110000000",
37894 => "0110001110000000",
37895 => "0110001110010000",
37896 => "0110001110010000",
37897 => "0110001110010000",
37898 => "0110001110010000",
37899 => "0110001110010000",
37900 => "0110001110010000",
37901 => "0110001110010000",
37902 => "0110001110010000",
37903 => "0110001110010000",
37904 => "0110001110010000",
37905 => "0110001110010000",
37906 => "0110001110100000",
37907 => "0110001110100000",
37908 => "0110001110100000",
37909 => "0110001110100000",
37910 => "0110001110100000",
37911 => "0110001110100000",
37912 => "0110001110100000",
37913 => "0110001110100000",
37914 => "0110001110100000",
37915 => "0110001110100000",
37916 => "0110001110100000",
37917 => "0110001110100000",
37918 => "0110001110110000",
37919 => "0110001110110000",
37920 => "0110001110110000",
37921 => "0110001110110000",
37922 => "0110001110110000",
37923 => "0110001110110000",
37924 => "0110001110110000",
37925 => "0110001110110000",
37926 => "0110001110110000",
37927 => "0110001110110000",
37928 => "0110001110110000",
37929 => "0110001110110000",
37930 => "0110001111000000",
37931 => "0110001111000000",
37932 => "0110001111000000",
37933 => "0110001111000000",
37934 => "0110001111000000",
37935 => "0110001111000000",
37936 => "0110001111000000",
37937 => "0110001111000000",
37938 => "0110001111000000",
37939 => "0110001111000000",
37940 => "0110001111000000",
37941 => "0110001111010000",
37942 => "0110001111010000",
37943 => "0110001111010000",
37944 => "0110001111010000",
37945 => "0110001111010000",
37946 => "0110001111010000",
37947 => "0110001111010000",
37948 => "0110001111010000",
37949 => "0110001111010000",
37950 => "0110001111010000",
37951 => "0110001111010000",
37952 => "0110001111010000",
37953 => "0110001111100000",
37954 => "0110001111100000",
37955 => "0110001111100000",
37956 => "0110001111100000",
37957 => "0110001111100000",
37958 => "0110001111100000",
37959 => "0110001111100000",
37960 => "0110001111100000",
37961 => "0110001111100000",
37962 => "0110001111100000",
37963 => "0110001111100000",
37964 => "0110001111110000",
37965 => "0110001111110000",
37966 => "0110001111110000",
37967 => "0110001111110000",
37968 => "0110001111110000",
37969 => "0110001111110000",
37970 => "0110001111110000",
37971 => "0110001111110000",
37972 => "0110001111110000",
37973 => "0110001111110000",
37974 => "0110001111110000",
37975 => "0110001111110000",
37976 => "0110010000000000",
37977 => "0110010000000000",
37978 => "0110010000000000",
37979 => "0110010000000000",
37980 => "0110010000000000",
37981 => "0110010000000000",
37982 => "0110010000000000",
37983 => "0110010000000000",
37984 => "0110010000000000",
37985 => "0110010000000000",
37986 => "0110010000000000",
37987 => "0110010000000000",
37988 => "0110010000010000",
37989 => "0110010000010000",
37990 => "0110010000010000",
37991 => "0110010000010000",
37992 => "0110010000010000",
37993 => "0110010000010000",
37994 => "0110010000010000",
37995 => "0110010000010000",
37996 => "0110010000010000",
37997 => "0110010000010000",
37998 => "0110010000010000",
37999 => "0110010000010000",
38000 => "0110010000100000",
38001 => "0110010000100000",
38002 => "0110010000100000",
38003 => "0110010000100000",
38004 => "0110010000100000",
38005 => "0110010000100000",
38006 => "0110010000100000",
38007 => "0110010000100000",
38008 => "0110010000100000",
38009 => "0110010000100000",
38010 => "0110010000100000",
38011 => "0110010000110000",
38012 => "0110010000110000",
38013 => "0110010000110000",
38014 => "0110010000110000",
38015 => "0110010000110000",
38016 => "0110010000110000",
38017 => "0110010000110000",
38018 => "0110010000110000",
38019 => "0110010000110000",
38020 => "0110010000110000",
38021 => "0110010000110000",
38022 => "0110010000110000",
38023 => "0110010001000000",
38024 => "0110010001000000",
38025 => "0110010001000000",
38026 => "0110010001000000",
38027 => "0110010001000000",
38028 => "0110010001000000",
38029 => "0110010001000000",
38030 => "0110010001000000",
38031 => "0110010001000000",
38032 => "0110010001000000",
38033 => "0110010001000000",
38034 => "0110010001000000",
38035 => "0110010001010000",
38036 => "0110010001010000",
38037 => "0110010001010000",
38038 => "0110010001010000",
38039 => "0110010001010000",
38040 => "0110010001010000",
38041 => "0110010001010000",
38042 => "0110010001010000",
38043 => "0110010001010000",
38044 => "0110010001010000",
38045 => "0110010001010000",
38046 => "0110010001010000",
38047 => "0110010001100000",
38048 => "0110010001100000",
38049 => "0110010001100000",
38050 => "0110010001100000",
38051 => "0110010001100000",
38052 => "0110010001100000",
38053 => "0110010001100000",
38054 => "0110010001100000",
38055 => "0110010001100000",
38056 => "0110010001100000",
38057 => "0110010001100000",
38058 => "0110010001110000",
38059 => "0110010001110000",
38060 => "0110010001110000",
38061 => "0110010001110000",
38062 => "0110010001110000",
38063 => "0110010001110000",
38064 => "0110010001110000",
38065 => "0110010001110000",
38066 => "0110010001110000",
38067 => "0110010001110000",
38068 => "0110010001110000",
38069 => "0110010001110000",
38070 => "0110010010000000",
38071 => "0110010010000000",
38072 => "0110010010000000",
38073 => "0110010010000000",
38074 => "0110010010000000",
38075 => "0110010010000000",
38076 => "0110010010000000",
38077 => "0110010010000000",
38078 => "0110010010000000",
38079 => "0110010010000000",
38080 => "0110010010000000",
38081 => "0110010010000000",
38082 => "0110010010010000",
38083 => "0110010010010000",
38084 => "0110010010010000",
38085 => "0110010010010000",
38086 => "0110010010010000",
38087 => "0110010010010000",
38088 => "0110010010010000",
38089 => "0110010010010000",
38090 => "0110010010010000",
38091 => "0110010010010000",
38092 => "0110010010010000",
38093 => "0110010010010000",
38094 => "0110010010100000",
38095 => "0110010010100000",
38096 => "0110010010100000",
38097 => "0110010010100000",
38098 => "0110010010100000",
38099 => "0110010010100000",
38100 => "0110010010100000",
38101 => "0110010010100000",
38102 => "0110010010100000",
38103 => "0110010010100000",
38104 => "0110010010100000",
38105 => "0110010010100000",
38106 => "0110010010110000",
38107 => "0110010010110000",
38108 => "0110010010110000",
38109 => "0110010010110000",
38110 => "0110010010110000",
38111 => "0110010010110000",
38112 => "0110010010110000",
38113 => "0110010010110000",
38114 => "0110010010110000",
38115 => "0110010010110000",
38116 => "0110010010110000",
38117 => "0110010010110000",
38118 => "0110010011000000",
38119 => "0110010011000000",
38120 => "0110010011000000",
38121 => "0110010011000000",
38122 => "0110010011000000",
38123 => "0110010011000000",
38124 => "0110010011000000",
38125 => "0110010011000000",
38126 => "0110010011000000",
38127 => "0110010011000000",
38128 => "0110010011000000",
38129 => "0110010011000000",
38130 => "0110010011010000",
38131 => "0110010011010000",
38132 => "0110010011010000",
38133 => "0110010011010000",
38134 => "0110010011010000",
38135 => "0110010011010000",
38136 => "0110010011010000",
38137 => "0110010011010000",
38138 => "0110010011010000",
38139 => "0110010011010000",
38140 => "0110010011010000",
38141 => "0110010011010000",
38142 => "0110010011100000",
38143 => "0110010011100000",
38144 => "0110010011100000",
38145 => "0110010011100000",
38146 => "0110010011100000",
38147 => "0110010011100000",
38148 => "0110010011100000",
38149 => "0110010011100000",
38150 => "0110010011100000",
38151 => "0110010011100000",
38152 => "0110010011100000",
38153 => "0110010011100000",
38154 => "0110010011110000",
38155 => "0110010011110000",
38156 => "0110010011110000",
38157 => "0110010011110000",
38158 => "0110010011110000",
38159 => "0110010011110000",
38160 => "0110010011110000",
38161 => "0110010011110000",
38162 => "0110010011110000",
38163 => "0110010011110000",
38164 => "0110010011110000",
38165 => "0110010011110000",
38166 => "0110010100000000",
38167 => "0110010100000000",
38168 => "0110010100000000",
38169 => "0110010100000000",
38170 => "0110010100000000",
38171 => "0110010100000000",
38172 => "0110010100000000",
38173 => "0110010100000000",
38174 => "0110010100000000",
38175 => "0110010100000000",
38176 => "0110010100000000",
38177 => "0110010100000000",
38178 => "0110010100010000",
38179 => "0110010100010000",
38180 => "0110010100010000",
38181 => "0110010100010000",
38182 => "0110010100010000",
38183 => "0110010100010000",
38184 => "0110010100010000",
38185 => "0110010100010000",
38186 => "0110010100010000",
38187 => "0110010100010000",
38188 => "0110010100010000",
38189 => "0110010100010000",
38190 => "0110010100100000",
38191 => "0110010100100000",
38192 => "0110010100100000",
38193 => "0110010100100000",
38194 => "0110010100100000",
38195 => "0110010100100000",
38196 => "0110010100100000",
38197 => "0110010100100000",
38198 => "0110010100100000",
38199 => "0110010100100000",
38200 => "0110010100100000",
38201 => "0110010100100000",
38202 => "0110010100110000",
38203 => "0110010100110000",
38204 => "0110010100110000",
38205 => "0110010100110000",
38206 => "0110010100110000",
38207 => "0110010100110000",
38208 => "0110010100110000",
38209 => "0110010100110000",
38210 => "0110010100110000",
38211 => "0110010100110000",
38212 => "0110010100110000",
38213 => "0110010100110000",
38214 => "0110010101000000",
38215 => "0110010101000000",
38216 => "0110010101000000",
38217 => "0110010101000000",
38218 => "0110010101000000",
38219 => "0110010101000000",
38220 => "0110010101000000",
38221 => "0110010101000000",
38222 => "0110010101000000",
38223 => "0110010101000000",
38224 => "0110010101000000",
38225 => "0110010101000000",
38226 => "0110010101010000",
38227 => "0110010101010000",
38228 => "0110010101010000",
38229 => "0110010101010000",
38230 => "0110010101010000",
38231 => "0110010101010000",
38232 => "0110010101010000",
38233 => "0110010101010000",
38234 => "0110010101010000",
38235 => "0110010101010000",
38236 => "0110010101010000",
38237 => "0110010101010000",
38238 => "0110010101100000",
38239 => "0110010101100000",
38240 => "0110010101100000",
38241 => "0110010101100000",
38242 => "0110010101100000",
38243 => "0110010101100000",
38244 => "0110010101100000",
38245 => "0110010101100000",
38246 => "0110010101100000",
38247 => "0110010101100000",
38248 => "0110010101100000",
38249 => "0110010101100000",
38250 => "0110010101110000",
38251 => "0110010101110000",
38252 => "0110010101110000",
38253 => "0110010101110000",
38254 => "0110010101110000",
38255 => "0110010101110000",
38256 => "0110010101110000",
38257 => "0110010101110000",
38258 => "0110010101110000",
38259 => "0110010101110000",
38260 => "0110010101110000",
38261 => "0110010101110000",
38262 => "0110010110000000",
38263 => "0110010110000000",
38264 => "0110010110000000",
38265 => "0110010110000000",
38266 => "0110010110000000",
38267 => "0110010110000000",
38268 => "0110010110000000",
38269 => "0110010110000000",
38270 => "0110010110000000",
38271 => "0110010110000000",
38272 => "0110010110000000",
38273 => "0110010110000000",
38274 => "0110010110000000",
38275 => "0110010110010000",
38276 => "0110010110010000",
38277 => "0110010110010000",
38278 => "0110010110010000",
38279 => "0110010110010000",
38280 => "0110010110010000",
38281 => "0110010110010000",
38282 => "0110010110010000",
38283 => "0110010110010000",
38284 => "0110010110010000",
38285 => "0110010110010000",
38286 => "0110010110010000",
38287 => "0110010110100000",
38288 => "0110010110100000",
38289 => "0110010110100000",
38290 => "0110010110100000",
38291 => "0110010110100000",
38292 => "0110010110100000",
38293 => "0110010110100000",
38294 => "0110010110100000",
38295 => "0110010110100000",
38296 => "0110010110100000",
38297 => "0110010110100000",
38298 => "0110010110100000",
38299 => "0110010110110000",
38300 => "0110010110110000",
38301 => "0110010110110000",
38302 => "0110010110110000",
38303 => "0110010110110000",
38304 => "0110010110110000",
38305 => "0110010110110000",
38306 => "0110010110110000",
38307 => "0110010110110000",
38308 => "0110010110110000",
38309 => "0110010110110000",
38310 => "0110010110110000",
38311 => "0110010111000000",
38312 => "0110010111000000",
38313 => "0110010111000000",
38314 => "0110010111000000",
38315 => "0110010111000000",
38316 => "0110010111000000",
38317 => "0110010111000000",
38318 => "0110010111000000",
38319 => "0110010111000000",
38320 => "0110010111000000",
38321 => "0110010111000000",
38322 => "0110010111000000",
38323 => "0110010111000000",
38324 => "0110010111010000",
38325 => "0110010111010000",
38326 => "0110010111010000",
38327 => "0110010111010000",
38328 => "0110010111010000",
38329 => "0110010111010000",
38330 => "0110010111010000",
38331 => "0110010111010000",
38332 => "0110010111010000",
38333 => "0110010111010000",
38334 => "0110010111010000",
38335 => "0110010111010000",
38336 => "0110010111100000",
38337 => "0110010111100000",
38338 => "0110010111100000",
38339 => "0110010111100000",
38340 => "0110010111100000",
38341 => "0110010111100000",
38342 => "0110010111100000",
38343 => "0110010111100000",
38344 => "0110010111100000",
38345 => "0110010111100000",
38346 => "0110010111100000",
38347 => "0110010111100000",
38348 => "0110010111110000",
38349 => "0110010111110000",
38350 => "0110010111110000",
38351 => "0110010111110000",
38352 => "0110010111110000",
38353 => "0110010111110000",
38354 => "0110010111110000",
38355 => "0110010111110000",
38356 => "0110010111110000",
38357 => "0110010111110000",
38358 => "0110010111110000",
38359 => "0110010111110000",
38360 => "0110011000000000",
38361 => "0110011000000000",
38362 => "0110011000000000",
38363 => "0110011000000000",
38364 => "0110011000000000",
38365 => "0110011000000000",
38366 => "0110011000000000",
38367 => "0110011000000000",
38368 => "0110011000000000",
38369 => "0110011000000000",
38370 => "0110011000000000",
38371 => "0110011000000000",
38372 => "0110011000000000",
38373 => "0110011000010000",
38374 => "0110011000010000",
38375 => "0110011000010000",
38376 => "0110011000010000",
38377 => "0110011000010000",
38378 => "0110011000010000",
38379 => "0110011000010000",
38380 => "0110011000010000",
38381 => "0110011000010000",
38382 => "0110011000010000",
38383 => "0110011000010000",
38384 => "0110011000010000",
38385 => "0110011000100000",
38386 => "0110011000100000",
38387 => "0110011000100000",
38388 => "0110011000100000",
38389 => "0110011000100000",
38390 => "0110011000100000",
38391 => "0110011000100000",
38392 => "0110011000100000",
38393 => "0110011000100000",
38394 => "0110011000100000",
38395 => "0110011000100000",
38396 => "0110011000100000",
38397 => "0110011000100000",
38398 => "0110011000110000",
38399 => "0110011000110000",
38400 => "0110011000110000",
38401 => "0110011000110000",
38402 => "0110011000110000",
38403 => "0110011000110000",
38404 => "0110011000110000",
38405 => "0110011000110000",
38406 => "0110011000110000",
38407 => "0110011000110000",
38408 => "0110011000110000",
38409 => "0110011000110000",
38410 => "0110011001000000",
38411 => "0110011001000000",
38412 => "0110011001000000",
38413 => "0110011001000000",
38414 => "0110011001000000",
38415 => "0110011001000000",
38416 => "0110011001000000",
38417 => "0110011001000000",
38418 => "0110011001000000",
38419 => "0110011001000000",
38420 => "0110011001000000",
38421 => "0110011001000000",
38422 => "0110011001010000",
38423 => "0110011001010000",
38424 => "0110011001010000",
38425 => "0110011001010000",
38426 => "0110011001010000",
38427 => "0110011001010000",
38428 => "0110011001010000",
38429 => "0110011001010000",
38430 => "0110011001010000",
38431 => "0110011001010000",
38432 => "0110011001010000",
38433 => "0110011001010000",
38434 => "0110011001010000",
38435 => "0110011001100000",
38436 => "0110011001100000",
38437 => "0110011001100000",
38438 => "0110011001100000",
38439 => "0110011001100000",
38440 => "0110011001100000",
38441 => "0110011001100000",
38442 => "0110011001100000",
38443 => "0110011001100000",
38444 => "0110011001100000",
38445 => "0110011001100000",
38446 => "0110011001100000",
38447 => "0110011001110000",
38448 => "0110011001110000",
38449 => "0110011001110000",
38450 => "0110011001110000",
38451 => "0110011001110000",
38452 => "0110011001110000",
38453 => "0110011001110000",
38454 => "0110011001110000",
38455 => "0110011001110000",
38456 => "0110011001110000",
38457 => "0110011001110000",
38458 => "0110011001110000",
38459 => "0110011001110000",
38460 => "0110011010000000",
38461 => "0110011010000000",
38462 => "0110011010000000",
38463 => "0110011010000000",
38464 => "0110011010000000",
38465 => "0110011010000000",
38466 => "0110011010000000",
38467 => "0110011010000000",
38468 => "0110011010000000",
38469 => "0110011010000000",
38470 => "0110011010000000",
38471 => "0110011010000000",
38472 => "0110011010010000",
38473 => "0110011010010000",
38474 => "0110011010010000",
38475 => "0110011010010000",
38476 => "0110011010010000",
38477 => "0110011010010000",
38478 => "0110011010010000",
38479 => "0110011010010000",
38480 => "0110011010010000",
38481 => "0110011010010000",
38482 => "0110011010010000",
38483 => "0110011010010000",
38484 => "0110011010010000",
38485 => "0110011010100000",
38486 => "0110011010100000",
38487 => "0110011010100000",
38488 => "0110011010100000",
38489 => "0110011010100000",
38490 => "0110011010100000",
38491 => "0110011010100000",
38492 => "0110011010100000",
38493 => "0110011010100000",
38494 => "0110011010100000",
38495 => "0110011010100000",
38496 => "0110011010100000",
38497 => "0110011010100000",
38498 => "0110011010110000",
38499 => "0110011010110000",
38500 => "0110011010110000",
38501 => "0110011010110000",
38502 => "0110011010110000",
38503 => "0110011010110000",
38504 => "0110011010110000",
38505 => "0110011010110000",
38506 => "0110011010110000",
38507 => "0110011010110000",
38508 => "0110011010110000",
38509 => "0110011010110000",
38510 => "0110011011000000",
38511 => "0110011011000000",
38512 => "0110011011000000",
38513 => "0110011011000000",
38514 => "0110011011000000",
38515 => "0110011011000000",
38516 => "0110011011000000",
38517 => "0110011011000000",
38518 => "0110011011000000",
38519 => "0110011011000000",
38520 => "0110011011000000",
38521 => "0110011011000000",
38522 => "0110011011000000",
38523 => "0110011011010000",
38524 => "0110011011010000",
38525 => "0110011011010000",
38526 => "0110011011010000",
38527 => "0110011011010000",
38528 => "0110011011010000",
38529 => "0110011011010000",
38530 => "0110011011010000",
38531 => "0110011011010000",
38532 => "0110011011010000",
38533 => "0110011011010000",
38534 => "0110011011010000",
38535 => "0110011011010000",
38536 => "0110011011100000",
38537 => "0110011011100000",
38538 => "0110011011100000",
38539 => "0110011011100000",
38540 => "0110011011100000",
38541 => "0110011011100000",
38542 => "0110011011100000",
38543 => "0110011011100000",
38544 => "0110011011100000",
38545 => "0110011011100000",
38546 => "0110011011100000",
38547 => "0110011011100000",
38548 => "0110011011110000",
38549 => "0110011011110000",
38550 => "0110011011110000",
38551 => "0110011011110000",
38552 => "0110011011110000",
38553 => "0110011011110000",
38554 => "0110011011110000",
38555 => "0110011011110000",
38556 => "0110011011110000",
38557 => "0110011011110000",
38558 => "0110011011110000",
38559 => "0110011011110000",
38560 => "0110011011110000",
38561 => "0110011100000000",
38562 => "0110011100000000",
38563 => "0110011100000000",
38564 => "0110011100000000",
38565 => "0110011100000000",
38566 => "0110011100000000",
38567 => "0110011100000000",
38568 => "0110011100000000",
38569 => "0110011100000000",
38570 => "0110011100000000",
38571 => "0110011100000000",
38572 => "0110011100000000",
38573 => "0110011100000000",
38574 => "0110011100010000",
38575 => "0110011100010000",
38576 => "0110011100010000",
38577 => "0110011100010000",
38578 => "0110011100010000",
38579 => "0110011100010000",
38580 => "0110011100010000",
38581 => "0110011100010000",
38582 => "0110011100010000",
38583 => "0110011100010000",
38584 => "0110011100010000",
38585 => "0110011100010000",
38586 => "0110011100100000",
38587 => "0110011100100000",
38588 => "0110011100100000",
38589 => "0110011100100000",
38590 => "0110011100100000",
38591 => "0110011100100000",
38592 => "0110011100100000",
38593 => "0110011100100000",
38594 => "0110011100100000",
38595 => "0110011100100000",
38596 => "0110011100100000",
38597 => "0110011100100000",
38598 => "0110011100100000",
38599 => "0110011100110000",
38600 => "0110011100110000",
38601 => "0110011100110000",
38602 => "0110011100110000",
38603 => "0110011100110000",
38604 => "0110011100110000",
38605 => "0110011100110000",
38606 => "0110011100110000",
38607 => "0110011100110000",
38608 => "0110011100110000",
38609 => "0110011100110000",
38610 => "0110011100110000",
38611 => "0110011100110000",
38612 => "0110011101000000",
38613 => "0110011101000000",
38614 => "0110011101000000",
38615 => "0110011101000000",
38616 => "0110011101000000",
38617 => "0110011101000000",
38618 => "0110011101000000",
38619 => "0110011101000000",
38620 => "0110011101000000",
38621 => "0110011101000000",
38622 => "0110011101000000",
38623 => "0110011101000000",
38624 => "0110011101000000",
38625 => "0110011101010000",
38626 => "0110011101010000",
38627 => "0110011101010000",
38628 => "0110011101010000",
38629 => "0110011101010000",
38630 => "0110011101010000",
38631 => "0110011101010000",
38632 => "0110011101010000",
38633 => "0110011101010000",
38634 => "0110011101010000",
38635 => "0110011101010000",
38636 => "0110011101010000",
38637 => "0110011101010000",
38638 => "0110011101100000",
38639 => "0110011101100000",
38640 => "0110011101100000",
38641 => "0110011101100000",
38642 => "0110011101100000",
38643 => "0110011101100000",
38644 => "0110011101100000",
38645 => "0110011101100000",
38646 => "0110011101100000",
38647 => "0110011101100000",
38648 => "0110011101100000",
38649 => "0110011101100000",
38650 => "0110011101110000",
38651 => "0110011101110000",
38652 => "0110011101110000",
38653 => "0110011101110000",
38654 => "0110011101110000",
38655 => "0110011101110000",
38656 => "0110011101110000",
38657 => "0110011101110000",
38658 => "0110011101110000",
38659 => "0110011101110000",
38660 => "0110011101110000",
38661 => "0110011101110000",
38662 => "0110011101110000",
38663 => "0110011110000000",
38664 => "0110011110000000",
38665 => "0110011110000000",
38666 => "0110011110000000",
38667 => "0110011110000000",
38668 => "0110011110000000",
38669 => "0110011110000000",
38670 => "0110011110000000",
38671 => "0110011110000000",
38672 => "0110011110000000",
38673 => "0110011110000000",
38674 => "0110011110000000",
38675 => "0110011110000000",
38676 => "0110011110010000",
38677 => "0110011110010000",
38678 => "0110011110010000",
38679 => "0110011110010000",
38680 => "0110011110010000",
38681 => "0110011110010000",
38682 => "0110011110010000",
38683 => "0110011110010000",
38684 => "0110011110010000",
38685 => "0110011110010000",
38686 => "0110011110010000",
38687 => "0110011110010000",
38688 => "0110011110010000",
38689 => "0110011110100000",
38690 => "0110011110100000",
38691 => "0110011110100000",
38692 => "0110011110100000",
38693 => "0110011110100000",
38694 => "0110011110100000",
38695 => "0110011110100000",
38696 => "0110011110100000",
38697 => "0110011110100000",
38698 => "0110011110100000",
38699 => "0110011110100000",
38700 => "0110011110100000",
38701 => "0110011110100000",
38702 => "0110011110110000",
38703 => "0110011110110000",
38704 => "0110011110110000",
38705 => "0110011110110000",
38706 => "0110011110110000",
38707 => "0110011110110000",
38708 => "0110011110110000",
38709 => "0110011110110000",
38710 => "0110011110110000",
38711 => "0110011110110000",
38712 => "0110011110110000",
38713 => "0110011110110000",
38714 => "0110011110110000",
38715 => "0110011111000000",
38716 => "0110011111000000",
38717 => "0110011111000000",
38718 => "0110011111000000",
38719 => "0110011111000000",
38720 => "0110011111000000",
38721 => "0110011111000000",
38722 => "0110011111000000",
38723 => "0110011111000000",
38724 => "0110011111000000",
38725 => "0110011111000000",
38726 => "0110011111000000",
38727 => "0110011111000000",
38728 => "0110011111010000",
38729 => "0110011111010000",
38730 => "0110011111010000",
38731 => "0110011111010000",
38732 => "0110011111010000",
38733 => "0110011111010000",
38734 => "0110011111010000",
38735 => "0110011111010000",
38736 => "0110011111010000",
38737 => "0110011111010000",
38738 => "0110011111010000",
38739 => "0110011111010000",
38740 => "0110011111010000",
38741 => "0110011111100000",
38742 => "0110011111100000",
38743 => "0110011111100000",
38744 => "0110011111100000",
38745 => "0110011111100000",
38746 => "0110011111100000",
38747 => "0110011111100000",
38748 => "0110011111100000",
38749 => "0110011111100000",
38750 => "0110011111100000",
38751 => "0110011111100000",
38752 => "0110011111100000",
38753 => "0110011111100000",
38754 => "0110011111110000",
38755 => "0110011111110000",
38756 => "0110011111110000",
38757 => "0110011111110000",
38758 => "0110011111110000",
38759 => "0110011111110000",
38760 => "0110011111110000",
38761 => "0110011111110000",
38762 => "0110011111110000",
38763 => "0110011111110000",
38764 => "0110011111110000",
38765 => "0110011111110000",
38766 => "0110011111110000",
38767 => "0110100000000000",
38768 => "0110100000000000",
38769 => "0110100000000000",
38770 => "0110100000000000",
38771 => "0110100000000000",
38772 => "0110100000000000",
38773 => "0110100000000000",
38774 => "0110100000000000",
38775 => "0110100000000000",
38776 => "0110100000000000",
38777 => "0110100000000000",
38778 => "0110100000000000",
38779 => "0110100000000000",
38780 => "0110100000000000",
38781 => "0110100000010000",
38782 => "0110100000010000",
38783 => "0110100000010000",
38784 => "0110100000010000",
38785 => "0110100000010000",
38786 => "0110100000010000",
38787 => "0110100000010000",
38788 => "0110100000010000",
38789 => "0110100000010000",
38790 => "0110100000010000",
38791 => "0110100000010000",
38792 => "0110100000010000",
38793 => "0110100000010000",
38794 => "0110100000100000",
38795 => "0110100000100000",
38796 => "0110100000100000",
38797 => "0110100000100000",
38798 => "0110100000100000",
38799 => "0110100000100000",
38800 => "0110100000100000",
38801 => "0110100000100000",
38802 => "0110100000100000",
38803 => "0110100000100000",
38804 => "0110100000100000",
38805 => "0110100000100000",
38806 => "0110100000100000",
38807 => "0110100000110000",
38808 => "0110100000110000",
38809 => "0110100000110000",
38810 => "0110100000110000",
38811 => "0110100000110000",
38812 => "0110100000110000",
38813 => "0110100000110000",
38814 => "0110100000110000",
38815 => "0110100000110000",
38816 => "0110100000110000",
38817 => "0110100000110000",
38818 => "0110100000110000",
38819 => "0110100000110000",
38820 => "0110100001000000",
38821 => "0110100001000000",
38822 => "0110100001000000",
38823 => "0110100001000000",
38824 => "0110100001000000",
38825 => "0110100001000000",
38826 => "0110100001000000",
38827 => "0110100001000000",
38828 => "0110100001000000",
38829 => "0110100001000000",
38830 => "0110100001000000",
38831 => "0110100001000000",
38832 => "0110100001000000",
38833 => "0110100001010000",
38834 => "0110100001010000",
38835 => "0110100001010000",
38836 => "0110100001010000",
38837 => "0110100001010000",
38838 => "0110100001010000",
38839 => "0110100001010000",
38840 => "0110100001010000",
38841 => "0110100001010000",
38842 => "0110100001010000",
38843 => "0110100001010000",
38844 => "0110100001010000",
38845 => "0110100001010000",
38846 => "0110100001010000",
38847 => "0110100001100000",
38848 => "0110100001100000",
38849 => "0110100001100000",
38850 => "0110100001100000",
38851 => "0110100001100000",
38852 => "0110100001100000",
38853 => "0110100001100000",
38854 => "0110100001100000",
38855 => "0110100001100000",
38856 => "0110100001100000",
38857 => "0110100001100000",
38858 => "0110100001100000",
38859 => "0110100001100000",
38860 => "0110100001110000",
38861 => "0110100001110000",
38862 => "0110100001110000",
38863 => "0110100001110000",
38864 => "0110100001110000",
38865 => "0110100001110000",
38866 => "0110100001110000",
38867 => "0110100001110000",
38868 => "0110100001110000",
38869 => "0110100001110000",
38870 => "0110100001110000",
38871 => "0110100001110000",
38872 => "0110100001110000",
38873 => "0110100010000000",
38874 => "0110100010000000",
38875 => "0110100010000000",
38876 => "0110100010000000",
38877 => "0110100010000000",
38878 => "0110100010000000",
38879 => "0110100010000000",
38880 => "0110100010000000",
38881 => "0110100010000000",
38882 => "0110100010000000",
38883 => "0110100010000000",
38884 => "0110100010000000",
38885 => "0110100010000000",
38886 => "0110100010000000",
38887 => "0110100010010000",
38888 => "0110100010010000",
38889 => "0110100010010000",
38890 => "0110100010010000",
38891 => "0110100010010000",
38892 => "0110100010010000",
38893 => "0110100010010000",
38894 => "0110100010010000",
38895 => "0110100010010000",
38896 => "0110100010010000",
38897 => "0110100010010000",
38898 => "0110100010010000",
38899 => "0110100010010000",
38900 => "0110100010100000",
38901 => "0110100010100000",
38902 => "0110100010100000",
38903 => "0110100010100000",
38904 => "0110100010100000",
38905 => "0110100010100000",
38906 => "0110100010100000",
38907 => "0110100010100000",
38908 => "0110100010100000",
38909 => "0110100010100000",
38910 => "0110100010100000",
38911 => "0110100010100000",
38912 => "0110100010100000",
38913 => "0110100010110000",
38914 => "0110100010110000",
38915 => "0110100010110000",
38916 => "0110100010110000",
38917 => "0110100010110000",
38918 => "0110100010110000",
38919 => "0110100010110000",
38920 => "0110100010110000",
38921 => "0110100010110000",
38922 => "0110100010110000",
38923 => "0110100010110000",
38924 => "0110100010110000",
38925 => "0110100010110000",
38926 => "0110100010110000",
38927 => "0110100011000000",
38928 => "0110100011000000",
38929 => "0110100011000000",
38930 => "0110100011000000",
38931 => "0110100011000000",
38932 => "0110100011000000",
38933 => "0110100011000000",
38934 => "0110100011000000",
38935 => "0110100011000000",
38936 => "0110100011000000",
38937 => "0110100011000000",
38938 => "0110100011000000",
38939 => "0110100011000000",
38940 => "0110100011010000",
38941 => "0110100011010000",
38942 => "0110100011010000",
38943 => "0110100011010000",
38944 => "0110100011010000",
38945 => "0110100011010000",
38946 => "0110100011010000",
38947 => "0110100011010000",
38948 => "0110100011010000",
38949 => "0110100011010000",
38950 => "0110100011010000",
38951 => "0110100011010000",
38952 => "0110100011010000",
38953 => "0110100011010000",
38954 => "0110100011100000",
38955 => "0110100011100000",
38956 => "0110100011100000",
38957 => "0110100011100000",
38958 => "0110100011100000",
38959 => "0110100011100000",
38960 => "0110100011100000",
38961 => "0110100011100000",
38962 => "0110100011100000",
38963 => "0110100011100000",
38964 => "0110100011100000",
38965 => "0110100011100000",
38966 => "0110100011100000",
38967 => "0110100011110000",
38968 => "0110100011110000",
38969 => "0110100011110000",
38970 => "0110100011110000",
38971 => "0110100011110000",
38972 => "0110100011110000",
38973 => "0110100011110000",
38974 => "0110100011110000",
38975 => "0110100011110000",
38976 => "0110100011110000",
38977 => "0110100011110000",
38978 => "0110100011110000",
38979 => "0110100011110000",
38980 => "0110100011110000",
38981 => "0110100100000000",
38982 => "0110100100000000",
38983 => "0110100100000000",
38984 => "0110100100000000",
38985 => "0110100100000000",
38986 => "0110100100000000",
38987 => "0110100100000000",
38988 => "0110100100000000",
38989 => "0110100100000000",
38990 => "0110100100000000",
38991 => "0110100100000000",
38992 => "0110100100000000",
38993 => "0110100100000000",
38994 => "0110100100010000",
38995 => "0110100100010000",
38996 => "0110100100010000",
38997 => "0110100100010000",
38998 => "0110100100010000",
38999 => "0110100100010000",
39000 => "0110100100010000",
39001 => "0110100100010000",
39002 => "0110100100010000",
39003 => "0110100100010000",
39004 => "0110100100010000",
39005 => "0110100100010000",
39006 => "0110100100010000",
39007 => "0110100100010000",
39008 => "0110100100100000",
39009 => "0110100100100000",
39010 => "0110100100100000",
39011 => "0110100100100000",
39012 => "0110100100100000",
39013 => "0110100100100000",
39014 => "0110100100100000",
39015 => "0110100100100000",
39016 => "0110100100100000",
39017 => "0110100100100000",
39018 => "0110100100100000",
39019 => "0110100100100000",
39020 => "0110100100100000",
39021 => "0110100100100000",
39022 => "0110100100110000",
39023 => "0110100100110000",
39024 => "0110100100110000",
39025 => "0110100100110000",
39026 => "0110100100110000",
39027 => "0110100100110000",
39028 => "0110100100110000",
39029 => "0110100100110000",
39030 => "0110100100110000",
39031 => "0110100100110000",
39032 => "0110100100110000",
39033 => "0110100100110000",
39034 => "0110100100110000",
39035 => "0110100101000000",
39036 => "0110100101000000",
39037 => "0110100101000000",
39038 => "0110100101000000",
39039 => "0110100101000000",
39040 => "0110100101000000",
39041 => "0110100101000000",
39042 => "0110100101000000",
39043 => "0110100101000000",
39044 => "0110100101000000",
39045 => "0110100101000000",
39046 => "0110100101000000",
39047 => "0110100101000000",
39048 => "0110100101000000",
39049 => "0110100101010000",
39050 => "0110100101010000",
39051 => "0110100101010000",
39052 => "0110100101010000",
39053 => "0110100101010000",
39054 => "0110100101010000",
39055 => "0110100101010000",
39056 => "0110100101010000",
39057 => "0110100101010000",
39058 => "0110100101010000",
39059 => "0110100101010000",
39060 => "0110100101010000",
39061 => "0110100101010000",
39062 => "0110100101010000",
39063 => "0110100101100000",
39064 => "0110100101100000",
39065 => "0110100101100000",
39066 => "0110100101100000",
39067 => "0110100101100000",
39068 => "0110100101100000",
39069 => "0110100101100000",
39070 => "0110100101100000",
39071 => "0110100101100000",
39072 => "0110100101100000",
39073 => "0110100101100000",
39074 => "0110100101100000",
39075 => "0110100101100000",
39076 => "0110100101110000",
39077 => "0110100101110000",
39078 => "0110100101110000",
39079 => "0110100101110000",
39080 => "0110100101110000",
39081 => "0110100101110000",
39082 => "0110100101110000",
39083 => "0110100101110000",
39084 => "0110100101110000",
39085 => "0110100101110000",
39086 => "0110100101110000",
39087 => "0110100101110000",
39088 => "0110100101110000",
39089 => "0110100101110000",
39090 => "0110100110000000",
39091 => "0110100110000000",
39092 => "0110100110000000",
39093 => "0110100110000000",
39094 => "0110100110000000",
39095 => "0110100110000000",
39096 => "0110100110000000",
39097 => "0110100110000000",
39098 => "0110100110000000",
39099 => "0110100110000000",
39100 => "0110100110000000",
39101 => "0110100110000000",
39102 => "0110100110000000",
39103 => "0110100110000000",
39104 => "0110100110010000",
39105 => "0110100110010000",
39106 => "0110100110010000",
39107 => "0110100110010000",
39108 => "0110100110010000",
39109 => "0110100110010000",
39110 => "0110100110010000",
39111 => "0110100110010000",
39112 => "0110100110010000",
39113 => "0110100110010000",
39114 => "0110100110010000",
39115 => "0110100110010000",
39116 => "0110100110010000",
39117 => "0110100110010000",
39118 => "0110100110100000",
39119 => "0110100110100000",
39120 => "0110100110100000",
39121 => "0110100110100000",
39122 => "0110100110100000",
39123 => "0110100110100000",
39124 => "0110100110100000",
39125 => "0110100110100000",
39126 => "0110100110100000",
39127 => "0110100110100000",
39128 => "0110100110100000",
39129 => "0110100110100000",
39130 => "0110100110100000",
39131 => "0110100110100000",
39132 => "0110100110110000",
39133 => "0110100110110000",
39134 => "0110100110110000",
39135 => "0110100110110000",
39136 => "0110100110110000",
39137 => "0110100110110000",
39138 => "0110100110110000",
39139 => "0110100110110000",
39140 => "0110100110110000",
39141 => "0110100110110000",
39142 => "0110100110110000",
39143 => "0110100110110000",
39144 => "0110100110110000",
39145 => "0110100110110000",
39146 => "0110100111000000",
39147 => "0110100111000000",
39148 => "0110100111000000",
39149 => "0110100111000000",
39150 => "0110100111000000",
39151 => "0110100111000000",
39152 => "0110100111000000",
39153 => "0110100111000000",
39154 => "0110100111000000",
39155 => "0110100111000000",
39156 => "0110100111000000",
39157 => "0110100111000000",
39158 => "0110100111000000",
39159 => "0110100111010000",
39160 => "0110100111010000",
39161 => "0110100111010000",
39162 => "0110100111010000",
39163 => "0110100111010000",
39164 => "0110100111010000",
39165 => "0110100111010000",
39166 => "0110100111010000",
39167 => "0110100111010000",
39168 => "0110100111010000",
39169 => "0110100111010000",
39170 => "0110100111010000",
39171 => "0110100111010000",
39172 => "0110100111010000",
39173 => "0110100111100000",
39174 => "0110100111100000",
39175 => "0110100111100000",
39176 => "0110100111100000",
39177 => "0110100111100000",
39178 => "0110100111100000",
39179 => "0110100111100000",
39180 => "0110100111100000",
39181 => "0110100111100000",
39182 => "0110100111100000",
39183 => "0110100111100000",
39184 => "0110100111100000",
39185 => "0110100111100000",
39186 => "0110100111100000",
39187 => "0110100111110000",
39188 => "0110100111110000",
39189 => "0110100111110000",
39190 => "0110100111110000",
39191 => "0110100111110000",
39192 => "0110100111110000",
39193 => "0110100111110000",
39194 => "0110100111110000",
39195 => "0110100111110000",
39196 => "0110100111110000",
39197 => "0110100111110000",
39198 => "0110100111110000",
39199 => "0110100111110000",
39200 => "0110100111110000",
39201 => "0110101000000000",
39202 => "0110101000000000",
39203 => "0110101000000000",
39204 => "0110101000000000",
39205 => "0110101000000000",
39206 => "0110101000000000",
39207 => "0110101000000000",
39208 => "0110101000000000",
39209 => "0110101000000000",
39210 => "0110101000000000",
39211 => "0110101000000000",
39212 => "0110101000000000",
39213 => "0110101000000000",
39214 => "0110101000000000",
39215 => "0110101000010000",
39216 => "0110101000010000",
39217 => "0110101000010000",
39218 => "0110101000010000",
39219 => "0110101000010000",
39220 => "0110101000010000",
39221 => "0110101000010000",
39222 => "0110101000010000",
39223 => "0110101000010000",
39224 => "0110101000010000",
39225 => "0110101000010000",
39226 => "0110101000010000",
39227 => "0110101000010000",
39228 => "0110101000010000",
39229 => "0110101000010000",
39230 => "0110101000100000",
39231 => "0110101000100000",
39232 => "0110101000100000",
39233 => "0110101000100000",
39234 => "0110101000100000",
39235 => "0110101000100000",
39236 => "0110101000100000",
39237 => "0110101000100000",
39238 => "0110101000100000",
39239 => "0110101000100000",
39240 => "0110101000100000",
39241 => "0110101000100000",
39242 => "0110101000100000",
39243 => "0110101000100000",
39244 => "0110101000110000",
39245 => "0110101000110000",
39246 => "0110101000110000",
39247 => "0110101000110000",
39248 => "0110101000110000",
39249 => "0110101000110000",
39250 => "0110101000110000",
39251 => "0110101000110000",
39252 => "0110101000110000",
39253 => "0110101000110000",
39254 => "0110101000110000",
39255 => "0110101000110000",
39256 => "0110101000110000",
39257 => "0110101000110000",
39258 => "0110101001000000",
39259 => "0110101001000000",
39260 => "0110101001000000",
39261 => "0110101001000000",
39262 => "0110101001000000",
39263 => "0110101001000000",
39264 => "0110101001000000",
39265 => "0110101001000000",
39266 => "0110101001000000",
39267 => "0110101001000000",
39268 => "0110101001000000",
39269 => "0110101001000000",
39270 => "0110101001000000",
39271 => "0110101001000000",
39272 => "0110101001010000",
39273 => "0110101001010000",
39274 => "0110101001010000",
39275 => "0110101001010000",
39276 => "0110101001010000",
39277 => "0110101001010000",
39278 => "0110101001010000",
39279 => "0110101001010000",
39280 => "0110101001010000",
39281 => "0110101001010000",
39282 => "0110101001010000",
39283 => "0110101001010000",
39284 => "0110101001010000",
39285 => "0110101001010000",
39286 => "0110101001100000",
39287 => "0110101001100000",
39288 => "0110101001100000",
39289 => "0110101001100000",
39290 => "0110101001100000",
39291 => "0110101001100000",
39292 => "0110101001100000",
39293 => "0110101001100000",
39294 => "0110101001100000",
39295 => "0110101001100000",
39296 => "0110101001100000",
39297 => "0110101001100000",
39298 => "0110101001100000",
39299 => "0110101001100000",
39300 => "0110101001110000",
39301 => "0110101001110000",
39302 => "0110101001110000",
39303 => "0110101001110000",
39304 => "0110101001110000",
39305 => "0110101001110000",
39306 => "0110101001110000",
39307 => "0110101001110000",
39308 => "0110101001110000",
39309 => "0110101001110000",
39310 => "0110101001110000",
39311 => "0110101001110000",
39312 => "0110101001110000",
39313 => "0110101001110000",
39314 => "0110101001110000",
39315 => "0110101010000000",
39316 => "0110101010000000",
39317 => "0110101010000000",
39318 => "0110101010000000",
39319 => "0110101010000000",
39320 => "0110101010000000",
39321 => "0110101010000000",
39322 => "0110101010000000",
39323 => "0110101010000000",
39324 => "0110101010000000",
39325 => "0110101010000000",
39326 => "0110101010000000",
39327 => "0110101010000000",
39328 => "0110101010000000",
39329 => "0110101010010000",
39330 => "0110101010010000",
39331 => "0110101010010000",
39332 => "0110101010010000",
39333 => "0110101010010000",
39334 => "0110101010010000",
39335 => "0110101010010000",
39336 => "0110101010010000",
39337 => "0110101010010000",
39338 => "0110101010010000",
39339 => "0110101010010000",
39340 => "0110101010010000",
39341 => "0110101010010000",
39342 => "0110101010010000",
39343 => "0110101010100000",
39344 => "0110101010100000",
39345 => "0110101010100000",
39346 => "0110101010100000",
39347 => "0110101010100000",
39348 => "0110101010100000",
39349 => "0110101010100000",
39350 => "0110101010100000",
39351 => "0110101010100000",
39352 => "0110101010100000",
39353 => "0110101010100000",
39354 => "0110101010100000",
39355 => "0110101010100000",
39356 => "0110101010100000",
39357 => "0110101010100000",
39358 => "0110101010110000",
39359 => "0110101010110000",
39360 => "0110101010110000",
39361 => "0110101010110000",
39362 => "0110101010110000",
39363 => "0110101010110000",
39364 => "0110101010110000",
39365 => "0110101010110000",
39366 => "0110101010110000",
39367 => "0110101010110000",
39368 => "0110101010110000",
39369 => "0110101010110000",
39370 => "0110101010110000",
39371 => "0110101010110000",
39372 => "0110101011000000",
39373 => "0110101011000000",
39374 => "0110101011000000",
39375 => "0110101011000000",
39376 => "0110101011000000",
39377 => "0110101011000000",
39378 => "0110101011000000",
39379 => "0110101011000000",
39380 => "0110101011000000",
39381 => "0110101011000000",
39382 => "0110101011000000",
39383 => "0110101011000000",
39384 => "0110101011000000",
39385 => "0110101011000000",
39386 => "0110101011000000",
39387 => "0110101011010000",
39388 => "0110101011010000",
39389 => "0110101011010000",
39390 => "0110101011010000",
39391 => "0110101011010000",
39392 => "0110101011010000",
39393 => "0110101011010000",
39394 => "0110101011010000",
39395 => "0110101011010000",
39396 => "0110101011010000",
39397 => "0110101011010000",
39398 => "0110101011010000",
39399 => "0110101011010000",
39400 => "0110101011010000",
39401 => "0110101011100000",
39402 => "0110101011100000",
39403 => "0110101011100000",
39404 => "0110101011100000",
39405 => "0110101011100000",
39406 => "0110101011100000",
39407 => "0110101011100000",
39408 => "0110101011100000",
39409 => "0110101011100000",
39410 => "0110101011100000",
39411 => "0110101011100000",
39412 => "0110101011100000",
39413 => "0110101011100000",
39414 => "0110101011100000",
39415 => "0110101011100000",
39416 => "0110101011110000",
39417 => "0110101011110000",
39418 => "0110101011110000",
39419 => "0110101011110000",
39420 => "0110101011110000",
39421 => "0110101011110000",
39422 => "0110101011110000",
39423 => "0110101011110000",
39424 => "0110101011110000",
39425 => "0110101011110000",
39426 => "0110101011110000",
39427 => "0110101011110000",
39428 => "0110101011110000",
39429 => "0110101011110000",
39430 => "0110101100000000",
39431 => "0110101100000000",
39432 => "0110101100000000",
39433 => "0110101100000000",
39434 => "0110101100000000",
39435 => "0110101100000000",
39436 => "0110101100000000",
39437 => "0110101100000000",
39438 => "0110101100000000",
39439 => "0110101100000000",
39440 => "0110101100000000",
39441 => "0110101100000000",
39442 => "0110101100000000",
39443 => "0110101100000000",
39444 => "0110101100000000",
39445 => "0110101100010000",
39446 => "0110101100010000",
39447 => "0110101100010000",
39448 => "0110101100010000",
39449 => "0110101100010000",
39450 => "0110101100010000",
39451 => "0110101100010000",
39452 => "0110101100010000",
39453 => "0110101100010000",
39454 => "0110101100010000",
39455 => "0110101100010000",
39456 => "0110101100010000",
39457 => "0110101100010000",
39458 => "0110101100010000",
39459 => "0110101100100000",
39460 => "0110101100100000",
39461 => "0110101100100000",
39462 => "0110101100100000",
39463 => "0110101100100000",
39464 => "0110101100100000",
39465 => "0110101100100000",
39466 => "0110101100100000",
39467 => "0110101100100000",
39468 => "0110101100100000",
39469 => "0110101100100000",
39470 => "0110101100100000",
39471 => "0110101100100000",
39472 => "0110101100100000",
39473 => "0110101100100000",
39474 => "0110101100110000",
39475 => "0110101100110000",
39476 => "0110101100110000",
39477 => "0110101100110000",
39478 => "0110101100110000",
39479 => "0110101100110000",
39480 => "0110101100110000",
39481 => "0110101100110000",
39482 => "0110101100110000",
39483 => "0110101100110000",
39484 => "0110101100110000",
39485 => "0110101100110000",
39486 => "0110101100110000",
39487 => "0110101100110000",
39488 => "0110101100110000",
39489 => "0110101101000000",
39490 => "0110101101000000",
39491 => "0110101101000000",
39492 => "0110101101000000",
39493 => "0110101101000000",
39494 => "0110101101000000",
39495 => "0110101101000000",
39496 => "0110101101000000",
39497 => "0110101101000000",
39498 => "0110101101000000",
39499 => "0110101101000000",
39500 => "0110101101000000",
39501 => "0110101101000000",
39502 => "0110101101000000",
39503 => "0110101101010000",
39504 => "0110101101010000",
39505 => "0110101101010000",
39506 => "0110101101010000",
39507 => "0110101101010000",
39508 => "0110101101010000",
39509 => "0110101101010000",
39510 => "0110101101010000",
39511 => "0110101101010000",
39512 => "0110101101010000",
39513 => "0110101101010000",
39514 => "0110101101010000",
39515 => "0110101101010000",
39516 => "0110101101010000",
39517 => "0110101101010000",
39518 => "0110101101100000",
39519 => "0110101101100000",
39520 => "0110101101100000",
39521 => "0110101101100000",
39522 => "0110101101100000",
39523 => "0110101101100000",
39524 => "0110101101100000",
39525 => "0110101101100000",
39526 => "0110101101100000",
39527 => "0110101101100000",
39528 => "0110101101100000",
39529 => "0110101101100000",
39530 => "0110101101100000",
39531 => "0110101101100000",
39532 => "0110101101100000",
39533 => "0110101101110000",
39534 => "0110101101110000",
39535 => "0110101101110000",
39536 => "0110101101110000",
39537 => "0110101101110000",
39538 => "0110101101110000",
39539 => "0110101101110000",
39540 => "0110101101110000",
39541 => "0110101101110000",
39542 => "0110101101110000",
39543 => "0110101101110000",
39544 => "0110101101110000",
39545 => "0110101101110000",
39546 => "0110101101110000",
39547 => "0110101101110000",
39548 => "0110101110000000",
39549 => "0110101110000000",
39550 => "0110101110000000",
39551 => "0110101110000000",
39552 => "0110101110000000",
39553 => "0110101110000000",
39554 => "0110101110000000",
39555 => "0110101110000000",
39556 => "0110101110000000",
39557 => "0110101110000000",
39558 => "0110101110000000",
39559 => "0110101110000000",
39560 => "0110101110000000",
39561 => "0110101110000000",
39562 => "0110101110000000",
39563 => "0110101110010000",
39564 => "0110101110010000",
39565 => "0110101110010000",
39566 => "0110101110010000",
39567 => "0110101110010000",
39568 => "0110101110010000",
39569 => "0110101110010000",
39570 => "0110101110010000",
39571 => "0110101110010000",
39572 => "0110101110010000",
39573 => "0110101110010000",
39574 => "0110101110010000",
39575 => "0110101110010000",
39576 => "0110101110010000",
39577 => "0110101110010000",
39578 => "0110101110100000",
39579 => "0110101110100000",
39580 => "0110101110100000",
39581 => "0110101110100000",
39582 => "0110101110100000",
39583 => "0110101110100000",
39584 => "0110101110100000",
39585 => "0110101110100000",
39586 => "0110101110100000",
39587 => "0110101110100000",
39588 => "0110101110100000",
39589 => "0110101110100000",
39590 => "0110101110100000",
39591 => "0110101110100000",
39592 => "0110101110100000",
39593 => "0110101110110000",
39594 => "0110101110110000",
39595 => "0110101110110000",
39596 => "0110101110110000",
39597 => "0110101110110000",
39598 => "0110101110110000",
39599 => "0110101110110000",
39600 => "0110101110110000",
39601 => "0110101110110000",
39602 => "0110101110110000",
39603 => "0110101110110000",
39604 => "0110101110110000",
39605 => "0110101110110000",
39606 => "0110101110110000",
39607 => "0110101110110000",
39608 => "0110101111000000",
39609 => "0110101111000000",
39610 => "0110101111000000",
39611 => "0110101111000000",
39612 => "0110101111000000",
39613 => "0110101111000000",
39614 => "0110101111000000",
39615 => "0110101111000000",
39616 => "0110101111000000",
39617 => "0110101111000000",
39618 => "0110101111000000",
39619 => "0110101111000000",
39620 => "0110101111000000",
39621 => "0110101111000000",
39622 => "0110101111000000",
39623 => "0110101111010000",
39624 => "0110101111010000",
39625 => "0110101111010000",
39626 => "0110101111010000",
39627 => "0110101111010000",
39628 => "0110101111010000",
39629 => "0110101111010000",
39630 => "0110101111010000",
39631 => "0110101111010000",
39632 => "0110101111010000",
39633 => "0110101111010000",
39634 => "0110101111010000",
39635 => "0110101111010000",
39636 => "0110101111010000",
39637 => "0110101111010000",
39638 => "0110101111100000",
39639 => "0110101111100000",
39640 => "0110101111100000",
39641 => "0110101111100000",
39642 => "0110101111100000",
39643 => "0110101111100000",
39644 => "0110101111100000",
39645 => "0110101111100000",
39646 => "0110101111100000",
39647 => "0110101111100000",
39648 => "0110101111100000",
39649 => "0110101111100000",
39650 => "0110101111100000",
39651 => "0110101111100000",
39652 => "0110101111100000",
39653 => "0110101111110000",
39654 => "0110101111110000",
39655 => "0110101111110000",
39656 => "0110101111110000",
39657 => "0110101111110000",
39658 => "0110101111110000",
39659 => "0110101111110000",
39660 => "0110101111110000",
39661 => "0110101111110000",
39662 => "0110101111110000",
39663 => "0110101111110000",
39664 => "0110101111110000",
39665 => "0110101111110000",
39666 => "0110101111110000",
39667 => "0110101111110000",
39668 => "0110110000000000",
39669 => "0110110000000000",
39670 => "0110110000000000",
39671 => "0110110000000000",
39672 => "0110110000000000",
39673 => "0110110000000000",
39674 => "0110110000000000",
39675 => "0110110000000000",
39676 => "0110110000000000",
39677 => "0110110000000000",
39678 => "0110110000000000",
39679 => "0110110000000000",
39680 => "0110110000000000",
39681 => "0110110000000000",
39682 => "0110110000000000",
39683 => "0110110000010000",
39684 => "0110110000010000",
39685 => "0110110000010000",
39686 => "0110110000010000",
39687 => "0110110000010000",
39688 => "0110110000010000",
39689 => "0110110000010000",
39690 => "0110110000010000",
39691 => "0110110000010000",
39692 => "0110110000010000",
39693 => "0110110000010000",
39694 => "0110110000010000",
39695 => "0110110000010000",
39696 => "0110110000010000",
39697 => "0110110000010000",
39698 => "0110110000100000",
39699 => "0110110000100000",
39700 => "0110110000100000",
39701 => "0110110000100000",
39702 => "0110110000100000",
39703 => "0110110000100000",
39704 => "0110110000100000",
39705 => "0110110000100000",
39706 => "0110110000100000",
39707 => "0110110000100000",
39708 => "0110110000100000",
39709 => "0110110000100000",
39710 => "0110110000100000",
39711 => "0110110000100000",
39712 => "0110110000100000",
39713 => "0110110000110000",
39714 => "0110110000110000",
39715 => "0110110000110000",
39716 => "0110110000110000",
39717 => "0110110000110000",
39718 => "0110110000110000",
39719 => "0110110000110000",
39720 => "0110110000110000",
39721 => "0110110000110000",
39722 => "0110110000110000",
39723 => "0110110000110000",
39724 => "0110110000110000",
39725 => "0110110000110000",
39726 => "0110110000110000",
39727 => "0110110000110000",
39728 => "0110110000110000",
39729 => "0110110001000000",
39730 => "0110110001000000",
39731 => "0110110001000000",
39732 => "0110110001000000",
39733 => "0110110001000000",
39734 => "0110110001000000",
39735 => "0110110001000000",
39736 => "0110110001000000",
39737 => "0110110001000000",
39738 => "0110110001000000",
39739 => "0110110001000000",
39740 => "0110110001000000",
39741 => "0110110001000000",
39742 => "0110110001000000",
39743 => "0110110001000000",
39744 => "0110110001010000",
39745 => "0110110001010000",
39746 => "0110110001010000",
39747 => "0110110001010000",
39748 => "0110110001010000",
39749 => "0110110001010000",
39750 => "0110110001010000",
39751 => "0110110001010000",
39752 => "0110110001010000",
39753 => "0110110001010000",
39754 => "0110110001010000",
39755 => "0110110001010000",
39756 => "0110110001010000",
39757 => "0110110001010000",
39758 => "0110110001010000",
39759 => "0110110001100000",
39760 => "0110110001100000",
39761 => "0110110001100000",
39762 => "0110110001100000",
39763 => "0110110001100000",
39764 => "0110110001100000",
39765 => "0110110001100000",
39766 => "0110110001100000",
39767 => "0110110001100000",
39768 => "0110110001100000",
39769 => "0110110001100000",
39770 => "0110110001100000",
39771 => "0110110001100000",
39772 => "0110110001100000",
39773 => "0110110001100000",
39774 => "0110110001100000",
39775 => "0110110001110000",
39776 => "0110110001110000",
39777 => "0110110001110000",
39778 => "0110110001110000",
39779 => "0110110001110000",
39780 => "0110110001110000",
39781 => "0110110001110000",
39782 => "0110110001110000",
39783 => "0110110001110000",
39784 => "0110110001110000",
39785 => "0110110001110000",
39786 => "0110110001110000",
39787 => "0110110001110000",
39788 => "0110110001110000",
39789 => "0110110001110000",
39790 => "0110110010000000",
39791 => "0110110010000000",
39792 => "0110110010000000",
39793 => "0110110010000000",
39794 => "0110110010000000",
39795 => "0110110010000000",
39796 => "0110110010000000",
39797 => "0110110010000000",
39798 => "0110110010000000",
39799 => "0110110010000000",
39800 => "0110110010000000",
39801 => "0110110010000000",
39802 => "0110110010000000",
39803 => "0110110010000000",
39804 => "0110110010000000",
39805 => "0110110010000000",
39806 => "0110110010010000",
39807 => "0110110010010000",
39808 => "0110110010010000",
39809 => "0110110010010000",
39810 => "0110110010010000",
39811 => "0110110010010000",
39812 => "0110110010010000",
39813 => "0110110010010000",
39814 => "0110110010010000",
39815 => "0110110010010000",
39816 => "0110110010010000",
39817 => "0110110010010000",
39818 => "0110110010010000",
39819 => "0110110010010000",
39820 => "0110110010010000",
39821 => "0110110010100000",
39822 => "0110110010100000",
39823 => "0110110010100000",
39824 => "0110110010100000",
39825 => "0110110010100000",
39826 => "0110110010100000",
39827 => "0110110010100000",
39828 => "0110110010100000",
39829 => "0110110010100000",
39830 => "0110110010100000",
39831 => "0110110010100000",
39832 => "0110110010100000",
39833 => "0110110010100000",
39834 => "0110110010100000",
39835 => "0110110010100000",
39836 => "0110110010100000",
39837 => "0110110010110000",
39838 => "0110110010110000",
39839 => "0110110010110000",
39840 => "0110110010110000",
39841 => "0110110010110000",
39842 => "0110110010110000",
39843 => "0110110010110000",
39844 => "0110110010110000",
39845 => "0110110010110000",
39846 => "0110110010110000",
39847 => "0110110010110000",
39848 => "0110110010110000",
39849 => "0110110010110000",
39850 => "0110110010110000",
39851 => "0110110010110000",
39852 => "0110110011000000",
39853 => "0110110011000000",
39854 => "0110110011000000",
39855 => "0110110011000000",
39856 => "0110110011000000",
39857 => "0110110011000000",
39858 => "0110110011000000",
39859 => "0110110011000000",
39860 => "0110110011000000",
39861 => "0110110011000000",
39862 => "0110110011000000",
39863 => "0110110011000000",
39864 => "0110110011000000",
39865 => "0110110011000000",
39866 => "0110110011000000",
39867 => "0110110011000000",
39868 => "0110110011010000",
39869 => "0110110011010000",
39870 => "0110110011010000",
39871 => "0110110011010000",
39872 => "0110110011010000",
39873 => "0110110011010000",
39874 => "0110110011010000",
39875 => "0110110011010000",
39876 => "0110110011010000",
39877 => "0110110011010000",
39878 => "0110110011010000",
39879 => "0110110011010000",
39880 => "0110110011010000",
39881 => "0110110011010000",
39882 => "0110110011010000",
39883 => "0110110011010000",
39884 => "0110110011100000",
39885 => "0110110011100000",
39886 => "0110110011100000",
39887 => "0110110011100000",
39888 => "0110110011100000",
39889 => "0110110011100000",
39890 => "0110110011100000",
39891 => "0110110011100000",
39892 => "0110110011100000",
39893 => "0110110011100000",
39894 => "0110110011100000",
39895 => "0110110011100000",
39896 => "0110110011100000",
39897 => "0110110011100000",
39898 => "0110110011100000",
39899 => "0110110011100000",
39900 => "0110110011110000",
39901 => "0110110011110000",
39902 => "0110110011110000",
39903 => "0110110011110000",
39904 => "0110110011110000",
39905 => "0110110011110000",
39906 => "0110110011110000",
39907 => "0110110011110000",
39908 => "0110110011110000",
39909 => "0110110011110000",
39910 => "0110110011110000",
39911 => "0110110011110000",
39912 => "0110110011110000",
39913 => "0110110011110000",
39914 => "0110110011110000",
39915 => "0110110100000000",
39916 => "0110110100000000",
39917 => "0110110100000000",
39918 => "0110110100000000",
39919 => "0110110100000000",
39920 => "0110110100000000",
39921 => "0110110100000000",
39922 => "0110110100000000",
39923 => "0110110100000000",
39924 => "0110110100000000",
39925 => "0110110100000000",
39926 => "0110110100000000",
39927 => "0110110100000000",
39928 => "0110110100000000",
39929 => "0110110100000000",
39930 => "0110110100000000",
39931 => "0110110100010000",
39932 => "0110110100010000",
39933 => "0110110100010000",
39934 => "0110110100010000",
39935 => "0110110100010000",
39936 => "0110110100010000",
39937 => "0110110100010000",
39938 => "0110110100010000",
39939 => "0110110100010000",
39940 => "0110110100010000",
39941 => "0110110100010000",
39942 => "0110110100010000",
39943 => "0110110100010000",
39944 => "0110110100010000",
39945 => "0110110100010000",
39946 => "0110110100010000",
39947 => "0110110100100000",
39948 => "0110110100100000",
39949 => "0110110100100000",
39950 => "0110110100100000",
39951 => "0110110100100000",
39952 => "0110110100100000",
39953 => "0110110100100000",
39954 => "0110110100100000",
39955 => "0110110100100000",
39956 => "0110110100100000",
39957 => "0110110100100000",
39958 => "0110110100100000",
39959 => "0110110100100000",
39960 => "0110110100100000",
39961 => "0110110100100000",
39962 => "0110110100100000",
39963 => "0110110100110000",
39964 => "0110110100110000",
39965 => "0110110100110000",
39966 => "0110110100110000",
39967 => "0110110100110000",
39968 => "0110110100110000",
39969 => "0110110100110000",
39970 => "0110110100110000",
39971 => "0110110100110000",
39972 => "0110110100110000",
39973 => "0110110100110000",
39974 => "0110110100110000",
39975 => "0110110100110000",
39976 => "0110110100110000",
39977 => "0110110100110000",
39978 => "0110110100110000",
39979 => "0110110101000000",
39980 => "0110110101000000",
39981 => "0110110101000000",
39982 => "0110110101000000",
39983 => "0110110101000000",
39984 => "0110110101000000",
39985 => "0110110101000000",
39986 => "0110110101000000",
39987 => "0110110101000000",
39988 => "0110110101000000",
39989 => "0110110101000000",
39990 => "0110110101000000",
39991 => "0110110101000000",
39992 => "0110110101000000",
39993 => "0110110101000000",
39994 => "0110110101000000",
39995 => "0110110101010000",
39996 => "0110110101010000",
39997 => "0110110101010000",
39998 => "0110110101010000",
39999 => "0110110101010000",
40000 => "0110110101010000",
40001 => "0110110101010000",
40002 => "0110110101010000",
40003 => "0110110101010000",
40004 => "0110110101010000",
40005 => "0110110101010000",
40006 => "0110110101010000",
40007 => "0110110101010000",
40008 => "0110110101010000",
40009 => "0110110101010000",
40010 => "0110110101010000",
40011 => "0110110101100000",
40012 => "0110110101100000",
40013 => "0110110101100000",
40014 => "0110110101100000",
40015 => "0110110101100000",
40016 => "0110110101100000",
40017 => "0110110101100000",
40018 => "0110110101100000",
40019 => "0110110101100000",
40020 => "0110110101100000",
40021 => "0110110101100000",
40022 => "0110110101100000",
40023 => "0110110101100000",
40024 => "0110110101100000",
40025 => "0110110101100000",
40026 => "0110110101100000",
40027 => "0110110101110000",
40028 => "0110110101110000",
40029 => "0110110101110000",
40030 => "0110110101110000",
40031 => "0110110101110000",
40032 => "0110110101110000",
40033 => "0110110101110000",
40034 => "0110110101110000",
40035 => "0110110101110000",
40036 => "0110110101110000",
40037 => "0110110101110000",
40038 => "0110110101110000",
40039 => "0110110101110000",
40040 => "0110110101110000",
40041 => "0110110101110000",
40042 => "0110110101110000",
40043 => "0110110110000000",
40044 => "0110110110000000",
40045 => "0110110110000000",
40046 => "0110110110000000",
40047 => "0110110110000000",
40048 => "0110110110000000",
40049 => "0110110110000000",
40050 => "0110110110000000",
40051 => "0110110110000000",
40052 => "0110110110000000",
40053 => "0110110110000000",
40054 => "0110110110000000",
40055 => "0110110110000000",
40056 => "0110110110000000",
40057 => "0110110110000000",
40058 => "0110110110000000",
40059 => "0110110110010000",
40060 => "0110110110010000",
40061 => "0110110110010000",
40062 => "0110110110010000",
40063 => "0110110110010000",
40064 => "0110110110010000",
40065 => "0110110110010000",
40066 => "0110110110010000",
40067 => "0110110110010000",
40068 => "0110110110010000",
40069 => "0110110110010000",
40070 => "0110110110010000",
40071 => "0110110110010000",
40072 => "0110110110010000",
40073 => "0110110110010000",
40074 => "0110110110010000",
40075 => "0110110110010000",
40076 => "0110110110100000",
40077 => "0110110110100000",
40078 => "0110110110100000",
40079 => "0110110110100000",
40080 => "0110110110100000",
40081 => "0110110110100000",
40082 => "0110110110100000",
40083 => "0110110110100000",
40084 => "0110110110100000",
40085 => "0110110110100000",
40086 => "0110110110100000",
40087 => "0110110110100000",
40088 => "0110110110100000",
40089 => "0110110110100000",
40090 => "0110110110100000",
40091 => "0110110110100000",
40092 => "0110110110110000",
40093 => "0110110110110000",
40094 => "0110110110110000",
40095 => "0110110110110000",
40096 => "0110110110110000",
40097 => "0110110110110000",
40098 => "0110110110110000",
40099 => "0110110110110000",
40100 => "0110110110110000",
40101 => "0110110110110000",
40102 => "0110110110110000",
40103 => "0110110110110000",
40104 => "0110110110110000",
40105 => "0110110110110000",
40106 => "0110110110110000",
40107 => "0110110110110000",
40108 => "0110110111000000",
40109 => "0110110111000000",
40110 => "0110110111000000",
40111 => "0110110111000000",
40112 => "0110110111000000",
40113 => "0110110111000000",
40114 => "0110110111000000",
40115 => "0110110111000000",
40116 => "0110110111000000",
40117 => "0110110111000000",
40118 => "0110110111000000",
40119 => "0110110111000000",
40120 => "0110110111000000",
40121 => "0110110111000000",
40122 => "0110110111000000",
40123 => "0110110111000000",
40124 => "0110110111010000",
40125 => "0110110111010000",
40126 => "0110110111010000",
40127 => "0110110111010000",
40128 => "0110110111010000",
40129 => "0110110111010000",
40130 => "0110110111010000",
40131 => "0110110111010000",
40132 => "0110110111010000",
40133 => "0110110111010000",
40134 => "0110110111010000",
40135 => "0110110111010000",
40136 => "0110110111010000",
40137 => "0110110111010000",
40138 => "0110110111010000",
40139 => "0110110111010000",
40140 => "0110110111010000",
40141 => "0110110111100000",
40142 => "0110110111100000",
40143 => "0110110111100000",
40144 => "0110110111100000",
40145 => "0110110111100000",
40146 => "0110110111100000",
40147 => "0110110111100000",
40148 => "0110110111100000",
40149 => "0110110111100000",
40150 => "0110110111100000",
40151 => "0110110111100000",
40152 => "0110110111100000",
40153 => "0110110111100000",
40154 => "0110110111100000",
40155 => "0110110111100000",
40156 => "0110110111100000",
40157 => "0110110111110000",
40158 => "0110110111110000",
40159 => "0110110111110000",
40160 => "0110110111110000",
40161 => "0110110111110000",
40162 => "0110110111110000",
40163 => "0110110111110000",
40164 => "0110110111110000",
40165 => "0110110111110000",
40166 => "0110110111110000",
40167 => "0110110111110000",
40168 => "0110110111110000",
40169 => "0110110111110000",
40170 => "0110110111110000",
40171 => "0110110111110000",
40172 => "0110110111110000",
40173 => "0110110111110000",
40174 => "0110111000000000",
40175 => "0110111000000000",
40176 => "0110111000000000",
40177 => "0110111000000000",
40178 => "0110111000000000",
40179 => "0110111000000000",
40180 => "0110111000000000",
40181 => "0110111000000000",
40182 => "0110111000000000",
40183 => "0110111000000000",
40184 => "0110111000000000",
40185 => "0110111000000000",
40186 => "0110111000000000",
40187 => "0110111000000000",
40188 => "0110111000000000",
40189 => "0110111000000000",
40190 => "0110111000010000",
40191 => "0110111000010000",
40192 => "0110111000010000",
40193 => "0110111000010000",
40194 => "0110111000010000",
40195 => "0110111000010000",
40196 => "0110111000010000",
40197 => "0110111000010000",
40198 => "0110111000010000",
40199 => "0110111000010000",
40200 => "0110111000010000",
40201 => "0110111000010000",
40202 => "0110111000010000",
40203 => "0110111000010000",
40204 => "0110111000010000",
40205 => "0110111000010000",
40206 => "0110111000010000",
40207 => "0110111000100000",
40208 => "0110111000100000",
40209 => "0110111000100000",
40210 => "0110111000100000",
40211 => "0110111000100000",
40212 => "0110111000100000",
40213 => "0110111000100000",
40214 => "0110111000100000",
40215 => "0110111000100000",
40216 => "0110111000100000",
40217 => "0110111000100000",
40218 => "0110111000100000",
40219 => "0110111000100000",
40220 => "0110111000100000",
40221 => "0110111000100000",
40222 => "0110111000100000",
40223 => "0110111000100000",
40224 => "0110111000110000",
40225 => "0110111000110000",
40226 => "0110111000110000",
40227 => "0110111000110000",
40228 => "0110111000110000",
40229 => "0110111000110000",
40230 => "0110111000110000",
40231 => "0110111000110000",
40232 => "0110111000110000",
40233 => "0110111000110000",
40234 => "0110111000110000",
40235 => "0110111000110000",
40236 => "0110111000110000",
40237 => "0110111000110000",
40238 => "0110111000110000",
40239 => "0110111000110000",
40240 => "0110111001000000",
40241 => "0110111001000000",
40242 => "0110111001000000",
40243 => "0110111001000000",
40244 => "0110111001000000",
40245 => "0110111001000000",
40246 => "0110111001000000",
40247 => "0110111001000000",
40248 => "0110111001000000",
40249 => "0110111001000000",
40250 => "0110111001000000",
40251 => "0110111001000000",
40252 => "0110111001000000",
40253 => "0110111001000000",
40254 => "0110111001000000",
40255 => "0110111001000000",
40256 => "0110111001000000",
40257 => "0110111001010000",
40258 => "0110111001010000",
40259 => "0110111001010000",
40260 => "0110111001010000",
40261 => "0110111001010000",
40262 => "0110111001010000",
40263 => "0110111001010000",
40264 => "0110111001010000",
40265 => "0110111001010000",
40266 => "0110111001010000",
40267 => "0110111001010000",
40268 => "0110111001010000",
40269 => "0110111001010000",
40270 => "0110111001010000",
40271 => "0110111001010000",
40272 => "0110111001010000",
40273 => "0110111001010000",
40274 => "0110111001100000",
40275 => "0110111001100000",
40276 => "0110111001100000",
40277 => "0110111001100000",
40278 => "0110111001100000",
40279 => "0110111001100000",
40280 => "0110111001100000",
40281 => "0110111001100000",
40282 => "0110111001100000",
40283 => "0110111001100000",
40284 => "0110111001100000",
40285 => "0110111001100000",
40286 => "0110111001100000",
40287 => "0110111001100000",
40288 => "0110111001100000",
40289 => "0110111001100000",
40290 => "0110111001100000",
40291 => "0110111001110000",
40292 => "0110111001110000",
40293 => "0110111001110000",
40294 => "0110111001110000",
40295 => "0110111001110000",
40296 => "0110111001110000",
40297 => "0110111001110000",
40298 => "0110111001110000",
40299 => "0110111001110000",
40300 => "0110111001110000",
40301 => "0110111001110000",
40302 => "0110111001110000",
40303 => "0110111001110000",
40304 => "0110111001110000",
40305 => "0110111001110000",
40306 => "0110111001110000",
40307 => "0110111001110000",
40308 => "0110111010000000",
40309 => "0110111010000000",
40310 => "0110111010000000",
40311 => "0110111010000000",
40312 => "0110111010000000",
40313 => "0110111010000000",
40314 => "0110111010000000",
40315 => "0110111010000000",
40316 => "0110111010000000",
40317 => "0110111010000000",
40318 => "0110111010000000",
40319 => "0110111010000000",
40320 => "0110111010000000",
40321 => "0110111010000000",
40322 => "0110111010000000",
40323 => "0110111010000000",
40324 => "0110111010000000",
40325 => "0110111010010000",
40326 => "0110111010010000",
40327 => "0110111010010000",
40328 => "0110111010010000",
40329 => "0110111010010000",
40330 => "0110111010010000",
40331 => "0110111010010000",
40332 => "0110111010010000",
40333 => "0110111010010000",
40334 => "0110111010010000",
40335 => "0110111010010000",
40336 => "0110111010010000",
40337 => "0110111010010000",
40338 => "0110111010010000",
40339 => "0110111010010000",
40340 => "0110111010010000",
40341 => "0110111010010000",
40342 => "0110111010100000",
40343 => "0110111010100000",
40344 => "0110111010100000",
40345 => "0110111010100000",
40346 => "0110111010100000",
40347 => "0110111010100000",
40348 => "0110111010100000",
40349 => "0110111010100000",
40350 => "0110111010100000",
40351 => "0110111010100000",
40352 => "0110111010100000",
40353 => "0110111010100000",
40354 => "0110111010100000",
40355 => "0110111010100000",
40356 => "0110111010100000",
40357 => "0110111010100000",
40358 => "0110111010100000",
40359 => "0110111010110000",
40360 => "0110111010110000",
40361 => "0110111010110000",
40362 => "0110111010110000",
40363 => "0110111010110000",
40364 => "0110111010110000",
40365 => "0110111010110000",
40366 => "0110111010110000",
40367 => "0110111010110000",
40368 => "0110111010110000",
40369 => "0110111010110000",
40370 => "0110111010110000",
40371 => "0110111010110000",
40372 => "0110111010110000",
40373 => "0110111010110000",
40374 => "0110111010110000",
40375 => "0110111010110000",
40376 => "0110111011000000",
40377 => "0110111011000000",
40378 => "0110111011000000",
40379 => "0110111011000000",
40380 => "0110111011000000",
40381 => "0110111011000000",
40382 => "0110111011000000",
40383 => "0110111011000000",
40384 => "0110111011000000",
40385 => "0110111011000000",
40386 => "0110111011000000",
40387 => "0110111011000000",
40388 => "0110111011000000",
40389 => "0110111011000000",
40390 => "0110111011000000",
40391 => "0110111011000000",
40392 => "0110111011000000",
40393 => "0110111011010000",
40394 => "0110111011010000",
40395 => "0110111011010000",
40396 => "0110111011010000",
40397 => "0110111011010000",
40398 => "0110111011010000",
40399 => "0110111011010000",
40400 => "0110111011010000",
40401 => "0110111011010000",
40402 => "0110111011010000",
40403 => "0110111011010000",
40404 => "0110111011010000",
40405 => "0110111011010000",
40406 => "0110111011010000",
40407 => "0110111011010000",
40408 => "0110111011010000",
40409 => "0110111011010000",
40410 => "0110111011100000",
40411 => "0110111011100000",
40412 => "0110111011100000",
40413 => "0110111011100000",
40414 => "0110111011100000",
40415 => "0110111011100000",
40416 => "0110111011100000",
40417 => "0110111011100000",
40418 => "0110111011100000",
40419 => "0110111011100000",
40420 => "0110111011100000",
40421 => "0110111011100000",
40422 => "0110111011100000",
40423 => "0110111011100000",
40424 => "0110111011100000",
40425 => "0110111011100000",
40426 => "0110111011100000",
40427 => "0110111011110000",
40428 => "0110111011110000",
40429 => "0110111011110000",
40430 => "0110111011110000",
40431 => "0110111011110000",
40432 => "0110111011110000",
40433 => "0110111011110000",
40434 => "0110111011110000",
40435 => "0110111011110000",
40436 => "0110111011110000",
40437 => "0110111011110000",
40438 => "0110111011110000",
40439 => "0110111011110000",
40440 => "0110111011110000",
40441 => "0110111011110000",
40442 => "0110111011110000",
40443 => "0110111011110000",
40444 => "0110111011110000",
40445 => "0110111100000000",
40446 => "0110111100000000",
40447 => "0110111100000000",
40448 => "0110111100000000",
40449 => "0110111100000000",
40450 => "0110111100000000",
40451 => "0110111100000000",
40452 => "0110111100000000",
40453 => "0110111100000000",
40454 => "0110111100000000",
40455 => "0110111100000000",
40456 => "0110111100000000",
40457 => "0110111100000000",
40458 => "0110111100000000",
40459 => "0110111100000000",
40460 => "0110111100000000",
40461 => "0110111100000000",
40462 => "0110111100010000",
40463 => "0110111100010000",
40464 => "0110111100010000",
40465 => "0110111100010000",
40466 => "0110111100010000",
40467 => "0110111100010000",
40468 => "0110111100010000",
40469 => "0110111100010000",
40470 => "0110111100010000",
40471 => "0110111100010000",
40472 => "0110111100010000",
40473 => "0110111100010000",
40474 => "0110111100010000",
40475 => "0110111100010000",
40476 => "0110111100010000",
40477 => "0110111100010000",
40478 => "0110111100010000",
40479 => "0110111100100000",
40480 => "0110111100100000",
40481 => "0110111100100000",
40482 => "0110111100100000",
40483 => "0110111100100000",
40484 => "0110111100100000",
40485 => "0110111100100000",
40486 => "0110111100100000",
40487 => "0110111100100000",
40488 => "0110111100100000",
40489 => "0110111100100000",
40490 => "0110111100100000",
40491 => "0110111100100000",
40492 => "0110111100100000",
40493 => "0110111100100000",
40494 => "0110111100100000",
40495 => "0110111100100000",
40496 => "0110111100100000",
40497 => "0110111100110000",
40498 => "0110111100110000",
40499 => "0110111100110000",
40500 => "0110111100110000",
40501 => "0110111100110000",
40502 => "0110111100110000",
40503 => "0110111100110000",
40504 => "0110111100110000",
40505 => "0110111100110000",
40506 => "0110111100110000",
40507 => "0110111100110000",
40508 => "0110111100110000",
40509 => "0110111100110000",
40510 => "0110111100110000",
40511 => "0110111100110000",
40512 => "0110111100110000",
40513 => "0110111100110000",
40514 => "0110111101000000",
40515 => "0110111101000000",
40516 => "0110111101000000",
40517 => "0110111101000000",
40518 => "0110111101000000",
40519 => "0110111101000000",
40520 => "0110111101000000",
40521 => "0110111101000000",
40522 => "0110111101000000",
40523 => "0110111101000000",
40524 => "0110111101000000",
40525 => "0110111101000000",
40526 => "0110111101000000",
40527 => "0110111101000000",
40528 => "0110111101000000",
40529 => "0110111101000000",
40530 => "0110111101000000",
40531 => "0110111101000000",
40532 => "0110111101010000",
40533 => "0110111101010000",
40534 => "0110111101010000",
40535 => "0110111101010000",
40536 => "0110111101010000",
40537 => "0110111101010000",
40538 => "0110111101010000",
40539 => "0110111101010000",
40540 => "0110111101010000",
40541 => "0110111101010000",
40542 => "0110111101010000",
40543 => "0110111101010000",
40544 => "0110111101010000",
40545 => "0110111101010000",
40546 => "0110111101010000",
40547 => "0110111101010000",
40548 => "0110111101010000",
40549 => "0110111101010000",
40550 => "0110111101100000",
40551 => "0110111101100000",
40552 => "0110111101100000",
40553 => "0110111101100000",
40554 => "0110111101100000",
40555 => "0110111101100000",
40556 => "0110111101100000",
40557 => "0110111101100000",
40558 => "0110111101100000",
40559 => "0110111101100000",
40560 => "0110111101100000",
40561 => "0110111101100000",
40562 => "0110111101100000",
40563 => "0110111101100000",
40564 => "0110111101100000",
40565 => "0110111101100000",
40566 => "0110111101100000",
40567 => "0110111101110000",
40568 => "0110111101110000",
40569 => "0110111101110000",
40570 => "0110111101110000",
40571 => "0110111101110000",
40572 => "0110111101110000",
40573 => "0110111101110000",
40574 => "0110111101110000",
40575 => "0110111101110000",
40576 => "0110111101110000",
40577 => "0110111101110000",
40578 => "0110111101110000",
40579 => "0110111101110000",
40580 => "0110111101110000",
40581 => "0110111101110000",
40582 => "0110111101110000",
40583 => "0110111101110000",
40584 => "0110111101110000",
40585 => "0110111110000000",
40586 => "0110111110000000",
40587 => "0110111110000000",
40588 => "0110111110000000",
40589 => "0110111110000000",
40590 => "0110111110000000",
40591 => "0110111110000000",
40592 => "0110111110000000",
40593 => "0110111110000000",
40594 => "0110111110000000",
40595 => "0110111110000000",
40596 => "0110111110000000",
40597 => "0110111110000000",
40598 => "0110111110000000",
40599 => "0110111110000000",
40600 => "0110111110000000",
40601 => "0110111110000000",
40602 => "0110111110000000",
40603 => "0110111110010000",
40604 => "0110111110010000",
40605 => "0110111110010000",
40606 => "0110111110010000",
40607 => "0110111110010000",
40608 => "0110111110010000",
40609 => "0110111110010000",
40610 => "0110111110010000",
40611 => "0110111110010000",
40612 => "0110111110010000",
40613 => "0110111110010000",
40614 => "0110111110010000",
40615 => "0110111110010000",
40616 => "0110111110010000",
40617 => "0110111110010000",
40618 => "0110111110010000",
40619 => "0110111110010000",
40620 => "0110111110010000",
40621 => "0110111110100000",
40622 => "0110111110100000",
40623 => "0110111110100000",
40624 => "0110111110100000",
40625 => "0110111110100000",
40626 => "0110111110100000",
40627 => "0110111110100000",
40628 => "0110111110100000",
40629 => "0110111110100000",
40630 => "0110111110100000",
40631 => "0110111110100000",
40632 => "0110111110100000",
40633 => "0110111110100000",
40634 => "0110111110100000",
40635 => "0110111110100000",
40636 => "0110111110100000",
40637 => "0110111110100000",
40638 => "0110111110100000",
40639 => "0110111110110000",
40640 => "0110111110110000",
40641 => "0110111110110000",
40642 => "0110111110110000",
40643 => "0110111110110000",
40644 => "0110111110110000",
40645 => "0110111110110000",
40646 => "0110111110110000",
40647 => "0110111110110000",
40648 => "0110111110110000",
40649 => "0110111110110000",
40650 => "0110111110110000",
40651 => "0110111110110000",
40652 => "0110111110110000",
40653 => "0110111110110000",
40654 => "0110111110110000",
40655 => "0110111110110000",
40656 => "0110111110110000",
40657 => "0110111111000000",
40658 => "0110111111000000",
40659 => "0110111111000000",
40660 => "0110111111000000",
40661 => "0110111111000000",
40662 => "0110111111000000",
40663 => "0110111111000000",
40664 => "0110111111000000",
40665 => "0110111111000000",
40666 => "0110111111000000",
40667 => "0110111111000000",
40668 => "0110111111000000",
40669 => "0110111111000000",
40670 => "0110111111000000",
40671 => "0110111111000000",
40672 => "0110111111000000",
40673 => "0110111111000000",
40674 => "0110111111000000",
40675 => "0110111111010000",
40676 => "0110111111010000",
40677 => "0110111111010000",
40678 => "0110111111010000",
40679 => "0110111111010000",
40680 => "0110111111010000",
40681 => "0110111111010000",
40682 => "0110111111010000",
40683 => "0110111111010000",
40684 => "0110111111010000",
40685 => "0110111111010000",
40686 => "0110111111010000",
40687 => "0110111111010000",
40688 => "0110111111010000",
40689 => "0110111111010000",
40690 => "0110111111010000",
40691 => "0110111111010000",
40692 => "0110111111010000",
40693 => "0110111111100000",
40694 => "0110111111100000",
40695 => "0110111111100000",
40696 => "0110111111100000",
40697 => "0110111111100000",
40698 => "0110111111100000",
40699 => "0110111111100000",
40700 => "0110111111100000",
40701 => "0110111111100000",
40702 => "0110111111100000",
40703 => "0110111111100000",
40704 => "0110111111100000",
40705 => "0110111111100000",
40706 => "0110111111100000",
40707 => "0110111111100000",
40708 => "0110111111100000",
40709 => "0110111111100000",
40710 => "0110111111100000",
40711 => "0110111111110000",
40712 => "0110111111110000",
40713 => "0110111111110000",
40714 => "0110111111110000",
40715 => "0110111111110000",
40716 => "0110111111110000",
40717 => "0110111111110000",
40718 => "0110111111110000",
40719 => "0110111111110000",
40720 => "0110111111110000",
40721 => "0110111111110000",
40722 => "0110111111110000",
40723 => "0110111111110000",
40724 => "0110111111110000",
40725 => "0110111111110000",
40726 => "0110111111110000",
40727 => "0110111111110000",
40728 => "0110111111110000",
40729 => "0111000000000000",
40730 => "0111000000000000",
40731 => "0111000000000000",
40732 => "0111000000000000",
40733 => "0111000000000000",
40734 => "0111000000000000",
40735 => "0111000000000000",
40736 => "0111000000000000",
40737 => "0111000000000000",
40738 => "0111000000000000",
40739 => "0111000000000000",
40740 => "0111000000000000",
40741 => "0111000000000000",
40742 => "0111000000000000",
40743 => "0111000000000000",
40744 => "0111000000000000",
40745 => "0111000000000000",
40746 => "0111000000000000",
40747 => "0111000000010000",
40748 => "0111000000010000",
40749 => "0111000000010000",
40750 => "0111000000010000",
40751 => "0111000000010000",
40752 => "0111000000010000",
40753 => "0111000000010000",
40754 => "0111000000010000",
40755 => "0111000000010000",
40756 => "0111000000010000",
40757 => "0111000000010000",
40758 => "0111000000010000",
40759 => "0111000000010000",
40760 => "0111000000010000",
40761 => "0111000000010000",
40762 => "0111000000010000",
40763 => "0111000000010000",
40764 => "0111000000010000",
40765 => "0111000000010000",
40766 => "0111000000100000",
40767 => "0111000000100000",
40768 => "0111000000100000",
40769 => "0111000000100000",
40770 => "0111000000100000",
40771 => "0111000000100000",
40772 => "0111000000100000",
40773 => "0111000000100000",
40774 => "0111000000100000",
40775 => "0111000000100000",
40776 => "0111000000100000",
40777 => "0111000000100000",
40778 => "0111000000100000",
40779 => "0111000000100000",
40780 => "0111000000100000",
40781 => "0111000000100000",
40782 => "0111000000100000",
40783 => "0111000000100000",
40784 => "0111000000110000",
40785 => "0111000000110000",
40786 => "0111000000110000",
40787 => "0111000000110000",
40788 => "0111000000110000",
40789 => "0111000000110000",
40790 => "0111000000110000",
40791 => "0111000000110000",
40792 => "0111000000110000",
40793 => "0111000000110000",
40794 => "0111000000110000",
40795 => "0111000000110000",
40796 => "0111000000110000",
40797 => "0111000000110000",
40798 => "0111000000110000",
40799 => "0111000000110000",
40800 => "0111000000110000",
40801 => "0111000000110000",
40802 => "0111000000110000",
40803 => "0111000001000000",
40804 => "0111000001000000",
40805 => "0111000001000000",
40806 => "0111000001000000",
40807 => "0111000001000000",
40808 => "0111000001000000",
40809 => "0111000001000000",
40810 => "0111000001000000",
40811 => "0111000001000000",
40812 => "0111000001000000",
40813 => "0111000001000000",
40814 => "0111000001000000",
40815 => "0111000001000000",
40816 => "0111000001000000",
40817 => "0111000001000000",
40818 => "0111000001000000",
40819 => "0111000001000000",
40820 => "0111000001000000",
40821 => "0111000001010000",
40822 => "0111000001010000",
40823 => "0111000001010000",
40824 => "0111000001010000",
40825 => "0111000001010000",
40826 => "0111000001010000",
40827 => "0111000001010000",
40828 => "0111000001010000",
40829 => "0111000001010000",
40830 => "0111000001010000",
40831 => "0111000001010000",
40832 => "0111000001010000",
40833 => "0111000001010000",
40834 => "0111000001010000",
40835 => "0111000001010000",
40836 => "0111000001010000",
40837 => "0111000001010000",
40838 => "0111000001010000",
40839 => "0111000001010000",
40840 => "0111000001100000",
40841 => "0111000001100000",
40842 => "0111000001100000",
40843 => "0111000001100000",
40844 => "0111000001100000",
40845 => "0111000001100000",
40846 => "0111000001100000",
40847 => "0111000001100000",
40848 => "0111000001100000",
40849 => "0111000001100000",
40850 => "0111000001100000",
40851 => "0111000001100000",
40852 => "0111000001100000",
40853 => "0111000001100000",
40854 => "0111000001100000",
40855 => "0111000001100000",
40856 => "0111000001100000",
40857 => "0111000001100000",
40858 => "0111000001110000",
40859 => "0111000001110000",
40860 => "0111000001110000",
40861 => "0111000001110000",
40862 => "0111000001110000",
40863 => "0111000001110000",
40864 => "0111000001110000",
40865 => "0111000001110000",
40866 => "0111000001110000",
40867 => "0111000001110000",
40868 => "0111000001110000",
40869 => "0111000001110000",
40870 => "0111000001110000",
40871 => "0111000001110000",
40872 => "0111000001110000",
40873 => "0111000001110000",
40874 => "0111000001110000",
40875 => "0111000001110000",
40876 => "0111000001110000",
40877 => "0111000010000000",
40878 => "0111000010000000",
40879 => "0111000010000000",
40880 => "0111000010000000",
40881 => "0111000010000000",
40882 => "0111000010000000",
40883 => "0111000010000000",
40884 => "0111000010000000",
40885 => "0111000010000000",
40886 => "0111000010000000",
40887 => "0111000010000000",
40888 => "0111000010000000",
40889 => "0111000010000000",
40890 => "0111000010000000",
40891 => "0111000010000000",
40892 => "0111000010000000",
40893 => "0111000010000000",
40894 => "0111000010000000",
40895 => "0111000010000000",
40896 => "0111000010010000",
40897 => "0111000010010000",
40898 => "0111000010010000",
40899 => "0111000010010000",
40900 => "0111000010010000",
40901 => "0111000010010000",
40902 => "0111000010010000",
40903 => "0111000010010000",
40904 => "0111000010010000",
40905 => "0111000010010000",
40906 => "0111000010010000",
40907 => "0111000010010000",
40908 => "0111000010010000",
40909 => "0111000010010000",
40910 => "0111000010010000",
40911 => "0111000010010000",
40912 => "0111000010010000",
40913 => "0111000010010000",
40914 => "0111000010010000",
40915 => "0111000010100000",
40916 => "0111000010100000",
40917 => "0111000010100000",
40918 => "0111000010100000",
40919 => "0111000010100000",
40920 => "0111000010100000",
40921 => "0111000010100000",
40922 => "0111000010100000",
40923 => "0111000010100000",
40924 => "0111000010100000",
40925 => "0111000010100000",
40926 => "0111000010100000",
40927 => "0111000010100000",
40928 => "0111000010100000",
40929 => "0111000010100000",
40930 => "0111000010100000",
40931 => "0111000010100000",
40932 => "0111000010100000",
40933 => "0111000010100000",
40934 => "0111000010110000",
40935 => "0111000010110000",
40936 => "0111000010110000",
40937 => "0111000010110000",
40938 => "0111000010110000",
40939 => "0111000010110000",
40940 => "0111000010110000",
40941 => "0111000010110000",
40942 => "0111000010110000",
40943 => "0111000010110000",
40944 => "0111000010110000",
40945 => "0111000010110000",
40946 => "0111000010110000",
40947 => "0111000010110000",
40948 => "0111000010110000",
40949 => "0111000010110000",
40950 => "0111000010110000",
40951 => "0111000010110000",
40952 => "0111000010110000",
40953 => "0111000011000000",
40954 => "0111000011000000",
40955 => "0111000011000000",
40956 => "0111000011000000",
40957 => "0111000011000000",
40958 => "0111000011000000",
40959 => "0111000011000000",
40960 => "0111000011000000",
40961 => "0111000011000000",
40962 => "0111000011000000",
40963 => "0111000011000000",
40964 => "0111000011000000",
40965 => "0111000011000000",
40966 => "0111000011000000",
40967 => "0111000011000000",
40968 => "0111000011000000",
40969 => "0111000011000000",
40970 => "0111000011000000",
40971 => "0111000011000000",
40972 => "0111000011010000",
40973 => "0111000011010000",
40974 => "0111000011010000",
40975 => "0111000011010000",
40976 => "0111000011010000",
40977 => "0111000011010000",
40978 => "0111000011010000",
40979 => "0111000011010000",
40980 => "0111000011010000",
40981 => "0111000011010000",
40982 => "0111000011010000",
40983 => "0111000011010000",
40984 => "0111000011010000",
40985 => "0111000011010000",
40986 => "0111000011010000",
40987 => "0111000011010000",
40988 => "0111000011010000",
40989 => "0111000011010000",
40990 => "0111000011010000",
40991 => "0111000011100000",
40992 => "0111000011100000",
40993 => "0111000011100000",
40994 => "0111000011100000",
40995 => "0111000011100000",
40996 => "0111000011100000",
40997 => "0111000011100000",
40998 => "0111000011100000",
40999 => "0111000011100000",
41000 => "0111000011100000",
41001 => "0111000011100000",
41002 => "0111000011100000",
41003 => "0111000011100000",
41004 => "0111000011100000",
41005 => "0111000011100000",
41006 => "0111000011100000",
41007 => "0111000011100000",
41008 => "0111000011100000",
41009 => "0111000011100000",
41010 => "0111000011110000",
41011 => "0111000011110000",
41012 => "0111000011110000",
41013 => "0111000011110000",
41014 => "0111000011110000",
41015 => "0111000011110000",
41016 => "0111000011110000",
41017 => "0111000011110000",
41018 => "0111000011110000",
41019 => "0111000011110000",
41020 => "0111000011110000",
41021 => "0111000011110000",
41022 => "0111000011110000",
41023 => "0111000011110000",
41024 => "0111000011110000",
41025 => "0111000011110000",
41026 => "0111000011110000",
41027 => "0111000011110000",
41028 => "0111000011110000",
41029 => "0111000100000000",
41030 => "0111000100000000",
41031 => "0111000100000000",
41032 => "0111000100000000",
41033 => "0111000100000000",
41034 => "0111000100000000",
41035 => "0111000100000000",
41036 => "0111000100000000",
41037 => "0111000100000000",
41038 => "0111000100000000",
41039 => "0111000100000000",
41040 => "0111000100000000",
41041 => "0111000100000000",
41042 => "0111000100000000",
41043 => "0111000100000000",
41044 => "0111000100000000",
41045 => "0111000100000000",
41046 => "0111000100000000",
41047 => "0111000100000000",
41048 => "0111000100000000",
41049 => "0111000100010000",
41050 => "0111000100010000",
41051 => "0111000100010000",
41052 => "0111000100010000",
41053 => "0111000100010000",
41054 => "0111000100010000",
41055 => "0111000100010000",
41056 => "0111000100010000",
41057 => "0111000100010000",
41058 => "0111000100010000",
41059 => "0111000100010000",
41060 => "0111000100010000",
41061 => "0111000100010000",
41062 => "0111000100010000",
41063 => "0111000100010000",
41064 => "0111000100010000",
41065 => "0111000100010000",
41066 => "0111000100010000",
41067 => "0111000100010000",
41068 => "0111000100100000",
41069 => "0111000100100000",
41070 => "0111000100100000",
41071 => "0111000100100000",
41072 => "0111000100100000",
41073 => "0111000100100000",
41074 => "0111000100100000",
41075 => "0111000100100000",
41076 => "0111000100100000",
41077 => "0111000100100000",
41078 => "0111000100100000",
41079 => "0111000100100000",
41080 => "0111000100100000",
41081 => "0111000100100000",
41082 => "0111000100100000",
41083 => "0111000100100000",
41084 => "0111000100100000",
41085 => "0111000100100000",
41086 => "0111000100100000",
41087 => "0111000100100000",
41088 => "0111000100110000",
41089 => "0111000100110000",
41090 => "0111000100110000",
41091 => "0111000100110000",
41092 => "0111000100110000",
41093 => "0111000100110000",
41094 => "0111000100110000",
41095 => "0111000100110000",
41096 => "0111000100110000",
41097 => "0111000100110000",
41098 => "0111000100110000",
41099 => "0111000100110000",
41100 => "0111000100110000",
41101 => "0111000100110000",
41102 => "0111000100110000",
41103 => "0111000100110000",
41104 => "0111000100110000",
41105 => "0111000100110000",
41106 => "0111000100110000",
41107 => "0111000101000000",
41108 => "0111000101000000",
41109 => "0111000101000000",
41110 => "0111000101000000",
41111 => "0111000101000000",
41112 => "0111000101000000",
41113 => "0111000101000000",
41114 => "0111000101000000",
41115 => "0111000101000000",
41116 => "0111000101000000",
41117 => "0111000101000000",
41118 => "0111000101000000",
41119 => "0111000101000000",
41120 => "0111000101000000",
41121 => "0111000101000000",
41122 => "0111000101000000",
41123 => "0111000101000000",
41124 => "0111000101000000",
41125 => "0111000101000000",
41126 => "0111000101000000",
41127 => "0111000101010000",
41128 => "0111000101010000",
41129 => "0111000101010000",
41130 => "0111000101010000",
41131 => "0111000101010000",
41132 => "0111000101010000",
41133 => "0111000101010000",
41134 => "0111000101010000",
41135 => "0111000101010000",
41136 => "0111000101010000",
41137 => "0111000101010000",
41138 => "0111000101010000",
41139 => "0111000101010000",
41140 => "0111000101010000",
41141 => "0111000101010000",
41142 => "0111000101010000",
41143 => "0111000101010000",
41144 => "0111000101010000",
41145 => "0111000101010000",
41146 => "0111000101100000",
41147 => "0111000101100000",
41148 => "0111000101100000",
41149 => "0111000101100000",
41150 => "0111000101100000",
41151 => "0111000101100000",
41152 => "0111000101100000",
41153 => "0111000101100000",
41154 => "0111000101100000",
41155 => "0111000101100000",
41156 => "0111000101100000",
41157 => "0111000101100000",
41158 => "0111000101100000",
41159 => "0111000101100000",
41160 => "0111000101100000",
41161 => "0111000101100000",
41162 => "0111000101100000",
41163 => "0111000101100000",
41164 => "0111000101100000",
41165 => "0111000101100000",
41166 => "0111000101110000",
41167 => "0111000101110000",
41168 => "0111000101110000",
41169 => "0111000101110000",
41170 => "0111000101110000",
41171 => "0111000101110000",
41172 => "0111000101110000",
41173 => "0111000101110000",
41174 => "0111000101110000",
41175 => "0111000101110000",
41176 => "0111000101110000",
41177 => "0111000101110000",
41178 => "0111000101110000",
41179 => "0111000101110000",
41180 => "0111000101110000",
41181 => "0111000101110000",
41182 => "0111000101110000",
41183 => "0111000101110000",
41184 => "0111000101110000",
41185 => "0111000101110000",
41186 => "0111000110000000",
41187 => "0111000110000000",
41188 => "0111000110000000",
41189 => "0111000110000000",
41190 => "0111000110000000",
41191 => "0111000110000000",
41192 => "0111000110000000",
41193 => "0111000110000000",
41194 => "0111000110000000",
41195 => "0111000110000000",
41196 => "0111000110000000",
41197 => "0111000110000000",
41198 => "0111000110000000",
41199 => "0111000110000000",
41200 => "0111000110000000",
41201 => "0111000110000000",
41202 => "0111000110000000",
41203 => "0111000110000000",
41204 => "0111000110000000",
41205 => "0111000110000000",
41206 => "0111000110010000",
41207 => "0111000110010000",
41208 => "0111000110010000",
41209 => "0111000110010000",
41210 => "0111000110010000",
41211 => "0111000110010000",
41212 => "0111000110010000",
41213 => "0111000110010000",
41214 => "0111000110010000",
41215 => "0111000110010000",
41216 => "0111000110010000",
41217 => "0111000110010000",
41218 => "0111000110010000",
41219 => "0111000110010000",
41220 => "0111000110010000",
41221 => "0111000110010000",
41222 => "0111000110010000",
41223 => "0111000110010000",
41224 => "0111000110010000",
41225 => "0111000110010000",
41226 => "0111000110100000",
41227 => "0111000110100000",
41228 => "0111000110100000",
41229 => "0111000110100000",
41230 => "0111000110100000",
41231 => "0111000110100000",
41232 => "0111000110100000",
41233 => "0111000110100000",
41234 => "0111000110100000",
41235 => "0111000110100000",
41236 => "0111000110100000",
41237 => "0111000110100000",
41238 => "0111000110100000",
41239 => "0111000110100000",
41240 => "0111000110100000",
41241 => "0111000110100000",
41242 => "0111000110100000",
41243 => "0111000110100000",
41244 => "0111000110100000",
41245 => "0111000110100000",
41246 => "0111000110110000",
41247 => "0111000110110000",
41248 => "0111000110110000",
41249 => "0111000110110000",
41250 => "0111000110110000",
41251 => "0111000110110000",
41252 => "0111000110110000",
41253 => "0111000110110000",
41254 => "0111000110110000",
41255 => "0111000110110000",
41256 => "0111000110110000",
41257 => "0111000110110000",
41258 => "0111000110110000",
41259 => "0111000110110000",
41260 => "0111000110110000",
41261 => "0111000110110000",
41262 => "0111000110110000",
41263 => "0111000110110000",
41264 => "0111000110110000",
41265 => "0111000110110000",
41266 => "0111000111000000",
41267 => "0111000111000000",
41268 => "0111000111000000",
41269 => "0111000111000000",
41270 => "0111000111000000",
41271 => "0111000111000000",
41272 => "0111000111000000",
41273 => "0111000111000000",
41274 => "0111000111000000",
41275 => "0111000111000000",
41276 => "0111000111000000",
41277 => "0111000111000000",
41278 => "0111000111000000",
41279 => "0111000111000000",
41280 => "0111000111000000",
41281 => "0111000111000000",
41282 => "0111000111000000",
41283 => "0111000111000000",
41284 => "0111000111000000",
41285 => "0111000111000000",
41286 => "0111000111010000",
41287 => "0111000111010000",
41288 => "0111000111010000",
41289 => "0111000111010000",
41290 => "0111000111010000",
41291 => "0111000111010000",
41292 => "0111000111010000",
41293 => "0111000111010000",
41294 => "0111000111010000",
41295 => "0111000111010000",
41296 => "0111000111010000",
41297 => "0111000111010000",
41298 => "0111000111010000",
41299 => "0111000111010000",
41300 => "0111000111010000",
41301 => "0111000111010000",
41302 => "0111000111010000",
41303 => "0111000111010000",
41304 => "0111000111010000",
41305 => "0111000111010000",
41306 => "0111000111010000",
41307 => "0111000111100000",
41308 => "0111000111100000",
41309 => "0111000111100000",
41310 => "0111000111100000",
41311 => "0111000111100000",
41312 => "0111000111100000",
41313 => "0111000111100000",
41314 => "0111000111100000",
41315 => "0111000111100000",
41316 => "0111000111100000",
41317 => "0111000111100000",
41318 => "0111000111100000",
41319 => "0111000111100000",
41320 => "0111000111100000",
41321 => "0111000111100000",
41322 => "0111000111100000",
41323 => "0111000111100000",
41324 => "0111000111100000",
41325 => "0111000111100000",
41326 => "0111000111100000",
41327 => "0111000111110000",
41328 => "0111000111110000",
41329 => "0111000111110000",
41330 => "0111000111110000",
41331 => "0111000111110000",
41332 => "0111000111110000",
41333 => "0111000111110000",
41334 => "0111000111110000",
41335 => "0111000111110000",
41336 => "0111000111110000",
41337 => "0111000111110000",
41338 => "0111000111110000",
41339 => "0111000111110000",
41340 => "0111000111110000",
41341 => "0111000111110000",
41342 => "0111000111110000",
41343 => "0111000111110000",
41344 => "0111000111110000",
41345 => "0111000111110000",
41346 => "0111000111110000",
41347 => "0111000111110000",
41348 => "0111001000000000",
41349 => "0111001000000000",
41350 => "0111001000000000",
41351 => "0111001000000000",
41352 => "0111001000000000",
41353 => "0111001000000000",
41354 => "0111001000000000",
41355 => "0111001000000000",
41356 => "0111001000000000",
41357 => "0111001000000000",
41358 => "0111001000000000",
41359 => "0111001000000000",
41360 => "0111001000000000",
41361 => "0111001000000000",
41362 => "0111001000000000",
41363 => "0111001000000000",
41364 => "0111001000000000",
41365 => "0111001000000000",
41366 => "0111001000000000",
41367 => "0111001000000000",
41368 => "0111001000010000",
41369 => "0111001000010000",
41370 => "0111001000010000",
41371 => "0111001000010000",
41372 => "0111001000010000",
41373 => "0111001000010000",
41374 => "0111001000010000",
41375 => "0111001000010000",
41376 => "0111001000010000",
41377 => "0111001000010000",
41378 => "0111001000010000",
41379 => "0111001000010000",
41380 => "0111001000010000",
41381 => "0111001000010000",
41382 => "0111001000010000",
41383 => "0111001000010000",
41384 => "0111001000010000",
41385 => "0111001000010000",
41386 => "0111001000010000",
41387 => "0111001000010000",
41388 => "0111001000010000",
41389 => "0111001000100000",
41390 => "0111001000100000",
41391 => "0111001000100000",
41392 => "0111001000100000",
41393 => "0111001000100000",
41394 => "0111001000100000",
41395 => "0111001000100000",
41396 => "0111001000100000",
41397 => "0111001000100000",
41398 => "0111001000100000",
41399 => "0111001000100000",
41400 => "0111001000100000",
41401 => "0111001000100000",
41402 => "0111001000100000",
41403 => "0111001000100000",
41404 => "0111001000100000",
41405 => "0111001000100000",
41406 => "0111001000100000",
41407 => "0111001000100000",
41408 => "0111001000100000",
41409 => "0111001000110000",
41410 => "0111001000110000",
41411 => "0111001000110000",
41412 => "0111001000110000",
41413 => "0111001000110000",
41414 => "0111001000110000",
41415 => "0111001000110000",
41416 => "0111001000110000",
41417 => "0111001000110000",
41418 => "0111001000110000",
41419 => "0111001000110000",
41420 => "0111001000110000",
41421 => "0111001000110000",
41422 => "0111001000110000",
41423 => "0111001000110000",
41424 => "0111001000110000",
41425 => "0111001000110000",
41426 => "0111001000110000",
41427 => "0111001000110000",
41428 => "0111001000110000",
41429 => "0111001000110000",
41430 => "0111001001000000",
41431 => "0111001001000000",
41432 => "0111001001000000",
41433 => "0111001001000000",
41434 => "0111001001000000",
41435 => "0111001001000000",
41436 => "0111001001000000",
41437 => "0111001001000000",
41438 => "0111001001000000",
41439 => "0111001001000000",
41440 => "0111001001000000",
41441 => "0111001001000000",
41442 => "0111001001000000",
41443 => "0111001001000000",
41444 => "0111001001000000",
41445 => "0111001001000000",
41446 => "0111001001000000",
41447 => "0111001001000000",
41448 => "0111001001000000",
41449 => "0111001001000000",
41450 => "0111001001000000",
41451 => "0111001001010000",
41452 => "0111001001010000",
41453 => "0111001001010000",
41454 => "0111001001010000",
41455 => "0111001001010000",
41456 => "0111001001010000",
41457 => "0111001001010000",
41458 => "0111001001010000",
41459 => "0111001001010000",
41460 => "0111001001010000",
41461 => "0111001001010000",
41462 => "0111001001010000",
41463 => "0111001001010000",
41464 => "0111001001010000",
41465 => "0111001001010000",
41466 => "0111001001010000",
41467 => "0111001001010000",
41468 => "0111001001010000",
41469 => "0111001001010000",
41470 => "0111001001010000",
41471 => "0111001001010000",
41472 => "0111001001100000",
41473 => "0111001001100000",
41474 => "0111001001100000",
41475 => "0111001001100000",
41476 => "0111001001100000",
41477 => "0111001001100000",
41478 => "0111001001100000",
41479 => "0111001001100000",
41480 => "0111001001100000",
41481 => "0111001001100000",
41482 => "0111001001100000",
41483 => "0111001001100000",
41484 => "0111001001100000",
41485 => "0111001001100000",
41486 => "0111001001100000",
41487 => "0111001001100000",
41488 => "0111001001100000",
41489 => "0111001001100000",
41490 => "0111001001100000",
41491 => "0111001001100000",
41492 => "0111001001100000",
41493 => "0111001001110000",
41494 => "0111001001110000",
41495 => "0111001001110000",
41496 => "0111001001110000",
41497 => "0111001001110000",
41498 => "0111001001110000",
41499 => "0111001001110000",
41500 => "0111001001110000",
41501 => "0111001001110000",
41502 => "0111001001110000",
41503 => "0111001001110000",
41504 => "0111001001110000",
41505 => "0111001001110000",
41506 => "0111001001110000",
41507 => "0111001001110000",
41508 => "0111001001110000",
41509 => "0111001001110000",
41510 => "0111001001110000",
41511 => "0111001001110000",
41512 => "0111001001110000",
41513 => "0111001001110000",
41514 => "0111001010000000",
41515 => "0111001010000000",
41516 => "0111001010000000",
41517 => "0111001010000000",
41518 => "0111001010000000",
41519 => "0111001010000000",
41520 => "0111001010000000",
41521 => "0111001010000000",
41522 => "0111001010000000",
41523 => "0111001010000000",
41524 => "0111001010000000",
41525 => "0111001010000000",
41526 => "0111001010000000",
41527 => "0111001010000000",
41528 => "0111001010000000",
41529 => "0111001010000000",
41530 => "0111001010000000",
41531 => "0111001010000000",
41532 => "0111001010000000",
41533 => "0111001010000000",
41534 => "0111001010000000",
41535 => "0111001010010000",
41536 => "0111001010010000",
41537 => "0111001010010000",
41538 => "0111001010010000",
41539 => "0111001010010000",
41540 => "0111001010010000",
41541 => "0111001010010000",
41542 => "0111001010010000",
41543 => "0111001010010000",
41544 => "0111001010010000",
41545 => "0111001010010000",
41546 => "0111001010010000",
41547 => "0111001010010000",
41548 => "0111001010010000",
41549 => "0111001010010000",
41550 => "0111001010010000",
41551 => "0111001010010000",
41552 => "0111001010010000",
41553 => "0111001010010000",
41554 => "0111001010010000",
41555 => "0111001010010000",
41556 => "0111001010010000",
41557 => "0111001010100000",
41558 => "0111001010100000",
41559 => "0111001010100000",
41560 => "0111001010100000",
41561 => "0111001010100000",
41562 => "0111001010100000",
41563 => "0111001010100000",
41564 => "0111001010100000",
41565 => "0111001010100000",
41566 => "0111001010100000",
41567 => "0111001010100000",
41568 => "0111001010100000",
41569 => "0111001010100000",
41570 => "0111001010100000",
41571 => "0111001010100000",
41572 => "0111001010100000",
41573 => "0111001010100000",
41574 => "0111001010100000",
41575 => "0111001010100000",
41576 => "0111001010100000",
41577 => "0111001010100000",
41578 => "0111001010110000",
41579 => "0111001010110000",
41580 => "0111001010110000",
41581 => "0111001010110000",
41582 => "0111001010110000",
41583 => "0111001010110000",
41584 => "0111001010110000",
41585 => "0111001010110000",
41586 => "0111001010110000",
41587 => "0111001010110000",
41588 => "0111001010110000",
41589 => "0111001010110000",
41590 => "0111001010110000",
41591 => "0111001010110000",
41592 => "0111001010110000",
41593 => "0111001010110000",
41594 => "0111001010110000",
41595 => "0111001010110000",
41596 => "0111001010110000",
41597 => "0111001010110000",
41598 => "0111001010110000",
41599 => "0111001011000000",
41600 => "0111001011000000",
41601 => "0111001011000000",
41602 => "0111001011000000",
41603 => "0111001011000000",
41604 => "0111001011000000",
41605 => "0111001011000000",
41606 => "0111001011000000",
41607 => "0111001011000000",
41608 => "0111001011000000",
41609 => "0111001011000000",
41610 => "0111001011000000",
41611 => "0111001011000000",
41612 => "0111001011000000",
41613 => "0111001011000000",
41614 => "0111001011000000",
41615 => "0111001011000000",
41616 => "0111001011000000",
41617 => "0111001011000000",
41618 => "0111001011000000",
41619 => "0111001011000000",
41620 => "0111001011000000",
41621 => "0111001011010000",
41622 => "0111001011010000",
41623 => "0111001011010000",
41624 => "0111001011010000",
41625 => "0111001011010000",
41626 => "0111001011010000",
41627 => "0111001011010000",
41628 => "0111001011010000",
41629 => "0111001011010000",
41630 => "0111001011010000",
41631 => "0111001011010000",
41632 => "0111001011010000",
41633 => "0111001011010000",
41634 => "0111001011010000",
41635 => "0111001011010000",
41636 => "0111001011010000",
41637 => "0111001011010000",
41638 => "0111001011010000",
41639 => "0111001011010000",
41640 => "0111001011010000",
41641 => "0111001011010000",
41642 => "0111001011010000",
41643 => "0111001011100000",
41644 => "0111001011100000",
41645 => "0111001011100000",
41646 => "0111001011100000",
41647 => "0111001011100000",
41648 => "0111001011100000",
41649 => "0111001011100000",
41650 => "0111001011100000",
41651 => "0111001011100000",
41652 => "0111001011100000",
41653 => "0111001011100000",
41654 => "0111001011100000",
41655 => "0111001011100000",
41656 => "0111001011100000",
41657 => "0111001011100000",
41658 => "0111001011100000",
41659 => "0111001011100000",
41660 => "0111001011100000",
41661 => "0111001011100000",
41662 => "0111001011100000",
41663 => "0111001011100000",
41664 => "0111001011110000",
41665 => "0111001011110000",
41666 => "0111001011110000",
41667 => "0111001011110000",
41668 => "0111001011110000",
41669 => "0111001011110000",
41670 => "0111001011110000",
41671 => "0111001011110000",
41672 => "0111001011110000",
41673 => "0111001011110000",
41674 => "0111001011110000",
41675 => "0111001011110000",
41676 => "0111001011110000",
41677 => "0111001011110000",
41678 => "0111001011110000",
41679 => "0111001011110000",
41680 => "0111001011110000",
41681 => "0111001011110000",
41682 => "0111001011110000",
41683 => "0111001011110000",
41684 => "0111001011110000",
41685 => "0111001011110000",
41686 => "0111001100000000",
41687 => "0111001100000000",
41688 => "0111001100000000",
41689 => "0111001100000000",
41690 => "0111001100000000",
41691 => "0111001100000000",
41692 => "0111001100000000",
41693 => "0111001100000000",
41694 => "0111001100000000",
41695 => "0111001100000000",
41696 => "0111001100000000",
41697 => "0111001100000000",
41698 => "0111001100000000",
41699 => "0111001100000000",
41700 => "0111001100000000",
41701 => "0111001100000000",
41702 => "0111001100000000",
41703 => "0111001100000000",
41704 => "0111001100000000",
41705 => "0111001100000000",
41706 => "0111001100000000",
41707 => "0111001100000000",
41708 => "0111001100010000",
41709 => "0111001100010000",
41710 => "0111001100010000",
41711 => "0111001100010000",
41712 => "0111001100010000",
41713 => "0111001100010000",
41714 => "0111001100010000",
41715 => "0111001100010000",
41716 => "0111001100010000",
41717 => "0111001100010000",
41718 => "0111001100010000",
41719 => "0111001100010000",
41720 => "0111001100010000",
41721 => "0111001100010000",
41722 => "0111001100010000",
41723 => "0111001100010000",
41724 => "0111001100010000",
41725 => "0111001100010000",
41726 => "0111001100010000",
41727 => "0111001100010000",
41728 => "0111001100010000",
41729 => "0111001100010000",
41730 => "0111001100100000",
41731 => "0111001100100000",
41732 => "0111001100100000",
41733 => "0111001100100000",
41734 => "0111001100100000",
41735 => "0111001100100000",
41736 => "0111001100100000",
41737 => "0111001100100000",
41738 => "0111001100100000",
41739 => "0111001100100000",
41740 => "0111001100100000",
41741 => "0111001100100000",
41742 => "0111001100100000",
41743 => "0111001100100000",
41744 => "0111001100100000",
41745 => "0111001100100000",
41746 => "0111001100100000",
41747 => "0111001100100000",
41748 => "0111001100100000",
41749 => "0111001100100000",
41750 => "0111001100100000",
41751 => "0111001100100000",
41752 => "0111001100110000",
41753 => "0111001100110000",
41754 => "0111001100110000",
41755 => "0111001100110000",
41756 => "0111001100110000",
41757 => "0111001100110000",
41758 => "0111001100110000",
41759 => "0111001100110000",
41760 => "0111001100110000",
41761 => "0111001100110000",
41762 => "0111001100110000",
41763 => "0111001100110000",
41764 => "0111001100110000",
41765 => "0111001100110000",
41766 => "0111001100110000",
41767 => "0111001100110000",
41768 => "0111001100110000",
41769 => "0111001100110000",
41770 => "0111001100110000",
41771 => "0111001100110000",
41772 => "0111001100110000",
41773 => "0111001100110000",
41774 => "0111001101000000",
41775 => "0111001101000000",
41776 => "0111001101000000",
41777 => "0111001101000000",
41778 => "0111001101000000",
41779 => "0111001101000000",
41780 => "0111001101000000",
41781 => "0111001101000000",
41782 => "0111001101000000",
41783 => "0111001101000000",
41784 => "0111001101000000",
41785 => "0111001101000000",
41786 => "0111001101000000",
41787 => "0111001101000000",
41788 => "0111001101000000",
41789 => "0111001101000000",
41790 => "0111001101000000",
41791 => "0111001101000000",
41792 => "0111001101000000",
41793 => "0111001101000000",
41794 => "0111001101000000",
41795 => "0111001101000000",
41796 => "0111001101000000",
41797 => "0111001101010000",
41798 => "0111001101010000",
41799 => "0111001101010000",
41800 => "0111001101010000",
41801 => "0111001101010000",
41802 => "0111001101010000",
41803 => "0111001101010000",
41804 => "0111001101010000",
41805 => "0111001101010000",
41806 => "0111001101010000",
41807 => "0111001101010000",
41808 => "0111001101010000",
41809 => "0111001101010000",
41810 => "0111001101010000",
41811 => "0111001101010000",
41812 => "0111001101010000",
41813 => "0111001101010000",
41814 => "0111001101010000",
41815 => "0111001101010000",
41816 => "0111001101010000",
41817 => "0111001101010000",
41818 => "0111001101010000",
41819 => "0111001101100000",
41820 => "0111001101100000",
41821 => "0111001101100000",
41822 => "0111001101100000",
41823 => "0111001101100000",
41824 => "0111001101100000",
41825 => "0111001101100000",
41826 => "0111001101100000",
41827 => "0111001101100000",
41828 => "0111001101100000",
41829 => "0111001101100000",
41830 => "0111001101100000",
41831 => "0111001101100000",
41832 => "0111001101100000",
41833 => "0111001101100000",
41834 => "0111001101100000",
41835 => "0111001101100000",
41836 => "0111001101100000",
41837 => "0111001101100000",
41838 => "0111001101100000",
41839 => "0111001101100000",
41840 => "0111001101100000",
41841 => "0111001101100000",
41842 => "0111001101110000",
41843 => "0111001101110000",
41844 => "0111001101110000",
41845 => "0111001101110000",
41846 => "0111001101110000",
41847 => "0111001101110000",
41848 => "0111001101110000",
41849 => "0111001101110000",
41850 => "0111001101110000",
41851 => "0111001101110000",
41852 => "0111001101110000",
41853 => "0111001101110000",
41854 => "0111001101110000",
41855 => "0111001101110000",
41856 => "0111001101110000",
41857 => "0111001101110000",
41858 => "0111001101110000",
41859 => "0111001101110000",
41860 => "0111001101110000",
41861 => "0111001101110000",
41862 => "0111001101110000",
41863 => "0111001101110000",
41864 => "0111001110000000",
41865 => "0111001110000000",
41866 => "0111001110000000",
41867 => "0111001110000000",
41868 => "0111001110000000",
41869 => "0111001110000000",
41870 => "0111001110000000",
41871 => "0111001110000000",
41872 => "0111001110000000",
41873 => "0111001110000000",
41874 => "0111001110000000",
41875 => "0111001110000000",
41876 => "0111001110000000",
41877 => "0111001110000000",
41878 => "0111001110000000",
41879 => "0111001110000000",
41880 => "0111001110000000",
41881 => "0111001110000000",
41882 => "0111001110000000",
41883 => "0111001110000000",
41884 => "0111001110000000",
41885 => "0111001110000000",
41886 => "0111001110000000",
41887 => "0111001110010000",
41888 => "0111001110010000",
41889 => "0111001110010000",
41890 => "0111001110010000",
41891 => "0111001110010000",
41892 => "0111001110010000",
41893 => "0111001110010000",
41894 => "0111001110010000",
41895 => "0111001110010000",
41896 => "0111001110010000",
41897 => "0111001110010000",
41898 => "0111001110010000",
41899 => "0111001110010000",
41900 => "0111001110010000",
41901 => "0111001110010000",
41902 => "0111001110010000",
41903 => "0111001110010000",
41904 => "0111001110010000",
41905 => "0111001110010000",
41906 => "0111001110010000",
41907 => "0111001110010000",
41908 => "0111001110010000",
41909 => "0111001110010000",
41910 => "0111001110100000",
41911 => "0111001110100000",
41912 => "0111001110100000",
41913 => "0111001110100000",
41914 => "0111001110100000",
41915 => "0111001110100000",
41916 => "0111001110100000",
41917 => "0111001110100000",
41918 => "0111001110100000",
41919 => "0111001110100000",
41920 => "0111001110100000",
41921 => "0111001110100000",
41922 => "0111001110100000",
41923 => "0111001110100000",
41924 => "0111001110100000",
41925 => "0111001110100000",
41926 => "0111001110100000",
41927 => "0111001110100000",
41928 => "0111001110100000",
41929 => "0111001110100000",
41930 => "0111001110100000",
41931 => "0111001110100000",
41932 => "0111001110100000",
41933 => "0111001110110000",
41934 => "0111001110110000",
41935 => "0111001110110000",
41936 => "0111001110110000",
41937 => "0111001110110000",
41938 => "0111001110110000",
41939 => "0111001110110000",
41940 => "0111001110110000",
41941 => "0111001110110000",
41942 => "0111001110110000",
41943 => "0111001110110000",
41944 => "0111001110110000",
41945 => "0111001110110000",
41946 => "0111001110110000",
41947 => "0111001110110000",
41948 => "0111001110110000",
41949 => "0111001110110000",
41950 => "0111001110110000",
41951 => "0111001110110000",
41952 => "0111001110110000",
41953 => "0111001110110000",
41954 => "0111001110110000",
41955 => "0111001110110000",
41956 => "0111001111000000",
41957 => "0111001111000000",
41958 => "0111001111000000",
41959 => "0111001111000000",
41960 => "0111001111000000",
41961 => "0111001111000000",
41962 => "0111001111000000",
41963 => "0111001111000000",
41964 => "0111001111000000",
41965 => "0111001111000000",
41966 => "0111001111000000",
41967 => "0111001111000000",
41968 => "0111001111000000",
41969 => "0111001111000000",
41970 => "0111001111000000",
41971 => "0111001111000000",
41972 => "0111001111000000",
41973 => "0111001111000000",
41974 => "0111001111000000",
41975 => "0111001111000000",
41976 => "0111001111000000",
41977 => "0111001111000000",
41978 => "0111001111000000",
41979 => "0111001111010000",
41980 => "0111001111010000",
41981 => "0111001111010000",
41982 => "0111001111010000",
41983 => "0111001111010000",
41984 => "0111001111010000",
41985 => "0111001111010000",
41986 => "0111001111010000",
41987 => "0111001111010000",
41988 => "0111001111010000",
41989 => "0111001111010000",
41990 => "0111001111010000",
41991 => "0111001111010000",
41992 => "0111001111010000",
41993 => "0111001111010000",
41994 => "0111001111010000",
41995 => "0111001111010000",
41996 => "0111001111010000",
41997 => "0111001111010000",
41998 => "0111001111010000",
41999 => "0111001111010000",
42000 => "0111001111010000",
42001 => "0111001111010000",
42002 => "0111001111100000",
42003 => "0111001111100000",
42004 => "0111001111100000",
42005 => "0111001111100000",
42006 => "0111001111100000",
42007 => "0111001111100000",
42008 => "0111001111100000",
42009 => "0111001111100000",
42010 => "0111001111100000",
42011 => "0111001111100000",
42012 => "0111001111100000",
42013 => "0111001111100000",
42014 => "0111001111100000",
42015 => "0111001111100000",
42016 => "0111001111100000",
42017 => "0111001111100000",
42018 => "0111001111100000",
42019 => "0111001111100000",
42020 => "0111001111100000",
42021 => "0111001111100000",
42022 => "0111001111100000",
42023 => "0111001111100000",
42024 => "0111001111100000",
42025 => "0111001111110000",
42026 => "0111001111110000",
42027 => "0111001111110000",
42028 => "0111001111110000",
42029 => "0111001111110000",
42030 => "0111001111110000",
42031 => "0111001111110000",
42032 => "0111001111110000",
42033 => "0111001111110000",
42034 => "0111001111110000",
42035 => "0111001111110000",
42036 => "0111001111110000",
42037 => "0111001111110000",
42038 => "0111001111110000",
42039 => "0111001111110000",
42040 => "0111001111110000",
42041 => "0111001111110000",
42042 => "0111001111110000",
42043 => "0111001111110000",
42044 => "0111001111110000",
42045 => "0111001111110000",
42046 => "0111001111110000",
42047 => "0111001111110000",
42048 => "0111001111110000",
42049 => "0111010000000000",
42050 => "0111010000000000",
42051 => "0111010000000000",
42052 => "0111010000000000",
42053 => "0111010000000000",
42054 => "0111010000000000",
42055 => "0111010000000000",
42056 => "0111010000000000",
42057 => "0111010000000000",
42058 => "0111010000000000",
42059 => "0111010000000000",
42060 => "0111010000000000",
42061 => "0111010000000000",
42062 => "0111010000000000",
42063 => "0111010000000000",
42064 => "0111010000000000",
42065 => "0111010000000000",
42066 => "0111010000000000",
42067 => "0111010000000000",
42068 => "0111010000000000",
42069 => "0111010000000000",
42070 => "0111010000000000",
42071 => "0111010000000000",
42072 => "0111010000010000",
42073 => "0111010000010000",
42074 => "0111010000010000",
42075 => "0111010000010000",
42076 => "0111010000010000",
42077 => "0111010000010000",
42078 => "0111010000010000",
42079 => "0111010000010000",
42080 => "0111010000010000",
42081 => "0111010000010000",
42082 => "0111010000010000",
42083 => "0111010000010000",
42084 => "0111010000010000",
42085 => "0111010000010000",
42086 => "0111010000010000",
42087 => "0111010000010000",
42088 => "0111010000010000",
42089 => "0111010000010000",
42090 => "0111010000010000",
42091 => "0111010000010000",
42092 => "0111010000010000",
42093 => "0111010000010000",
42094 => "0111010000010000",
42095 => "0111010000010000",
42096 => "0111010000100000",
42097 => "0111010000100000",
42098 => "0111010000100000",
42099 => "0111010000100000",
42100 => "0111010000100000",
42101 => "0111010000100000",
42102 => "0111010000100000",
42103 => "0111010000100000",
42104 => "0111010000100000",
42105 => "0111010000100000",
42106 => "0111010000100000",
42107 => "0111010000100000",
42108 => "0111010000100000",
42109 => "0111010000100000",
42110 => "0111010000100000",
42111 => "0111010000100000",
42112 => "0111010000100000",
42113 => "0111010000100000",
42114 => "0111010000100000",
42115 => "0111010000100000",
42116 => "0111010000100000",
42117 => "0111010000100000",
42118 => "0111010000100000",
42119 => "0111010000100000",
42120 => "0111010000110000",
42121 => "0111010000110000",
42122 => "0111010000110000",
42123 => "0111010000110000",
42124 => "0111010000110000",
42125 => "0111010000110000",
42126 => "0111010000110000",
42127 => "0111010000110000",
42128 => "0111010000110000",
42129 => "0111010000110000",
42130 => "0111010000110000",
42131 => "0111010000110000",
42132 => "0111010000110000",
42133 => "0111010000110000",
42134 => "0111010000110000",
42135 => "0111010000110000",
42136 => "0111010000110000",
42137 => "0111010000110000",
42138 => "0111010000110000",
42139 => "0111010000110000",
42140 => "0111010000110000",
42141 => "0111010000110000",
42142 => "0111010000110000",
42143 => "0111010001000000",
42144 => "0111010001000000",
42145 => "0111010001000000",
42146 => "0111010001000000",
42147 => "0111010001000000",
42148 => "0111010001000000",
42149 => "0111010001000000",
42150 => "0111010001000000",
42151 => "0111010001000000",
42152 => "0111010001000000",
42153 => "0111010001000000",
42154 => "0111010001000000",
42155 => "0111010001000000",
42156 => "0111010001000000",
42157 => "0111010001000000",
42158 => "0111010001000000",
42159 => "0111010001000000",
42160 => "0111010001000000",
42161 => "0111010001000000",
42162 => "0111010001000000",
42163 => "0111010001000000",
42164 => "0111010001000000",
42165 => "0111010001000000",
42166 => "0111010001000000",
42167 => "0111010001010000",
42168 => "0111010001010000",
42169 => "0111010001010000",
42170 => "0111010001010000",
42171 => "0111010001010000",
42172 => "0111010001010000",
42173 => "0111010001010000",
42174 => "0111010001010000",
42175 => "0111010001010000",
42176 => "0111010001010000",
42177 => "0111010001010000",
42178 => "0111010001010000",
42179 => "0111010001010000",
42180 => "0111010001010000",
42181 => "0111010001010000",
42182 => "0111010001010000",
42183 => "0111010001010000",
42184 => "0111010001010000",
42185 => "0111010001010000",
42186 => "0111010001010000",
42187 => "0111010001010000",
42188 => "0111010001010000",
42189 => "0111010001010000",
42190 => "0111010001010000",
42191 => "0111010001010000",
42192 => "0111010001100000",
42193 => "0111010001100000",
42194 => "0111010001100000",
42195 => "0111010001100000",
42196 => "0111010001100000",
42197 => "0111010001100000",
42198 => "0111010001100000",
42199 => "0111010001100000",
42200 => "0111010001100000",
42201 => "0111010001100000",
42202 => "0111010001100000",
42203 => "0111010001100000",
42204 => "0111010001100000",
42205 => "0111010001100000",
42206 => "0111010001100000",
42207 => "0111010001100000",
42208 => "0111010001100000",
42209 => "0111010001100000",
42210 => "0111010001100000",
42211 => "0111010001100000",
42212 => "0111010001100000",
42213 => "0111010001100000",
42214 => "0111010001100000",
42215 => "0111010001100000",
42216 => "0111010001110000",
42217 => "0111010001110000",
42218 => "0111010001110000",
42219 => "0111010001110000",
42220 => "0111010001110000",
42221 => "0111010001110000",
42222 => "0111010001110000",
42223 => "0111010001110000",
42224 => "0111010001110000",
42225 => "0111010001110000",
42226 => "0111010001110000",
42227 => "0111010001110000",
42228 => "0111010001110000",
42229 => "0111010001110000",
42230 => "0111010001110000",
42231 => "0111010001110000",
42232 => "0111010001110000",
42233 => "0111010001110000",
42234 => "0111010001110000",
42235 => "0111010001110000",
42236 => "0111010001110000",
42237 => "0111010001110000",
42238 => "0111010001110000",
42239 => "0111010001110000",
42240 => "0111010010000000",
42241 => "0111010010000000",
42242 => "0111010010000000",
42243 => "0111010010000000",
42244 => "0111010010000000",
42245 => "0111010010000000",
42246 => "0111010010000000",
42247 => "0111010010000000",
42248 => "0111010010000000",
42249 => "0111010010000000",
42250 => "0111010010000000",
42251 => "0111010010000000",
42252 => "0111010010000000",
42253 => "0111010010000000",
42254 => "0111010010000000",
42255 => "0111010010000000",
42256 => "0111010010000000",
42257 => "0111010010000000",
42258 => "0111010010000000",
42259 => "0111010010000000",
42260 => "0111010010000000",
42261 => "0111010010000000",
42262 => "0111010010000000",
42263 => "0111010010000000",
42264 => "0111010010000000",
42265 => "0111010010010000",
42266 => "0111010010010000",
42267 => "0111010010010000",
42268 => "0111010010010000",
42269 => "0111010010010000",
42270 => "0111010010010000",
42271 => "0111010010010000",
42272 => "0111010010010000",
42273 => "0111010010010000",
42274 => "0111010010010000",
42275 => "0111010010010000",
42276 => "0111010010010000",
42277 => "0111010010010000",
42278 => "0111010010010000",
42279 => "0111010010010000",
42280 => "0111010010010000",
42281 => "0111010010010000",
42282 => "0111010010010000",
42283 => "0111010010010000",
42284 => "0111010010010000",
42285 => "0111010010010000",
42286 => "0111010010010000",
42287 => "0111010010010000",
42288 => "0111010010010000",
42289 => "0111010010100000",
42290 => "0111010010100000",
42291 => "0111010010100000",
42292 => "0111010010100000",
42293 => "0111010010100000",
42294 => "0111010010100000",
42295 => "0111010010100000",
42296 => "0111010010100000",
42297 => "0111010010100000",
42298 => "0111010010100000",
42299 => "0111010010100000",
42300 => "0111010010100000",
42301 => "0111010010100000",
42302 => "0111010010100000",
42303 => "0111010010100000",
42304 => "0111010010100000",
42305 => "0111010010100000",
42306 => "0111010010100000",
42307 => "0111010010100000",
42308 => "0111010010100000",
42309 => "0111010010100000",
42310 => "0111010010100000",
42311 => "0111010010100000",
42312 => "0111010010100000",
42313 => "0111010010100000",
42314 => "0111010010110000",
42315 => "0111010010110000",
42316 => "0111010010110000",
42317 => "0111010010110000",
42318 => "0111010010110000",
42319 => "0111010010110000",
42320 => "0111010010110000",
42321 => "0111010010110000",
42322 => "0111010010110000",
42323 => "0111010010110000",
42324 => "0111010010110000",
42325 => "0111010010110000",
42326 => "0111010010110000",
42327 => "0111010010110000",
42328 => "0111010010110000",
42329 => "0111010010110000",
42330 => "0111010010110000",
42331 => "0111010010110000",
42332 => "0111010010110000",
42333 => "0111010010110000",
42334 => "0111010010110000",
42335 => "0111010010110000",
42336 => "0111010010110000",
42337 => "0111010010110000",
42338 => "0111010010110000",
42339 => "0111010011000000",
42340 => "0111010011000000",
42341 => "0111010011000000",
42342 => "0111010011000000",
42343 => "0111010011000000",
42344 => "0111010011000000",
42345 => "0111010011000000",
42346 => "0111010011000000",
42347 => "0111010011000000",
42348 => "0111010011000000",
42349 => "0111010011000000",
42350 => "0111010011000000",
42351 => "0111010011000000",
42352 => "0111010011000000",
42353 => "0111010011000000",
42354 => "0111010011000000",
42355 => "0111010011000000",
42356 => "0111010011000000",
42357 => "0111010011000000",
42358 => "0111010011000000",
42359 => "0111010011000000",
42360 => "0111010011000000",
42361 => "0111010011000000",
42362 => "0111010011000000",
42363 => "0111010011000000",
42364 => "0111010011010000",
42365 => "0111010011010000",
42366 => "0111010011010000",
42367 => "0111010011010000",
42368 => "0111010011010000",
42369 => "0111010011010000",
42370 => "0111010011010000",
42371 => "0111010011010000",
42372 => "0111010011010000",
42373 => "0111010011010000",
42374 => "0111010011010000",
42375 => "0111010011010000",
42376 => "0111010011010000",
42377 => "0111010011010000",
42378 => "0111010011010000",
42379 => "0111010011010000",
42380 => "0111010011010000",
42381 => "0111010011010000",
42382 => "0111010011010000",
42383 => "0111010011010000",
42384 => "0111010011010000",
42385 => "0111010011010000",
42386 => "0111010011010000",
42387 => "0111010011010000",
42388 => "0111010011010000",
42389 => "0111010011100000",
42390 => "0111010011100000",
42391 => "0111010011100000",
42392 => "0111010011100000",
42393 => "0111010011100000",
42394 => "0111010011100000",
42395 => "0111010011100000",
42396 => "0111010011100000",
42397 => "0111010011100000",
42398 => "0111010011100000",
42399 => "0111010011100000",
42400 => "0111010011100000",
42401 => "0111010011100000",
42402 => "0111010011100000",
42403 => "0111010011100000",
42404 => "0111010011100000",
42405 => "0111010011100000",
42406 => "0111010011100000",
42407 => "0111010011100000",
42408 => "0111010011100000",
42409 => "0111010011100000",
42410 => "0111010011100000",
42411 => "0111010011100000",
42412 => "0111010011100000",
42413 => "0111010011100000",
42414 => "0111010011110000",
42415 => "0111010011110000",
42416 => "0111010011110000",
42417 => "0111010011110000",
42418 => "0111010011110000",
42419 => "0111010011110000",
42420 => "0111010011110000",
42421 => "0111010011110000",
42422 => "0111010011110000",
42423 => "0111010011110000",
42424 => "0111010011110000",
42425 => "0111010011110000",
42426 => "0111010011110000",
42427 => "0111010011110000",
42428 => "0111010011110000",
42429 => "0111010011110000",
42430 => "0111010011110000",
42431 => "0111010011110000",
42432 => "0111010011110000",
42433 => "0111010011110000",
42434 => "0111010011110000",
42435 => "0111010011110000",
42436 => "0111010011110000",
42437 => "0111010011110000",
42438 => "0111010011110000",
42439 => "0111010100000000",
42440 => "0111010100000000",
42441 => "0111010100000000",
42442 => "0111010100000000",
42443 => "0111010100000000",
42444 => "0111010100000000",
42445 => "0111010100000000",
42446 => "0111010100000000",
42447 => "0111010100000000",
42448 => "0111010100000000",
42449 => "0111010100000000",
42450 => "0111010100000000",
42451 => "0111010100000000",
42452 => "0111010100000000",
42453 => "0111010100000000",
42454 => "0111010100000000",
42455 => "0111010100000000",
42456 => "0111010100000000",
42457 => "0111010100000000",
42458 => "0111010100000000",
42459 => "0111010100000000",
42460 => "0111010100000000",
42461 => "0111010100000000",
42462 => "0111010100000000",
42463 => "0111010100000000",
42464 => "0111010100000000",
42465 => "0111010100010000",
42466 => "0111010100010000",
42467 => "0111010100010000",
42468 => "0111010100010000",
42469 => "0111010100010000",
42470 => "0111010100010000",
42471 => "0111010100010000",
42472 => "0111010100010000",
42473 => "0111010100010000",
42474 => "0111010100010000",
42475 => "0111010100010000",
42476 => "0111010100010000",
42477 => "0111010100010000",
42478 => "0111010100010000",
42479 => "0111010100010000",
42480 => "0111010100010000",
42481 => "0111010100010000",
42482 => "0111010100010000",
42483 => "0111010100010000",
42484 => "0111010100010000",
42485 => "0111010100010000",
42486 => "0111010100010000",
42487 => "0111010100010000",
42488 => "0111010100010000",
42489 => "0111010100010000",
42490 => "0111010100100000",
42491 => "0111010100100000",
42492 => "0111010100100000",
42493 => "0111010100100000",
42494 => "0111010100100000",
42495 => "0111010100100000",
42496 => "0111010100100000",
42497 => "0111010100100000",
42498 => "0111010100100000",
42499 => "0111010100100000",
42500 => "0111010100100000",
42501 => "0111010100100000",
42502 => "0111010100100000",
42503 => "0111010100100000",
42504 => "0111010100100000",
42505 => "0111010100100000",
42506 => "0111010100100000",
42507 => "0111010100100000",
42508 => "0111010100100000",
42509 => "0111010100100000",
42510 => "0111010100100000",
42511 => "0111010100100000",
42512 => "0111010100100000",
42513 => "0111010100100000",
42514 => "0111010100100000",
42515 => "0111010100100000",
42516 => "0111010100110000",
42517 => "0111010100110000",
42518 => "0111010100110000",
42519 => "0111010100110000",
42520 => "0111010100110000",
42521 => "0111010100110000",
42522 => "0111010100110000",
42523 => "0111010100110000",
42524 => "0111010100110000",
42525 => "0111010100110000",
42526 => "0111010100110000",
42527 => "0111010100110000",
42528 => "0111010100110000",
42529 => "0111010100110000",
42530 => "0111010100110000",
42531 => "0111010100110000",
42532 => "0111010100110000",
42533 => "0111010100110000",
42534 => "0111010100110000",
42535 => "0111010100110000",
42536 => "0111010100110000",
42537 => "0111010100110000",
42538 => "0111010100110000",
42539 => "0111010100110000",
42540 => "0111010100110000",
42541 => "0111010100110000",
42542 => "0111010101000000",
42543 => "0111010101000000",
42544 => "0111010101000000",
42545 => "0111010101000000",
42546 => "0111010101000000",
42547 => "0111010101000000",
42548 => "0111010101000000",
42549 => "0111010101000000",
42550 => "0111010101000000",
42551 => "0111010101000000",
42552 => "0111010101000000",
42553 => "0111010101000000",
42554 => "0111010101000000",
42555 => "0111010101000000",
42556 => "0111010101000000",
42557 => "0111010101000000",
42558 => "0111010101000000",
42559 => "0111010101000000",
42560 => "0111010101000000",
42561 => "0111010101000000",
42562 => "0111010101000000",
42563 => "0111010101000000",
42564 => "0111010101000000",
42565 => "0111010101000000",
42566 => "0111010101000000",
42567 => "0111010101000000",
42568 => "0111010101010000",
42569 => "0111010101010000",
42570 => "0111010101010000",
42571 => "0111010101010000",
42572 => "0111010101010000",
42573 => "0111010101010000",
42574 => "0111010101010000",
42575 => "0111010101010000",
42576 => "0111010101010000",
42577 => "0111010101010000",
42578 => "0111010101010000",
42579 => "0111010101010000",
42580 => "0111010101010000",
42581 => "0111010101010000",
42582 => "0111010101010000",
42583 => "0111010101010000",
42584 => "0111010101010000",
42585 => "0111010101010000",
42586 => "0111010101010000",
42587 => "0111010101010000",
42588 => "0111010101010000",
42589 => "0111010101010000",
42590 => "0111010101010000",
42591 => "0111010101010000",
42592 => "0111010101010000",
42593 => "0111010101010000",
42594 => "0111010101100000",
42595 => "0111010101100000",
42596 => "0111010101100000",
42597 => "0111010101100000",
42598 => "0111010101100000",
42599 => "0111010101100000",
42600 => "0111010101100000",
42601 => "0111010101100000",
42602 => "0111010101100000",
42603 => "0111010101100000",
42604 => "0111010101100000",
42605 => "0111010101100000",
42606 => "0111010101100000",
42607 => "0111010101100000",
42608 => "0111010101100000",
42609 => "0111010101100000",
42610 => "0111010101100000",
42611 => "0111010101100000",
42612 => "0111010101100000",
42613 => "0111010101100000",
42614 => "0111010101100000",
42615 => "0111010101100000",
42616 => "0111010101100000",
42617 => "0111010101100000",
42618 => "0111010101100000",
42619 => "0111010101100000",
42620 => "0111010101110000",
42621 => "0111010101110000",
42622 => "0111010101110000",
42623 => "0111010101110000",
42624 => "0111010101110000",
42625 => "0111010101110000",
42626 => "0111010101110000",
42627 => "0111010101110000",
42628 => "0111010101110000",
42629 => "0111010101110000",
42630 => "0111010101110000",
42631 => "0111010101110000",
42632 => "0111010101110000",
42633 => "0111010101110000",
42634 => "0111010101110000",
42635 => "0111010101110000",
42636 => "0111010101110000",
42637 => "0111010101110000",
42638 => "0111010101110000",
42639 => "0111010101110000",
42640 => "0111010101110000",
42641 => "0111010101110000",
42642 => "0111010101110000",
42643 => "0111010101110000",
42644 => "0111010101110000",
42645 => "0111010101110000",
42646 => "0111010101110000",
42647 => "0111010110000000",
42648 => "0111010110000000",
42649 => "0111010110000000",
42650 => "0111010110000000",
42651 => "0111010110000000",
42652 => "0111010110000000",
42653 => "0111010110000000",
42654 => "0111010110000000",
42655 => "0111010110000000",
42656 => "0111010110000000",
42657 => "0111010110000000",
42658 => "0111010110000000",
42659 => "0111010110000000",
42660 => "0111010110000000",
42661 => "0111010110000000",
42662 => "0111010110000000",
42663 => "0111010110000000",
42664 => "0111010110000000",
42665 => "0111010110000000",
42666 => "0111010110000000",
42667 => "0111010110000000",
42668 => "0111010110000000",
42669 => "0111010110000000",
42670 => "0111010110000000",
42671 => "0111010110000000",
42672 => "0111010110000000",
42673 => "0111010110010000",
42674 => "0111010110010000",
42675 => "0111010110010000",
42676 => "0111010110010000",
42677 => "0111010110010000",
42678 => "0111010110010000",
42679 => "0111010110010000",
42680 => "0111010110010000",
42681 => "0111010110010000",
42682 => "0111010110010000",
42683 => "0111010110010000",
42684 => "0111010110010000",
42685 => "0111010110010000",
42686 => "0111010110010000",
42687 => "0111010110010000",
42688 => "0111010110010000",
42689 => "0111010110010000",
42690 => "0111010110010000",
42691 => "0111010110010000",
42692 => "0111010110010000",
42693 => "0111010110010000",
42694 => "0111010110010000",
42695 => "0111010110010000",
42696 => "0111010110010000",
42697 => "0111010110010000",
42698 => "0111010110010000",
42699 => "0111010110010000",
42700 => "0111010110100000",
42701 => "0111010110100000",
42702 => "0111010110100000",
42703 => "0111010110100000",
42704 => "0111010110100000",
42705 => "0111010110100000",
42706 => "0111010110100000",
42707 => "0111010110100000",
42708 => "0111010110100000",
42709 => "0111010110100000",
42710 => "0111010110100000",
42711 => "0111010110100000",
42712 => "0111010110100000",
42713 => "0111010110100000",
42714 => "0111010110100000",
42715 => "0111010110100000",
42716 => "0111010110100000",
42717 => "0111010110100000",
42718 => "0111010110100000",
42719 => "0111010110100000",
42720 => "0111010110100000",
42721 => "0111010110100000",
42722 => "0111010110100000",
42723 => "0111010110100000",
42724 => "0111010110100000",
42725 => "0111010110100000",
42726 => "0111010110100000",
42727 => "0111010110110000",
42728 => "0111010110110000",
42729 => "0111010110110000",
42730 => "0111010110110000",
42731 => "0111010110110000",
42732 => "0111010110110000",
42733 => "0111010110110000",
42734 => "0111010110110000",
42735 => "0111010110110000",
42736 => "0111010110110000",
42737 => "0111010110110000",
42738 => "0111010110110000",
42739 => "0111010110110000",
42740 => "0111010110110000",
42741 => "0111010110110000",
42742 => "0111010110110000",
42743 => "0111010110110000",
42744 => "0111010110110000",
42745 => "0111010110110000",
42746 => "0111010110110000",
42747 => "0111010110110000",
42748 => "0111010110110000",
42749 => "0111010110110000",
42750 => "0111010110110000",
42751 => "0111010110110000",
42752 => "0111010110110000",
42753 => "0111010110110000",
42754 => "0111010111000000",
42755 => "0111010111000000",
42756 => "0111010111000000",
42757 => "0111010111000000",
42758 => "0111010111000000",
42759 => "0111010111000000",
42760 => "0111010111000000",
42761 => "0111010111000000",
42762 => "0111010111000000",
42763 => "0111010111000000",
42764 => "0111010111000000",
42765 => "0111010111000000",
42766 => "0111010111000000",
42767 => "0111010111000000",
42768 => "0111010111000000",
42769 => "0111010111000000",
42770 => "0111010111000000",
42771 => "0111010111000000",
42772 => "0111010111000000",
42773 => "0111010111000000",
42774 => "0111010111000000",
42775 => "0111010111000000",
42776 => "0111010111000000",
42777 => "0111010111000000",
42778 => "0111010111000000",
42779 => "0111010111000000",
42780 => "0111010111000000",
42781 => "0111010111010000",
42782 => "0111010111010000",
42783 => "0111010111010000",
42784 => "0111010111010000",
42785 => "0111010111010000",
42786 => "0111010111010000",
42787 => "0111010111010000",
42788 => "0111010111010000",
42789 => "0111010111010000",
42790 => "0111010111010000",
42791 => "0111010111010000",
42792 => "0111010111010000",
42793 => "0111010111010000",
42794 => "0111010111010000",
42795 => "0111010111010000",
42796 => "0111010111010000",
42797 => "0111010111010000",
42798 => "0111010111010000",
42799 => "0111010111010000",
42800 => "0111010111010000",
42801 => "0111010111010000",
42802 => "0111010111010000",
42803 => "0111010111010000",
42804 => "0111010111010000",
42805 => "0111010111010000",
42806 => "0111010111010000",
42807 => "0111010111010000",
42808 => "0111010111100000",
42809 => "0111010111100000",
42810 => "0111010111100000",
42811 => "0111010111100000",
42812 => "0111010111100000",
42813 => "0111010111100000",
42814 => "0111010111100000",
42815 => "0111010111100000",
42816 => "0111010111100000",
42817 => "0111010111100000",
42818 => "0111010111100000",
42819 => "0111010111100000",
42820 => "0111010111100000",
42821 => "0111010111100000",
42822 => "0111010111100000",
42823 => "0111010111100000",
42824 => "0111010111100000",
42825 => "0111010111100000",
42826 => "0111010111100000",
42827 => "0111010111100000",
42828 => "0111010111100000",
42829 => "0111010111100000",
42830 => "0111010111100000",
42831 => "0111010111100000",
42832 => "0111010111100000",
42833 => "0111010111100000",
42834 => "0111010111100000",
42835 => "0111010111100000",
42836 => "0111010111110000",
42837 => "0111010111110000",
42838 => "0111010111110000",
42839 => "0111010111110000",
42840 => "0111010111110000",
42841 => "0111010111110000",
42842 => "0111010111110000",
42843 => "0111010111110000",
42844 => "0111010111110000",
42845 => "0111010111110000",
42846 => "0111010111110000",
42847 => "0111010111110000",
42848 => "0111010111110000",
42849 => "0111010111110000",
42850 => "0111010111110000",
42851 => "0111010111110000",
42852 => "0111010111110000",
42853 => "0111010111110000",
42854 => "0111010111110000",
42855 => "0111010111110000",
42856 => "0111010111110000",
42857 => "0111010111110000",
42858 => "0111010111110000",
42859 => "0111010111110000",
42860 => "0111010111110000",
42861 => "0111010111110000",
42862 => "0111010111110000",
42863 => "0111011000000000",
42864 => "0111011000000000",
42865 => "0111011000000000",
42866 => "0111011000000000",
42867 => "0111011000000000",
42868 => "0111011000000000",
42869 => "0111011000000000",
42870 => "0111011000000000",
42871 => "0111011000000000",
42872 => "0111011000000000",
42873 => "0111011000000000",
42874 => "0111011000000000",
42875 => "0111011000000000",
42876 => "0111011000000000",
42877 => "0111011000000000",
42878 => "0111011000000000",
42879 => "0111011000000000",
42880 => "0111011000000000",
42881 => "0111011000000000",
42882 => "0111011000000000",
42883 => "0111011000000000",
42884 => "0111011000000000",
42885 => "0111011000000000",
42886 => "0111011000000000",
42887 => "0111011000000000",
42888 => "0111011000000000",
42889 => "0111011000000000",
42890 => "0111011000000000",
42891 => "0111011000010000",
42892 => "0111011000010000",
42893 => "0111011000010000",
42894 => "0111011000010000",
42895 => "0111011000010000",
42896 => "0111011000010000",
42897 => "0111011000010000",
42898 => "0111011000010000",
42899 => "0111011000010000",
42900 => "0111011000010000",
42901 => "0111011000010000",
42902 => "0111011000010000",
42903 => "0111011000010000",
42904 => "0111011000010000",
42905 => "0111011000010000",
42906 => "0111011000010000",
42907 => "0111011000010000",
42908 => "0111011000010000",
42909 => "0111011000010000",
42910 => "0111011000010000",
42911 => "0111011000010000",
42912 => "0111011000010000",
42913 => "0111011000010000",
42914 => "0111011000010000",
42915 => "0111011000010000",
42916 => "0111011000010000",
42917 => "0111011000010000",
42918 => "0111011000010000",
42919 => "0111011000100000",
42920 => "0111011000100000",
42921 => "0111011000100000",
42922 => "0111011000100000",
42923 => "0111011000100000",
42924 => "0111011000100000",
42925 => "0111011000100000",
42926 => "0111011000100000",
42927 => "0111011000100000",
42928 => "0111011000100000",
42929 => "0111011000100000",
42930 => "0111011000100000",
42931 => "0111011000100000",
42932 => "0111011000100000",
42933 => "0111011000100000",
42934 => "0111011000100000",
42935 => "0111011000100000",
42936 => "0111011000100000",
42937 => "0111011000100000",
42938 => "0111011000100000",
42939 => "0111011000100000",
42940 => "0111011000100000",
42941 => "0111011000100000",
42942 => "0111011000100000",
42943 => "0111011000100000",
42944 => "0111011000100000",
42945 => "0111011000100000",
42946 => "0111011000100000",
42947 => "0111011000110000",
42948 => "0111011000110000",
42949 => "0111011000110000",
42950 => "0111011000110000",
42951 => "0111011000110000",
42952 => "0111011000110000",
42953 => "0111011000110000",
42954 => "0111011000110000",
42955 => "0111011000110000",
42956 => "0111011000110000",
42957 => "0111011000110000",
42958 => "0111011000110000",
42959 => "0111011000110000",
42960 => "0111011000110000",
42961 => "0111011000110000",
42962 => "0111011000110000",
42963 => "0111011000110000",
42964 => "0111011000110000",
42965 => "0111011000110000",
42966 => "0111011000110000",
42967 => "0111011000110000",
42968 => "0111011000110000",
42969 => "0111011000110000",
42970 => "0111011000110000",
42971 => "0111011000110000",
42972 => "0111011000110000",
42973 => "0111011000110000",
42974 => "0111011000110000",
42975 => "0111011001000000",
42976 => "0111011001000000",
42977 => "0111011001000000",
42978 => "0111011001000000",
42979 => "0111011001000000",
42980 => "0111011001000000",
42981 => "0111011001000000",
42982 => "0111011001000000",
42983 => "0111011001000000",
42984 => "0111011001000000",
42985 => "0111011001000000",
42986 => "0111011001000000",
42987 => "0111011001000000",
42988 => "0111011001000000",
42989 => "0111011001000000",
42990 => "0111011001000000",
42991 => "0111011001000000",
42992 => "0111011001000000",
42993 => "0111011001000000",
42994 => "0111011001000000",
42995 => "0111011001000000",
42996 => "0111011001000000",
42997 => "0111011001000000",
42998 => "0111011001000000",
42999 => "0111011001000000",
43000 => "0111011001000000",
43001 => "0111011001000000",
43002 => "0111011001000000",
43003 => "0111011001000000",
43004 => "0111011001010000",
43005 => "0111011001010000",
43006 => "0111011001010000",
43007 => "0111011001010000",
43008 => "0111011001010000",
43009 => "0111011001010000",
43010 => "0111011001010000",
43011 => "0111011001010000",
43012 => "0111011001010000",
43013 => "0111011001010000",
43014 => "0111011001010000",
43015 => "0111011001010000",
43016 => "0111011001010000",
43017 => "0111011001010000",
43018 => "0111011001010000",
43019 => "0111011001010000",
43020 => "0111011001010000",
43021 => "0111011001010000",
43022 => "0111011001010000",
43023 => "0111011001010000",
43024 => "0111011001010000",
43025 => "0111011001010000",
43026 => "0111011001010000",
43027 => "0111011001010000",
43028 => "0111011001010000",
43029 => "0111011001010000",
43030 => "0111011001010000",
43031 => "0111011001010000",
43032 => "0111011001100000",
43033 => "0111011001100000",
43034 => "0111011001100000",
43035 => "0111011001100000",
43036 => "0111011001100000",
43037 => "0111011001100000",
43038 => "0111011001100000",
43039 => "0111011001100000",
43040 => "0111011001100000",
43041 => "0111011001100000",
43042 => "0111011001100000",
43043 => "0111011001100000",
43044 => "0111011001100000",
43045 => "0111011001100000",
43046 => "0111011001100000",
43047 => "0111011001100000",
43048 => "0111011001100000",
43049 => "0111011001100000",
43050 => "0111011001100000",
43051 => "0111011001100000",
43052 => "0111011001100000",
43053 => "0111011001100000",
43054 => "0111011001100000",
43055 => "0111011001100000",
43056 => "0111011001100000",
43057 => "0111011001100000",
43058 => "0111011001100000",
43059 => "0111011001100000",
43060 => "0111011001100000",
43061 => "0111011001110000",
43062 => "0111011001110000",
43063 => "0111011001110000",
43064 => "0111011001110000",
43065 => "0111011001110000",
43066 => "0111011001110000",
43067 => "0111011001110000",
43068 => "0111011001110000",
43069 => "0111011001110000",
43070 => "0111011001110000",
43071 => "0111011001110000",
43072 => "0111011001110000",
43073 => "0111011001110000",
43074 => "0111011001110000",
43075 => "0111011001110000",
43076 => "0111011001110000",
43077 => "0111011001110000",
43078 => "0111011001110000",
43079 => "0111011001110000",
43080 => "0111011001110000",
43081 => "0111011001110000",
43082 => "0111011001110000",
43083 => "0111011001110000",
43084 => "0111011001110000",
43085 => "0111011001110000",
43086 => "0111011001110000",
43087 => "0111011001110000",
43088 => "0111011001110000",
43089 => "0111011001110000",
43090 => "0111011010000000",
43091 => "0111011010000000",
43092 => "0111011010000000",
43093 => "0111011010000000",
43094 => "0111011010000000",
43095 => "0111011010000000",
43096 => "0111011010000000",
43097 => "0111011010000000",
43098 => "0111011010000000",
43099 => "0111011010000000",
43100 => "0111011010000000",
43101 => "0111011010000000",
43102 => "0111011010000000",
43103 => "0111011010000000",
43104 => "0111011010000000",
43105 => "0111011010000000",
43106 => "0111011010000000",
43107 => "0111011010000000",
43108 => "0111011010000000",
43109 => "0111011010000000",
43110 => "0111011010000000",
43111 => "0111011010000000",
43112 => "0111011010000000",
43113 => "0111011010000000",
43114 => "0111011010000000",
43115 => "0111011010000000",
43116 => "0111011010000000",
43117 => "0111011010000000",
43118 => "0111011010000000",
43119 => "0111011010010000",
43120 => "0111011010010000",
43121 => "0111011010010000",
43122 => "0111011010010000",
43123 => "0111011010010000",
43124 => "0111011010010000",
43125 => "0111011010010000",
43126 => "0111011010010000",
43127 => "0111011010010000",
43128 => "0111011010010000",
43129 => "0111011010010000",
43130 => "0111011010010000",
43131 => "0111011010010000",
43132 => "0111011010010000",
43133 => "0111011010010000",
43134 => "0111011010010000",
43135 => "0111011010010000",
43136 => "0111011010010000",
43137 => "0111011010010000",
43138 => "0111011010010000",
43139 => "0111011010010000",
43140 => "0111011010010000",
43141 => "0111011010010000",
43142 => "0111011010010000",
43143 => "0111011010010000",
43144 => "0111011010010000",
43145 => "0111011010010000",
43146 => "0111011010010000",
43147 => "0111011010010000",
43148 => "0111011010100000",
43149 => "0111011010100000",
43150 => "0111011010100000",
43151 => "0111011010100000",
43152 => "0111011010100000",
43153 => "0111011010100000",
43154 => "0111011010100000",
43155 => "0111011010100000",
43156 => "0111011010100000",
43157 => "0111011010100000",
43158 => "0111011010100000",
43159 => "0111011010100000",
43160 => "0111011010100000",
43161 => "0111011010100000",
43162 => "0111011010100000",
43163 => "0111011010100000",
43164 => "0111011010100000",
43165 => "0111011010100000",
43166 => "0111011010100000",
43167 => "0111011010100000",
43168 => "0111011010100000",
43169 => "0111011010100000",
43170 => "0111011010100000",
43171 => "0111011010100000",
43172 => "0111011010100000",
43173 => "0111011010100000",
43174 => "0111011010100000",
43175 => "0111011010100000",
43176 => "0111011010100000",
43177 => "0111011010100000",
43178 => "0111011010110000",
43179 => "0111011010110000",
43180 => "0111011010110000",
43181 => "0111011010110000",
43182 => "0111011010110000",
43183 => "0111011010110000",
43184 => "0111011010110000",
43185 => "0111011010110000",
43186 => "0111011010110000",
43187 => "0111011010110000",
43188 => "0111011010110000",
43189 => "0111011010110000",
43190 => "0111011010110000",
43191 => "0111011010110000",
43192 => "0111011010110000",
43193 => "0111011010110000",
43194 => "0111011010110000",
43195 => "0111011010110000",
43196 => "0111011010110000",
43197 => "0111011010110000",
43198 => "0111011010110000",
43199 => "0111011010110000",
43200 => "0111011010110000",
43201 => "0111011010110000",
43202 => "0111011010110000",
43203 => "0111011010110000",
43204 => "0111011010110000",
43205 => "0111011010110000",
43206 => "0111011010110000",
43207 => "0111011010110000",
43208 => "0111011011000000",
43209 => "0111011011000000",
43210 => "0111011011000000",
43211 => "0111011011000000",
43212 => "0111011011000000",
43213 => "0111011011000000",
43214 => "0111011011000000",
43215 => "0111011011000000",
43216 => "0111011011000000",
43217 => "0111011011000000",
43218 => "0111011011000000",
43219 => "0111011011000000",
43220 => "0111011011000000",
43221 => "0111011011000000",
43222 => "0111011011000000",
43223 => "0111011011000000",
43224 => "0111011011000000",
43225 => "0111011011000000",
43226 => "0111011011000000",
43227 => "0111011011000000",
43228 => "0111011011000000",
43229 => "0111011011000000",
43230 => "0111011011000000",
43231 => "0111011011000000",
43232 => "0111011011000000",
43233 => "0111011011000000",
43234 => "0111011011000000",
43235 => "0111011011000000",
43236 => "0111011011000000",
43237 => "0111011011010000",
43238 => "0111011011010000",
43239 => "0111011011010000",
43240 => "0111011011010000",
43241 => "0111011011010000",
43242 => "0111011011010000",
43243 => "0111011011010000",
43244 => "0111011011010000",
43245 => "0111011011010000",
43246 => "0111011011010000",
43247 => "0111011011010000",
43248 => "0111011011010000",
43249 => "0111011011010000",
43250 => "0111011011010000",
43251 => "0111011011010000",
43252 => "0111011011010000",
43253 => "0111011011010000",
43254 => "0111011011010000",
43255 => "0111011011010000",
43256 => "0111011011010000",
43257 => "0111011011010000",
43258 => "0111011011010000",
43259 => "0111011011010000",
43260 => "0111011011010000",
43261 => "0111011011010000",
43262 => "0111011011010000",
43263 => "0111011011010000",
43264 => "0111011011010000",
43265 => "0111011011010000",
43266 => "0111011011010000",
43267 => "0111011011100000",
43268 => "0111011011100000",
43269 => "0111011011100000",
43270 => "0111011011100000",
43271 => "0111011011100000",
43272 => "0111011011100000",
43273 => "0111011011100000",
43274 => "0111011011100000",
43275 => "0111011011100000",
43276 => "0111011011100000",
43277 => "0111011011100000",
43278 => "0111011011100000",
43279 => "0111011011100000",
43280 => "0111011011100000",
43281 => "0111011011100000",
43282 => "0111011011100000",
43283 => "0111011011100000",
43284 => "0111011011100000",
43285 => "0111011011100000",
43286 => "0111011011100000",
43287 => "0111011011100000",
43288 => "0111011011100000",
43289 => "0111011011100000",
43290 => "0111011011100000",
43291 => "0111011011100000",
43292 => "0111011011100000",
43293 => "0111011011100000",
43294 => "0111011011100000",
43295 => "0111011011100000",
43296 => "0111011011100000",
43297 => "0111011011100000",
43298 => "0111011011110000",
43299 => "0111011011110000",
43300 => "0111011011110000",
43301 => "0111011011110000",
43302 => "0111011011110000",
43303 => "0111011011110000",
43304 => "0111011011110000",
43305 => "0111011011110000",
43306 => "0111011011110000",
43307 => "0111011011110000",
43308 => "0111011011110000",
43309 => "0111011011110000",
43310 => "0111011011110000",
43311 => "0111011011110000",
43312 => "0111011011110000",
43313 => "0111011011110000",
43314 => "0111011011110000",
43315 => "0111011011110000",
43316 => "0111011011110000",
43317 => "0111011011110000",
43318 => "0111011011110000",
43319 => "0111011011110000",
43320 => "0111011011110000",
43321 => "0111011011110000",
43322 => "0111011011110000",
43323 => "0111011011110000",
43324 => "0111011011110000",
43325 => "0111011011110000",
43326 => "0111011011110000",
43327 => "0111011011110000",
43328 => "0111011100000000",
43329 => "0111011100000000",
43330 => "0111011100000000",
43331 => "0111011100000000",
43332 => "0111011100000000",
43333 => "0111011100000000",
43334 => "0111011100000000",
43335 => "0111011100000000",
43336 => "0111011100000000",
43337 => "0111011100000000",
43338 => "0111011100000000",
43339 => "0111011100000000",
43340 => "0111011100000000",
43341 => "0111011100000000",
43342 => "0111011100000000",
43343 => "0111011100000000",
43344 => "0111011100000000",
43345 => "0111011100000000",
43346 => "0111011100000000",
43347 => "0111011100000000",
43348 => "0111011100000000",
43349 => "0111011100000000",
43350 => "0111011100000000",
43351 => "0111011100000000",
43352 => "0111011100000000",
43353 => "0111011100000000",
43354 => "0111011100000000",
43355 => "0111011100000000",
43356 => "0111011100000000",
43357 => "0111011100000000",
43358 => "0111011100000000",
43359 => "0111011100010000",
43360 => "0111011100010000",
43361 => "0111011100010000",
43362 => "0111011100010000",
43363 => "0111011100010000",
43364 => "0111011100010000",
43365 => "0111011100010000",
43366 => "0111011100010000",
43367 => "0111011100010000",
43368 => "0111011100010000",
43369 => "0111011100010000",
43370 => "0111011100010000",
43371 => "0111011100010000",
43372 => "0111011100010000",
43373 => "0111011100010000",
43374 => "0111011100010000",
43375 => "0111011100010000",
43376 => "0111011100010000",
43377 => "0111011100010000",
43378 => "0111011100010000",
43379 => "0111011100010000",
43380 => "0111011100010000",
43381 => "0111011100010000",
43382 => "0111011100010000",
43383 => "0111011100010000",
43384 => "0111011100010000",
43385 => "0111011100010000",
43386 => "0111011100010000",
43387 => "0111011100010000",
43388 => "0111011100010000",
43389 => "0111011100100000",
43390 => "0111011100100000",
43391 => "0111011100100000",
43392 => "0111011100100000",
43393 => "0111011100100000",
43394 => "0111011100100000",
43395 => "0111011100100000",
43396 => "0111011100100000",
43397 => "0111011100100000",
43398 => "0111011100100000",
43399 => "0111011100100000",
43400 => "0111011100100000",
43401 => "0111011100100000",
43402 => "0111011100100000",
43403 => "0111011100100000",
43404 => "0111011100100000",
43405 => "0111011100100000",
43406 => "0111011100100000",
43407 => "0111011100100000",
43408 => "0111011100100000",
43409 => "0111011100100000",
43410 => "0111011100100000",
43411 => "0111011100100000",
43412 => "0111011100100000",
43413 => "0111011100100000",
43414 => "0111011100100000",
43415 => "0111011100100000",
43416 => "0111011100100000",
43417 => "0111011100100000",
43418 => "0111011100100000",
43419 => "0111011100100000",
43420 => "0111011100110000",
43421 => "0111011100110000",
43422 => "0111011100110000",
43423 => "0111011100110000",
43424 => "0111011100110000",
43425 => "0111011100110000",
43426 => "0111011100110000",
43427 => "0111011100110000",
43428 => "0111011100110000",
43429 => "0111011100110000",
43430 => "0111011100110000",
43431 => "0111011100110000",
43432 => "0111011100110000",
43433 => "0111011100110000",
43434 => "0111011100110000",
43435 => "0111011100110000",
43436 => "0111011100110000",
43437 => "0111011100110000",
43438 => "0111011100110000",
43439 => "0111011100110000",
43440 => "0111011100110000",
43441 => "0111011100110000",
43442 => "0111011100110000",
43443 => "0111011100110000",
43444 => "0111011100110000",
43445 => "0111011100110000",
43446 => "0111011100110000",
43447 => "0111011100110000",
43448 => "0111011100110000",
43449 => "0111011100110000",
43450 => "0111011100110000",
43451 => "0111011100110000",
43452 => "0111011101000000",
43453 => "0111011101000000",
43454 => "0111011101000000",
43455 => "0111011101000000",
43456 => "0111011101000000",
43457 => "0111011101000000",
43458 => "0111011101000000",
43459 => "0111011101000000",
43460 => "0111011101000000",
43461 => "0111011101000000",
43462 => "0111011101000000",
43463 => "0111011101000000",
43464 => "0111011101000000",
43465 => "0111011101000000",
43466 => "0111011101000000",
43467 => "0111011101000000",
43468 => "0111011101000000",
43469 => "0111011101000000",
43470 => "0111011101000000",
43471 => "0111011101000000",
43472 => "0111011101000000",
43473 => "0111011101000000",
43474 => "0111011101000000",
43475 => "0111011101000000",
43476 => "0111011101000000",
43477 => "0111011101000000",
43478 => "0111011101000000",
43479 => "0111011101000000",
43480 => "0111011101000000",
43481 => "0111011101000000",
43482 => "0111011101000000",
43483 => "0111011101010000",
43484 => "0111011101010000",
43485 => "0111011101010000",
43486 => "0111011101010000",
43487 => "0111011101010000",
43488 => "0111011101010000",
43489 => "0111011101010000",
43490 => "0111011101010000",
43491 => "0111011101010000",
43492 => "0111011101010000",
43493 => "0111011101010000",
43494 => "0111011101010000",
43495 => "0111011101010000",
43496 => "0111011101010000",
43497 => "0111011101010000",
43498 => "0111011101010000",
43499 => "0111011101010000",
43500 => "0111011101010000",
43501 => "0111011101010000",
43502 => "0111011101010000",
43503 => "0111011101010000",
43504 => "0111011101010000",
43505 => "0111011101010000",
43506 => "0111011101010000",
43507 => "0111011101010000",
43508 => "0111011101010000",
43509 => "0111011101010000",
43510 => "0111011101010000",
43511 => "0111011101010000",
43512 => "0111011101010000",
43513 => "0111011101010000",
43514 => "0111011101010000",
43515 => "0111011101100000",
43516 => "0111011101100000",
43517 => "0111011101100000",
43518 => "0111011101100000",
43519 => "0111011101100000",
43520 => "0111011101100000",
43521 => "0111011101100000",
43522 => "0111011101100000",
43523 => "0111011101100000",
43524 => "0111011101100000",
43525 => "0111011101100000",
43526 => "0111011101100000",
43527 => "0111011101100000",
43528 => "0111011101100000",
43529 => "0111011101100000",
43530 => "0111011101100000",
43531 => "0111011101100000",
43532 => "0111011101100000",
43533 => "0111011101100000",
43534 => "0111011101100000",
43535 => "0111011101100000",
43536 => "0111011101100000",
43537 => "0111011101100000",
43538 => "0111011101100000",
43539 => "0111011101100000",
43540 => "0111011101100000",
43541 => "0111011101100000",
43542 => "0111011101100000",
43543 => "0111011101100000",
43544 => "0111011101100000",
43545 => "0111011101100000",
43546 => "0111011101110000",
43547 => "0111011101110000",
43548 => "0111011101110000",
43549 => "0111011101110000",
43550 => "0111011101110000",
43551 => "0111011101110000",
43552 => "0111011101110000",
43553 => "0111011101110000",
43554 => "0111011101110000",
43555 => "0111011101110000",
43556 => "0111011101110000",
43557 => "0111011101110000",
43558 => "0111011101110000",
43559 => "0111011101110000",
43560 => "0111011101110000",
43561 => "0111011101110000",
43562 => "0111011101110000",
43563 => "0111011101110000",
43564 => "0111011101110000",
43565 => "0111011101110000",
43566 => "0111011101110000",
43567 => "0111011101110000",
43568 => "0111011101110000",
43569 => "0111011101110000",
43570 => "0111011101110000",
43571 => "0111011101110000",
43572 => "0111011101110000",
43573 => "0111011101110000",
43574 => "0111011101110000",
43575 => "0111011101110000",
43576 => "0111011101110000",
43577 => "0111011101110000",
43578 => "0111011110000000",
43579 => "0111011110000000",
43580 => "0111011110000000",
43581 => "0111011110000000",
43582 => "0111011110000000",
43583 => "0111011110000000",
43584 => "0111011110000000",
43585 => "0111011110000000",
43586 => "0111011110000000",
43587 => "0111011110000000",
43588 => "0111011110000000",
43589 => "0111011110000000",
43590 => "0111011110000000",
43591 => "0111011110000000",
43592 => "0111011110000000",
43593 => "0111011110000000",
43594 => "0111011110000000",
43595 => "0111011110000000",
43596 => "0111011110000000",
43597 => "0111011110000000",
43598 => "0111011110000000",
43599 => "0111011110000000",
43600 => "0111011110000000",
43601 => "0111011110000000",
43602 => "0111011110000000",
43603 => "0111011110000000",
43604 => "0111011110000000",
43605 => "0111011110000000",
43606 => "0111011110000000",
43607 => "0111011110000000",
43608 => "0111011110000000",
43609 => "0111011110000000",
43610 => "0111011110000000",
43611 => "0111011110010000",
43612 => "0111011110010000",
43613 => "0111011110010000",
43614 => "0111011110010000",
43615 => "0111011110010000",
43616 => "0111011110010000",
43617 => "0111011110010000",
43618 => "0111011110010000",
43619 => "0111011110010000",
43620 => "0111011110010000",
43621 => "0111011110010000",
43622 => "0111011110010000",
43623 => "0111011110010000",
43624 => "0111011110010000",
43625 => "0111011110010000",
43626 => "0111011110010000",
43627 => "0111011110010000",
43628 => "0111011110010000",
43629 => "0111011110010000",
43630 => "0111011110010000",
43631 => "0111011110010000",
43632 => "0111011110010000",
43633 => "0111011110010000",
43634 => "0111011110010000",
43635 => "0111011110010000",
43636 => "0111011110010000",
43637 => "0111011110010000",
43638 => "0111011110010000",
43639 => "0111011110010000",
43640 => "0111011110010000",
43641 => "0111011110010000",
43642 => "0111011110010000",
43643 => "0111011110100000",
43644 => "0111011110100000",
43645 => "0111011110100000",
43646 => "0111011110100000",
43647 => "0111011110100000",
43648 => "0111011110100000",
43649 => "0111011110100000",
43650 => "0111011110100000",
43651 => "0111011110100000",
43652 => "0111011110100000",
43653 => "0111011110100000",
43654 => "0111011110100000",
43655 => "0111011110100000",
43656 => "0111011110100000",
43657 => "0111011110100000",
43658 => "0111011110100000",
43659 => "0111011110100000",
43660 => "0111011110100000",
43661 => "0111011110100000",
43662 => "0111011110100000",
43663 => "0111011110100000",
43664 => "0111011110100000",
43665 => "0111011110100000",
43666 => "0111011110100000",
43667 => "0111011110100000",
43668 => "0111011110100000",
43669 => "0111011110100000",
43670 => "0111011110100000",
43671 => "0111011110100000",
43672 => "0111011110100000",
43673 => "0111011110100000",
43674 => "0111011110100000",
43675 => "0111011110100000",
43676 => "0111011110110000",
43677 => "0111011110110000",
43678 => "0111011110110000",
43679 => "0111011110110000",
43680 => "0111011110110000",
43681 => "0111011110110000",
43682 => "0111011110110000",
43683 => "0111011110110000",
43684 => "0111011110110000",
43685 => "0111011110110000",
43686 => "0111011110110000",
43687 => "0111011110110000",
43688 => "0111011110110000",
43689 => "0111011110110000",
43690 => "0111011110110000",
43691 => "0111011110110000",
43692 => "0111011110110000",
43693 => "0111011110110000",
43694 => "0111011110110000",
43695 => "0111011110110000",
43696 => "0111011110110000",
43697 => "0111011110110000",
43698 => "0111011110110000",
43699 => "0111011110110000",
43700 => "0111011110110000",
43701 => "0111011110110000",
43702 => "0111011110110000",
43703 => "0111011110110000",
43704 => "0111011110110000",
43705 => "0111011110110000",
43706 => "0111011110110000",
43707 => "0111011110110000",
43708 => "0111011110110000",
43709 => "0111011111000000",
43710 => "0111011111000000",
43711 => "0111011111000000",
43712 => "0111011111000000",
43713 => "0111011111000000",
43714 => "0111011111000000",
43715 => "0111011111000000",
43716 => "0111011111000000",
43717 => "0111011111000000",
43718 => "0111011111000000",
43719 => "0111011111000000",
43720 => "0111011111000000",
43721 => "0111011111000000",
43722 => "0111011111000000",
43723 => "0111011111000000",
43724 => "0111011111000000",
43725 => "0111011111000000",
43726 => "0111011111000000",
43727 => "0111011111000000",
43728 => "0111011111000000",
43729 => "0111011111000000",
43730 => "0111011111000000",
43731 => "0111011111000000",
43732 => "0111011111000000",
43733 => "0111011111000000",
43734 => "0111011111000000",
43735 => "0111011111000000",
43736 => "0111011111000000",
43737 => "0111011111000000",
43738 => "0111011111000000",
43739 => "0111011111000000",
43740 => "0111011111000000",
43741 => "0111011111000000",
43742 => "0111011111010000",
43743 => "0111011111010000",
43744 => "0111011111010000",
43745 => "0111011111010000",
43746 => "0111011111010000",
43747 => "0111011111010000",
43748 => "0111011111010000",
43749 => "0111011111010000",
43750 => "0111011111010000",
43751 => "0111011111010000",
43752 => "0111011111010000",
43753 => "0111011111010000",
43754 => "0111011111010000",
43755 => "0111011111010000",
43756 => "0111011111010000",
43757 => "0111011111010000",
43758 => "0111011111010000",
43759 => "0111011111010000",
43760 => "0111011111010000",
43761 => "0111011111010000",
43762 => "0111011111010000",
43763 => "0111011111010000",
43764 => "0111011111010000",
43765 => "0111011111010000",
43766 => "0111011111010000",
43767 => "0111011111010000",
43768 => "0111011111010000",
43769 => "0111011111010000",
43770 => "0111011111010000",
43771 => "0111011111010000",
43772 => "0111011111010000",
43773 => "0111011111010000",
43774 => "0111011111010000",
43775 => "0111011111100000",
43776 => "0111011111100000",
43777 => "0111011111100000",
43778 => "0111011111100000",
43779 => "0111011111100000",
43780 => "0111011111100000",
43781 => "0111011111100000",
43782 => "0111011111100000",
43783 => "0111011111100000",
43784 => "0111011111100000",
43785 => "0111011111100000",
43786 => "0111011111100000",
43787 => "0111011111100000",
43788 => "0111011111100000",
43789 => "0111011111100000",
43790 => "0111011111100000",
43791 => "0111011111100000",
43792 => "0111011111100000",
43793 => "0111011111100000",
43794 => "0111011111100000",
43795 => "0111011111100000",
43796 => "0111011111100000",
43797 => "0111011111100000",
43798 => "0111011111100000",
43799 => "0111011111100000",
43800 => "0111011111100000",
43801 => "0111011111100000",
43802 => "0111011111100000",
43803 => "0111011111100000",
43804 => "0111011111100000",
43805 => "0111011111100000",
43806 => "0111011111100000",
43807 => "0111011111100000",
43808 => "0111011111100000",
43809 => "0111011111110000",
43810 => "0111011111110000",
43811 => "0111011111110000",
43812 => "0111011111110000",
43813 => "0111011111110000",
43814 => "0111011111110000",
43815 => "0111011111110000",
43816 => "0111011111110000",
43817 => "0111011111110000",
43818 => "0111011111110000",
43819 => "0111011111110000",
43820 => "0111011111110000",
43821 => "0111011111110000",
43822 => "0111011111110000",
43823 => "0111011111110000",
43824 => "0111011111110000",
43825 => "0111011111110000",
43826 => "0111011111110000",
43827 => "0111011111110000",
43828 => "0111011111110000",
43829 => "0111011111110000",
43830 => "0111011111110000",
43831 => "0111011111110000",
43832 => "0111011111110000",
43833 => "0111011111110000",
43834 => "0111011111110000",
43835 => "0111011111110000",
43836 => "0111011111110000",
43837 => "0111011111110000",
43838 => "0111011111110000",
43839 => "0111011111110000",
43840 => "0111011111110000",
43841 => "0111011111110000",
43842 => "0111011111110000",
43843 => "0111100000000000",
43844 => "0111100000000000",
43845 => "0111100000000000",
43846 => "0111100000000000",
43847 => "0111100000000000",
43848 => "0111100000000000",
43849 => "0111100000000000",
43850 => "0111100000000000",
43851 => "0111100000000000",
43852 => "0111100000000000",
43853 => "0111100000000000",
43854 => "0111100000000000",
43855 => "0111100000000000",
43856 => "0111100000000000",
43857 => "0111100000000000",
43858 => "0111100000000000",
43859 => "0111100000000000",
43860 => "0111100000000000",
43861 => "0111100000000000",
43862 => "0111100000000000",
43863 => "0111100000000000",
43864 => "0111100000000000",
43865 => "0111100000000000",
43866 => "0111100000000000",
43867 => "0111100000000000",
43868 => "0111100000000000",
43869 => "0111100000000000",
43870 => "0111100000000000",
43871 => "0111100000000000",
43872 => "0111100000000000",
43873 => "0111100000000000",
43874 => "0111100000000000",
43875 => "0111100000000000",
43876 => "0111100000000000",
43877 => "0111100000010000",
43878 => "0111100000010000",
43879 => "0111100000010000",
43880 => "0111100000010000",
43881 => "0111100000010000",
43882 => "0111100000010000",
43883 => "0111100000010000",
43884 => "0111100000010000",
43885 => "0111100000010000",
43886 => "0111100000010000",
43887 => "0111100000010000",
43888 => "0111100000010000",
43889 => "0111100000010000",
43890 => "0111100000010000",
43891 => "0111100000010000",
43892 => "0111100000010000",
43893 => "0111100000010000",
43894 => "0111100000010000",
43895 => "0111100000010000",
43896 => "0111100000010000",
43897 => "0111100000010000",
43898 => "0111100000010000",
43899 => "0111100000010000",
43900 => "0111100000010000",
43901 => "0111100000010000",
43902 => "0111100000010000",
43903 => "0111100000010000",
43904 => "0111100000010000",
43905 => "0111100000010000",
43906 => "0111100000010000",
43907 => "0111100000010000",
43908 => "0111100000010000",
43909 => "0111100000010000",
43910 => "0111100000010000",
43911 => "0111100000100000",
43912 => "0111100000100000",
43913 => "0111100000100000",
43914 => "0111100000100000",
43915 => "0111100000100000",
43916 => "0111100000100000",
43917 => "0111100000100000",
43918 => "0111100000100000",
43919 => "0111100000100000",
43920 => "0111100000100000",
43921 => "0111100000100000",
43922 => "0111100000100000",
43923 => "0111100000100000",
43924 => "0111100000100000",
43925 => "0111100000100000",
43926 => "0111100000100000",
43927 => "0111100000100000",
43928 => "0111100000100000",
43929 => "0111100000100000",
43930 => "0111100000100000",
43931 => "0111100000100000",
43932 => "0111100000100000",
43933 => "0111100000100000",
43934 => "0111100000100000",
43935 => "0111100000100000",
43936 => "0111100000100000",
43937 => "0111100000100000",
43938 => "0111100000100000",
43939 => "0111100000100000",
43940 => "0111100000100000",
43941 => "0111100000100000",
43942 => "0111100000100000",
43943 => "0111100000100000",
43944 => "0111100000100000",
43945 => "0111100000100000",
43946 => "0111100000110000",
43947 => "0111100000110000",
43948 => "0111100000110000",
43949 => "0111100000110000",
43950 => "0111100000110000",
43951 => "0111100000110000",
43952 => "0111100000110000",
43953 => "0111100000110000",
43954 => "0111100000110000",
43955 => "0111100000110000",
43956 => "0111100000110000",
43957 => "0111100000110000",
43958 => "0111100000110000",
43959 => "0111100000110000",
43960 => "0111100000110000",
43961 => "0111100000110000",
43962 => "0111100000110000",
43963 => "0111100000110000",
43964 => "0111100000110000",
43965 => "0111100000110000",
43966 => "0111100000110000",
43967 => "0111100000110000",
43968 => "0111100000110000",
43969 => "0111100000110000",
43970 => "0111100000110000",
43971 => "0111100000110000",
43972 => "0111100000110000",
43973 => "0111100000110000",
43974 => "0111100000110000",
43975 => "0111100000110000",
43976 => "0111100000110000",
43977 => "0111100000110000",
43978 => "0111100000110000",
43979 => "0111100000110000",
43980 => "0111100000110000",
43981 => "0111100001000000",
43982 => "0111100001000000",
43983 => "0111100001000000",
43984 => "0111100001000000",
43985 => "0111100001000000",
43986 => "0111100001000000",
43987 => "0111100001000000",
43988 => "0111100001000000",
43989 => "0111100001000000",
43990 => "0111100001000000",
43991 => "0111100001000000",
43992 => "0111100001000000",
43993 => "0111100001000000",
43994 => "0111100001000000",
43995 => "0111100001000000",
43996 => "0111100001000000",
43997 => "0111100001000000",
43998 => "0111100001000000",
43999 => "0111100001000000",
44000 => "0111100001000000",
44001 => "0111100001000000",
44002 => "0111100001000000",
44003 => "0111100001000000",
44004 => "0111100001000000",
44005 => "0111100001000000",
44006 => "0111100001000000",
44007 => "0111100001000000",
44008 => "0111100001000000",
44009 => "0111100001000000",
44010 => "0111100001000000",
44011 => "0111100001000000",
44012 => "0111100001000000",
44013 => "0111100001000000",
44014 => "0111100001000000",
44015 => "0111100001000000",
44016 => "0111100001010000",
44017 => "0111100001010000",
44018 => "0111100001010000",
44019 => "0111100001010000",
44020 => "0111100001010000",
44021 => "0111100001010000",
44022 => "0111100001010000",
44023 => "0111100001010000",
44024 => "0111100001010000",
44025 => "0111100001010000",
44026 => "0111100001010000",
44027 => "0111100001010000",
44028 => "0111100001010000",
44029 => "0111100001010000",
44030 => "0111100001010000",
44031 => "0111100001010000",
44032 => "0111100001010000",
44033 => "0111100001010000",
44034 => "0111100001010000",
44035 => "0111100001010000",
44036 => "0111100001010000",
44037 => "0111100001010000",
44038 => "0111100001010000",
44039 => "0111100001010000",
44040 => "0111100001010000",
44041 => "0111100001010000",
44042 => "0111100001010000",
44043 => "0111100001010000",
44044 => "0111100001010000",
44045 => "0111100001010000",
44046 => "0111100001010000",
44047 => "0111100001010000",
44048 => "0111100001010000",
44049 => "0111100001010000",
44050 => "0111100001010000",
44051 => "0111100001010000",
44052 => "0111100001100000",
44053 => "0111100001100000",
44054 => "0111100001100000",
44055 => "0111100001100000",
44056 => "0111100001100000",
44057 => "0111100001100000",
44058 => "0111100001100000",
44059 => "0111100001100000",
44060 => "0111100001100000",
44061 => "0111100001100000",
44062 => "0111100001100000",
44063 => "0111100001100000",
44064 => "0111100001100000",
44065 => "0111100001100000",
44066 => "0111100001100000",
44067 => "0111100001100000",
44068 => "0111100001100000",
44069 => "0111100001100000",
44070 => "0111100001100000",
44071 => "0111100001100000",
44072 => "0111100001100000",
44073 => "0111100001100000",
44074 => "0111100001100000",
44075 => "0111100001100000",
44076 => "0111100001100000",
44077 => "0111100001100000",
44078 => "0111100001100000",
44079 => "0111100001100000",
44080 => "0111100001100000",
44081 => "0111100001100000",
44082 => "0111100001100000",
44083 => "0111100001100000",
44084 => "0111100001100000",
44085 => "0111100001100000",
44086 => "0111100001100000",
44087 => "0111100001110000",
44088 => "0111100001110000",
44089 => "0111100001110000",
44090 => "0111100001110000",
44091 => "0111100001110000",
44092 => "0111100001110000",
44093 => "0111100001110000",
44094 => "0111100001110000",
44095 => "0111100001110000",
44096 => "0111100001110000",
44097 => "0111100001110000",
44098 => "0111100001110000",
44099 => "0111100001110000",
44100 => "0111100001110000",
44101 => "0111100001110000",
44102 => "0111100001110000",
44103 => "0111100001110000",
44104 => "0111100001110000",
44105 => "0111100001110000",
44106 => "0111100001110000",
44107 => "0111100001110000",
44108 => "0111100001110000",
44109 => "0111100001110000",
44110 => "0111100001110000",
44111 => "0111100001110000",
44112 => "0111100001110000",
44113 => "0111100001110000",
44114 => "0111100001110000",
44115 => "0111100001110000",
44116 => "0111100001110000",
44117 => "0111100001110000",
44118 => "0111100001110000",
44119 => "0111100001110000",
44120 => "0111100001110000",
44121 => "0111100001110000",
44122 => "0111100001110000",
44123 => "0111100010000000",
44124 => "0111100010000000",
44125 => "0111100010000000",
44126 => "0111100010000000",
44127 => "0111100010000000",
44128 => "0111100010000000",
44129 => "0111100010000000",
44130 => "0111100010000000",
44131 => "0111100010000000",
44132 => "0111100010000000",
44133 => "0111100010000000",
44134 => "0111100010000000",
44135 => "0111100010000000",
44136 => "0111100010000000",
44137 => "0111100010000000",
44138 => "0111100010000000",
44139 => "0111100010000000",
44140 => "0111100010000000",
44141 => "0111100010000000",
44142 => "0111100010000000",
44143 => "0111100010000000",
44144 => "0111100010000000",
44145 => "0111100010000000",
44146 => "0111100010000000",
44147 => "0111100010000000",
44148 => "0111100010000000",
44149 => "0111100010000000",
44150 => "0111100010000000",
44151 => "0111100010000000",
44152 => "0111100010000000",
44153 => "0111100010000000",
44154 => "0111100010000000",
44155 => "0111100010000000",
44156 => "0111100010000000",
44157 => "0111100010000000",
44158 => "0111100010000000",
44159 => "0111100010000000",
44160 => "0111100010010000",
44161 => "0111100010010000",
44162 => "0111100010010000",
44163 => "0111100010010000",
44164 => "0111100010010000",
44165 => "0111100010010000",
44166 => "0111100010010000",
44167 => "0111100010010000",
44168 => "0111100010010000",
44169 => "0111100010010000",
44170 => "0111100010010000",
44171 => "0111100010010000",
44172 => "0111100010010000",
44173 => "0111100010010000",
44174 => "0111100010010000",
44175 => "0111100010010000",
44176 => "0111100010010000",
44177 => "0111100010010000",
44178 => "0111100010010000",
44179 => "0111100010010000",
44180 => "0111100010010000",
44181 => "0111100010010000",
44182 => "0111100010010000",
44183 => "0111100010010000",
44184 => "0111100010010000",
44185 => "0111100010010000",
44186 => "0111100010010000",
44187 => "0111100010010000",
44188 => "0111100010010000",
44189 => "0111100010010000",
44190 => "0111100010010000",
44191 => "0111100010010000",
44192 => "0111100010010000",
44193 => "0111100010010000",
44194 => "0111100010010000",
44195 => "0111100010010000",
44196 => "0111100010100000",
44197 => "0111100010100000",
44198 => "0111100010100000",
44199 => "0111100010100000",
44200 => "0111100010100000",
44201 => "0111100010100000",
44202 => "0111100010100000",
44203 => "0111100010100000",
44204 => "0111100010100000",
44205 => "0111100010100000",
44206 => "0111100010100000",
44207 => "0111100010100000",
44208 => "0111100010100000",
44209 => "0111100010100000",
44210 => "0111100010100000",
44211 => "0111100010100000",
44212 => "0111100010100000",
44213 => "0111100010100000",
44214 => "0111100010100000",
44215 => "0111100010100000",
44216 => "0111100010100000",
44217 => "0111100010100000",
44218 => "0111100010100000",
44219 => "0111100010100000",
44220 => "0111100010100000",
44221 => "0111100010100000",
44222 => "0111100010100000",
44223 => "0111100010100000",
44224 => "0111100010100000",
44225 => "0111100010100000",
44226 => "0111100010100000",
44227 => "0111100010100000",
44228 => "0111100010100000",
44229 => "0111100010100000",
44230 => "0111100010100000",
44231 => "0111100010100000",
44232 => "0111100010100000",
44233 => "0111100010110000",
44234 => "0111100010110000",
44235 => "0111100010110000",
44236 => "0111100010110000",
44237 => "0111100010110000",
44238 => "0111100010110000",
44239 => "0111100010110000",
44240 => "0111100010110000",
44241 => "0111100010110000",
44242 => "0111100010110000",
44243 => "0111100010110000",
44244 => "0111100010110000",
44245 => "0111100010110000",
44246 => "0111100010110000",
44247 => "0111100010110000",
44248 => "0111100010110000",
44249 => "0111100010110000",
44250 => "0111100010110000",
44251 => "0111100010110000",
44252 => "0111100010110000",
44253 => "0111100010110000",
44254 => "0111100010110000",
44255 => "0111100010110000",
44256 => "0111100010110000",
44257 => "0111100010110000",
44258 => "0111100010110000",
44259 => "0111100010110000",
44260 => "0111100010110000",
44261 => "0111100010110000",
44262 => "0111100010110000",
44263 => "0111100010110000",
44264 => "0111100010110000",
44265 => "0111100010110000",
44266 => "0111100010110000",
44267 => "0111100010110000",
44268 => "0111100010110000",
44269 => "0111100010110000",
44270 => "0111100011000000",
44271 => "0111100011000000",
44272 => "0111100011000000",
44273 => "0111100011000000",
44274 => "0111100011000000",
44275 => "0111100011000000",
44276 => "0111100011000000",
44277 => "0111100011000000",
44278 => "0111100011000000",
44279 => "0111100011000000",
44280 => "0111100011000000",
44281 => "0111100011000000",
44282 => "0111100011000000",
44283 => "0111100011000000",
44284 => "0111100011000000",
44285 => "0111100011000000",
44286 => "0111100011000000",
44287 => "0111100011000000",
44288 => "0111100011000000",
44289 => "0111100011000000",
44290 => "0111100011000000",
44291 => "0111100011000000",
44292 => "0111100011000000",
44293 => "0111100011000000",
44294 => "0111100011000000",
44295 => "0111100011000000",
44296 => "0111100011000000",
44297 => "0111100011000000",
44298 => "0111100011000000",
44299 => "0111100011000000",
44300 => "0111100011000000",
44301 => "0111100011000000",
44302 => "0111100011000000",
44303 => "0111100011000000",
44304 => "0111100011000000",
44305 => "0111100011000000",
44306 => "0111100011000000",
44307 => "0111100011010000",
44308 => "0111100011010000",
44309 => "0111100011010000",
44310 => "0111100011010000",
44311 => "0111100011010000",
44312 => "0111100011010000",
44313 => "0111100011010000",
44314 => "0111100011010000",
44315 => "0111100011010000",
44316 => "0111100011010000",
44317 => "0111100011010000",
44318 => "0111100011010000",
44319 => "0111100011010000",
44320 => "0111100011010000",
44321 => "0111100011010000",
44322 => "0111100011010000",
44323 => "0111100011010000",
44324 => "0111100011010000",
44325 => "0111100011010000",
44326 => "0111100011010000",
44327 => "0111100011010000",
44328 => "0111100011010000",
44329 => "0111100011010000",
44330 => "0111100011010000",
44331 => "0111100011010000",
44332 => "0111100011010000",
44333 => "0111100011010000",
44334 => "0111100011010000",
44335 => "0111100011010000",
44336 => "0111100011010000",
44337 => "0111100011010000",
44338 => "0111100011010000",
44339 => "0111100011010000",
44340 => "0111100011010000",
44341 => "0111100011010000",
44342 => "0111100011010000",
44343 => "0111100011010000",
44344 => "0111100011010000",
44345 => "0111100011100000",
44346 => "0111100011100000",
44347 => "0111100011100000",
44348 => "0111100011100000",
44349 => "0111100011100000",
44350 => "0111100011100000",
44351 => "0111100011100000",
44352 => "0111100011100000",
44353 => "0111100011100000",
44354 => "0111100011100000",
44355 => "0111100011100000",
44356 => "0111100011100000",
44357 => "0111100011100000",
44358 => "0111100011100000",
44359 => "0111100011100000",
44360 => "0111100011100000",
44361 => "0111100011100000",
44362 => "0111100011100000",
44363 => "0111100011100000",
44364 => "0111100011100000",
44365 => "0111100011100000",
44366 => "0111100011100000",
44367 => "0111100011100000",
44368 => "0111100011100000",
44369 => "0111100011100000",
44370 => "0111100011100000",
44371 => "0111100011100000",
44372 => "0111100011100000",
44373 => "0111100011100000",
44374 => "0111100011100000",
44375 => "0111100011100000",
44376 => "0111100011100000",
44377 => "0111100011100000",
44378 => "0111100011100000",
44379 => "0111100011100000",
44380 => "0111100011100000",
44381 => "0111100011100000",
44382 => "0111100011100000",
44383 => "0111100011110000",
44384 => "0111100011110000",
44385 => "0111100011110000",
44386 => "0111100011110000",
44387 => "0111100011110000",
44388 => "0111100011110000",
44389 => "0111100011110000",
44390 => "0111100011110000",
44391 => "0111100011110000",
44392 => "0111100011110000",
44393 => "0111100011110000",
44394 => "0111100011110000",
44395 => "0111100011110000",
44396 => "0111100011110000",
44397 => "0111100011110000",
44398 => "0111100011110000",
44399 => "0111100011110000",
44400 => "0111100011110000",
44401 => "0111100011110000",
44402 => "0111100011110000",
44403 => "0111100011110000",
44404 => "0111100011110000",
44405 => "0111100011110000",
44406 => "0111100011110000",
44407 => "0111100011110000",
44408 => "0111100011110000",
44409 => "0111100011110000",
44410 => "0111100011110000",
44411 => "0111100011110000",
44412 => "0111100011110000",
44413 => "0111100011110000",
44414 => "0111100011110000",
44415 => "0111100011110000",
44416 => "0111100011110000",
44417 => "0111100011110000",
44418 => "0111100011110000",
44419 => "0111100011110000",
44420 => "0111100011110000",
44421 => "0111100011110000",
44422 => "0111100100000000",
44423 => "0111100100000000",
44424 => "0111100100000000",
44425 => "0111100100000000",
44426 => "0111100100000000",
44427 => "0111100100000000",
44428 => "0111100100000000",
44429 => "0111100100000000",
44430 => "0111100100000000",
44431 => "0111100100000000",
44432 => "0111100100000000",
44433 => "0111100100000000",
44434 => "0111100100000000",
44435 => "0111100100000000",
44436 => "0111100100000000",
44437 => "0111100100000000",
44438 => "0111100100000000",
44439 => "0111100100000000",
44440 => "0111100100000000",
44441 => "0111100100000000",
44442 => "0111100100000000",
44443 => "0111100100000000",
44444 => "0111100100000000",
44445 => "0111100100000000",
44446 => "0111100100000000",
44447 => "0111100100000000",
44448 => "0111100100000000",
44449 => "0111100100000000",
44450 => "0111100100000000",
44451 => "0111100100000000",
44452 => "0111100100000000",
44453 => "0111100100000000",
44454 => "0111100100000000",
44455 => "0111100100000000",
44456 => "0111100100000000",
44457 => "0111100100000000",
44458 => "0111100100000000",
44459 => "0111100100000000",
44460 => "0111100100010000",
44461 => "0111100100010000",
44462 => "0111100100010000",
44463 => "0111100100010000",
44464 => "0111100100010000",
44465 => "0111100100010000",
44466 => "0111100100010000",
44467 => "0111100100010000",
44468 => "0111100100010000",
44469 => "0111100100010000",
44470 => "0111100100010000",
44471 => "0111100100010000",
44472 => "0111100100010000",
44473 => "0111100100010000",
44474 => "0111100100010000",
44475 => "0111100100010000",
44476 => "0111100100010000",
44477 => "0111100100010000",
44478 => "0111100100010000",
44479 => "0111100100010000",
44480 => "0111100100010000",
44481 => "0111100100010000",
44482 => "0111100100010000",
44483 => "0111100100010000",
44484 => "0111100100010000",
44485 => "0111100100010000",
44486 => "0111100100010000",
44487 => "0111100100010000",
44488 => "0111100100010000",
44489 => "0111100100010000",
44490 => "0111100100010000",
44491 => "0111100100010000",
44492 => "0111100100010000",
44493 => "0111100100010000",
44494 => "0111100100010000",
44495 => "0111100100010000",
44496 => "0111100100010000",
44497 => "0111100100010000",
44498 => "0111100100010000",
44499 => "0111100100100000",
44500 => "0111100100100000",
44501 => "0111100100100000",
44502 => "0111100100100000",
44503 => "0111100100100000",
44504 => "0111100100100000",
44505 => "0111100100100000",
44506 => "0111100100100000",
44507 => "0111100100100000",
44508 => "0111100100100000",
44509 => "0111100100100000",
44510 => "0111100100100000",
44511 => "0111100100100000",
44512 => "0111100100100000",
44513 => "0111100100100000",
44514 => "0111100100100000",
44515 => "0111100100100000",
44516 => "0111100100100000",
44517 => "0111100100100000",
44518 => "0111100100100000",
44519 => "0111100100100000",
44520 => "0111100100100000",
44521 => "0111100100100000",
44522 => "0111100100100000",
44523 => "0111100100100000",
44524 => "0111100100100000",
44525 => "0111100100100000",
44526 => "0111100100100000",
44527 => "0111100100100000",
44528 => "0111100100100000",
44529 => "0111100100100000",
44530 => "0111100100100000",
44531 => "0111100100100000",
44532 => "0111100100100000",
44533 => "0111100100100000",
44534 => "0111100100100000",
44535 => "0111100100100000",
44536 => "0111100100100000",
44537 => "0111100100100000",
44538 => "0111100100100000",
44539 => "0111100100110000",
44540 => "0111100100110000",
44541 => "0111100100110000",
44542 => "0111100100110000",
44543 => "0111100100110000",
44544 => "0111100100110000",
44545 => "0111100100110000",
44546 => "0111100100110000",
44547 => "0111100100110000",
44548 => "0111100100110000",
44549 => "0111100100110000",
44550 => "0111100100110000",
44551 => "0111100100110000",
44552 => "0111100100110000",
44553 => "0111100100110000",
44554 => "0111100100110000",
44555 => "0111100100110000",
44556 => "0111100100110000",
44557 => "0111100100110000",
44558 => "0111100100110000",
44559 => "0111100100110000",
44560 => "0111100100110000",
44561 => "0111100100110000",
44562 => "0111100100110000",
44563 => "0111100100110000",
44564 => "0111100100110000",
44565 => "0111100100110000",
44566 => "0111100100110000",
44567 => "0111100100110000",
44568 => "0111100100110000",
44569 => "0111100100110000",
44570 => "0111100100110000",
44571 => "0111100100110000",
44572 => "0111100100110000",
44573 => "0111100100110000",
44574 => "0111100100110000",
44575 => "0111100100110000",
44576 => "0111100100110000",
44577 => "0111100100110000",
44578 => "0111100101000000",
44579 => "0111100101000000",
44580 => "0111100101000000",
44581 => "0111100101000000",
44582 => "0111100101000000",
44583 => "0111100101000000",
44584 => "0111100101000000",
44585 => "0111100101000000",
44586 => "0111100101000000",
44587 => "0111100101000000",
44588 => "0111100101000000",
44589 => "0111100101000000",
44590 => "0111100101000000",
44591 => "0111100101000000",
44592 => "0111100101000000",
44593 => "0111100101000000",
44594 => "0111100101000000",
44595 => "0111100101000000",
44596 => "0111100101000000",
44597 => "0111100101000000",
44598 => "0111100101000000",
44599 => "0111100101000000",
44600 => "0111100101000000",
44601 => "0111100101000000",
44602 => "0111100101000000",
44603 => "0111100101000000",
44604 => "0111100101000000",
44605 => "0111100101000000",
44606 => "0111100101000000",
44607 => "0111100101000000",
44608 => "0111100101000000",
44609 => "0111100101000000",
44610 => "0111100101000000",
44611 => "0111100101000000",
44612 => "0111100101000000",
44613 => "0111100101000000",
44614 => "0111100101000000",
44615 => "0111100101000000",
44616 => "0111100101000000",
44617 => "0111100101000000",
44618 => "0111100101010000",
44619 => "0111100101010000",
44620 => "0111100101010000",
44621 => "0111100101010000",
44622 => "0111100101010000",
44623 => "0111100101010000",
44624 => "0111100101010000",
44625 => "0111100101010000",
44626 => "0111100101010000",
44627 => "0111100101010000",
44628 => "0111100101010000",
44629 => "0111100101010000",
44630 => "0111100101010000",
44631 => "0111100101010000",
44632 => "0111100101010000",
44633 => "0111100101010000",
44634 => "0111100101010000",
44635 => "0111100101010000",
44636 => "0111100101010000",
44637 => "0111100101010000",
44638 => "0111100101010000",
44639 => "0111100101010000",
44640 => "0111100101010000",
44641 => "0111100101010000",
44642 => "0111100101010000",
44643 => "0111100101010000",
44644 => "0111100101010000",
44645 => "0111100101010000",
44646 => "0111100101010000",
44647 => "0111100101010000",
44648 => "0111100101010000",
44649 => "0111100101010000",
44650 => "0111100101010000",
44651 => "0111100101010000",
44652 => "0111100101010000",
44653 => "0111100101010000",
44654 => "0111100101010000",
44655 => "0111100101010000",
44656 => "0111100101010000",
44657 => "0111100101010000",
44658 => "0111100101010000",
44659 => "0111100101100000",
44660 => "0111100101100000",
44661 => "0111100101100000",
44662 => "0111100101100000",
44663 => "0111100101100000",
44664 => "0111100101100000",
44665 => "0111100101100000",
44666 => "0111100101100000",
44667 => "0111100101100000",
44668 => "0111100101100000",
44669 => "0111100101100000",
44670 => "0111100101100000",
44671 => "0111100101100000",
44672 => "0111100101100000",
44673 => "0111100101100000",
44674 => "0111100101100000",
44675 => "0111100101100000",
44676 => "0111100101100000",
44677 => "0111100101100000",
44678 => "0111100101100000",
44679 => "0111100101100000",
44680 => "0111100101100000",
44681 => "0111100101100000",
44682 => "0111100101100000",
44683 => "0111100101100000",
44684 => "0111100101100000",
44685 => "0111100101100000",
44686 => "0111100101100000",
44687 => "0111100101100000",
44688 => "0111100101100000",
44689 => "0111100101100000",
44690 => "0111100101100000",
44691 => "0111100101100000",
44692 => "0111100101100000",
44693 => "0111100101100000",
44694 => "0111100101100000",
44695 => "0111100101100000",
44696 => "0111100101100000",
44697 => "0111100101100000",
44698 => "0111100101100000",
44699 => "0111100101100000",
44700 => "0111100101110000",
44701 => "0111100101110000",
44702 => "0111100101110000",
44703 => "0111100101110000",
44704 => "0111100101110000",
44705 => "0111100101110000",
44706 => "0111100101110000",
44707 => "0111100101110000",
44708 => "0111100101110000",
44709 => "0111100101110000",
44710 => "0111100101110000",
44711 => "0111100101110000",
44712 => "0111100101110000",
44713 => "0111100101110000",
44714 => "0111100101110000",
44715 => "0111100101110000",
44716 => "0111100101110000",
44717 => "0111100101110000",
44718 => "0111100101110000",
44719 => "0111100101110000",
44720 => "0111100101110000",
44721 => "0111100101110000",
44722 => "0111100101110000",
44723 => "0111100101110000",
44724 => "0111100101110000",
44725 => "0111100101110000",
44726 => "0111100101110000",
44727 => "0111100101110000",
44728 => "0111100101110000",
44729 => "0111100101110000",
44730 => "0111100101110000",
44731 => "0111100101110000",
44732 => "0111100101110000",
44733 => "0111100101110000",
44734 => "0111100101110000",
44735 => "0111100101110000",
44736 => "0111100101110000",
44737 => "0111100101110000",
44738 => "0111100101110000",
44739 => "0111100101110000",
44740 => "0111100101110000",
44741 => "0111100110000000",
44742 => "0111100110000000",
44743 => "0111100110000000",
44744 => "0111100110000000",
44745 => "0111100110000000",
44746 => "0111100110000000",
44747 => "0111100110000000",
44748 => "0111100110000000",
44749 => "0111100110000000",
44750 => "0111100110000000",
44751 => "0111100110000000",
44752 => "0111100110000000",
44753 => "0111100110000000",
44754 => "0111100110000000",
44755 => "0111100110000000",
44756 => "0111100110000000",
44757 => "0111100110000000",
44758 => "0111100110000000",
44759 => "0111100110000000",
44760 => "0111100110000000",
44761 => "0111100110000000",
44762 => "0111100110000000",
44763 => "0111100110000000",
44764 => "0111100110000000",
44765 => "0111100110000000",
44766 => "0111100110000000",
44767 => "0111100110000000",
44768 => "0111100110000000",
44769 => "0111100110000000",
44770 => "0111100110000000",
44771 => "0111100110000000",
44772 => "0111100110000000",
44773 => "0111100110000000",
44774 => "0111100110000000",
44775 => "0111100110000000",
44776 => "0111100110000000",
44777 => "0111100110000000",
44778 => "0111100110000000",
44779 => "0111100110000000",
44780 => "0111100110000000",
44781 => "0111100110000000",
44782 => "0111100110010000",
44783 => "0111100110010000",
44784 => "0111100110010000",
44785 => "0111100110010000",
44786 => "0111100110010000",
44787 => "0111100110010000",
44788 => "0111100110010000",
44789 => "0111100110010000",
44790 => "0111100110010000",
44791 => "0111100110010000",
44792 => "0111100110010000",
44793 => "0111100110010000",
44794 => "0111100110010000",
44795 => "0111100110010000",
44796 => "0111100110010000",
44797 => "0111100110010000",
44798 => "0111100110010000",
44799 => "0111100110010000",
44800 => "0111100110010000",
44801 => "0111100110010000",
44802 => "0111100110010000",
44803 => "0111100110010000",
44804 => "0111100110010000",
44805 => "0111100110010000",
44806 => "0111100110010000",
44807 => "0111100110010000",
44808 => "0111100110010000",
44809 => "0111100110010000",
44810 => "0111100110010000",
44811 => "0111100110010000",
44812 => "0111100110010000",
44813 => "0111100110010000",
44814 => "0111100110010000",
44815 => "0111100110010000",
44816 => "0111100110010000",
44817 => "0111100110010000",
44818 => "0111100110010000",
44819 => "0111100110010000",
44820 => "0111100110010000",
44821 => "0111100110010000",
44822 => "0111100110010000",
44823 => "0111100110010000",
44824 => "0111100110100000",
44825 => "0111100110100000",
44826 => "0111100110100000",
44827 => "0111100110100000",
44828 => "0111100110100000",
44829 => "0111100110100000",
44830 => "0111100110100000",
44831 => "0111100110100000",
44832 => "0111100110100000",
44833 => "0111100110100000",
44834 => "0111100110100000",
44835 => "0111100110100000",
44836 => "0111100110100000",
44837 => "0111100110100000",
44838 => "0111100110100000",
44839 => "0111100110100000",
44840 => "0111100110100000",
44841 => "0111100110100000",
44842 => "0111100110100000",
44843 => "0111100110100000",
44844 => "0111100110100000",
44845 => "0111100110100000",
44846 => "0111100110100000",
44847 => "0111100110100000",
44848 => "0111100110100000",
44849 => "0111100110100000",
44850 => "0111100110100000",
44851 => "0111100110100000",
44852 => "0111100110100000",
44853 => "0111100110100000",
44854 => "0111100110100000",
44855 => "0111100110100000",
44856 => "0111100110100000",
44857 => "0111100110100000",
44858 => "0111100110100000",
44859 => "0111100110100000",
44860 => "0111100110100000",
44861 => "0111100110100000",
44862 => "0111100110100000",
44863 => "0111100110100000",
44864 => "0111100110100000",
44865 => "0111100110100000",
44866 => "0111100110110000",
44867 => "0111100110110000",
44868 => "0111100110110000",
44869 => "0111100110110000",
44870 => "0111100110110000",
44871 => "0111100110110000",
44872 => "0111100110110000",
44873 => "0111100110110000",
44874 => "0111100110110000",
44875 => "0111100110110000",
44876 => "0111100110110000",
44877 => "0111100110110000",
44878 => "0111100110110000",
44879 => "0111100110110000",
44880 => "0111100110110000",
44881 => "0111100110110000",
44882 => "0111100110110000",
44883 => "0111100110110000",
44884 => "0111100110110000",
44885 => "0111100110110000",
44886 => "0111100110110000",
44887 => "0111100110110000",
44888 => "0111100110110000",
44889 => "0111100110110000",
44890 => "0111100110110000",
44891 => "0111100110110000",
44892 => "0111100110110000",
44893 => "0111100110110000",
44894 => "0111100110110000",
44895 => "0111100110110000",
44896 => "0111100110110000",
44897 => "0111100110110000",
44898 => "0111100110110000",
44899 => "0111100110110000",
44900 => "0111100110110000",
44901 => "0111100110110000",
44902 => "0111100110110000",
44903 => "0111100110110000",
44904 => "0111100110110000",
44905 => "0111100110110000",
44906 => "0111100110110000",
44907 => "0111100110110000",
44908 => "0111100110110000",
44909 => "0111100111000000",
44910 => "0111100111000000",
44911 => "0111100111000000",
44912 => "0111100111000000",
44913 => "0111100111000000",
44914 => "0111100111000000",
44915 => "0111100111000000",
44916 => "0111100111000000",
44917 => "0111100111000000",
44918 => "0111100111000000",
44919 => "0111100111000000",
44920 => "0111100111000000",
44921 => "0111100111000000",
44922 => "0111100111000000",
44923 => "0111100111000000",
44924 => "0111100111000000",
44925 => "0111100111000000",
44926 => "0111100111000000",
44927 => "0111100111000000",
44928 => "0111100111000000",
44929 => "0111100111000000",
44930 => "0111100111000000",
44931 => "0111100111000000",
44932 => "0111100111000000",
44933 => "0111100111000000",
44934 => "0111100111000000",
44935 => "0111100111000000",
44936 => "0111100111000000",
44937 => "0111100111000000",
44938 => "0111100111000000",
44939 => "0111100111000000",
44940 => "0111100111000000",
44941 => "0111100111000000",
44942 => "0111100111000000",
44943 => "0111100111000000",
44944 => "0111100111000000",
44945 => "0111100111000000",
44946 => "0111100111000000",
44947 => "0111100111000000",
44948 => "0111100111000000",
44949 => "0111100111000000",
44950 => "0111100111000000",
44951 => "0111100111000000",
44952 => "0111100111010000",
44953 => "0111100111010000",
44954 => "0111100111010000",
44955 => "0111100111010000",
44956 => "0111100111010000",
44957 => "0111100111010000",
44958 => "0111100111010000",
44959 => "0111100111010000",
44960 => "0111100111010000",
44961 => "0111100111010000",
44962 => "0111100111010000",
44963 => "0111100111010000",
44964 => "0111100111010000",
44965 => "0111100111010000",
44966 => "0111100111010000",
44967 => "0111100111010000",
44968 => "0111100111010000",
44969 => "0111100111010000",
44970 => "0111100111010000",
44971 => "0111100111010000",
44972 => "0111100111010000",
44973 => "0111100111010000",
44974 => "0111100111010000",
44975 => "0111100111010000",
44976 => "0111100111010000",
44977 => "0111100111010000",
44978 => "0111100111010000",
44979 => "0111100111010000",
44980 => "0111100111010000",
44981 => "0111100111010000",
44982 => "0111100111010000",
44983 => "0111100111010000",
44984 => "0111100111010000",
44985 => "0111100111010000",
44986 => "0111100111010000",
44987 => "0111100111010000",
44988 => "0111100111010000",
44989 => "0111100111010000",
44990 => "0111100111010000",
44991 => "0111100111010000",
44992 => "0111100111010000",
44993 => "0111100111010000",
44994 => "0111100111010000",
44995 => "0111100111100000",
44996 => "0111100111100000",
44997 => "0111100111100000",
44998 => "0111100111100000",
44999 => "0111100111100000",
45000 => "0111100111100000",
45001 => "0111100111100000",
45002 => "0111100111100000",
45003 => "0111100111100000",
45004 => "0111100111100000",
45005 => "0111100111100000",
45006 => "0111100111100000",
45007 => "0111100111100000",
45008 => "0111100111100000",
45009 => "0111100111100000",
45010 => "0111100111100000",
45011 => "0111100111100000",
45012 => "0111100111100000",
45013 => "0111100111100000",
45014 => "0111100111100000",
45015 => "0111100111100000",
45016 => "0111100111100000",
45017 => "0111100111100000",
45018 => "0111100111100000",
45019 => "0111100111100000",
45020 => "0111100111100000",
45021 => "0111100111100000",
45022 => "0111100111100000",
45023 => "0111100111100000",
45024 => "0111100111100000",
45025 => "0111100111100000",
45026 => "0111100111100000",
45027 => "0111100111100000",
45028 => "0111100111100000",
45029 => "0111100111100000",
45030 => "0111100111100000",
45031 => "0111100111100000",
45032 => "0111100111100000",
45033 => "0111100111100000",
45034 => "0111100111100000",
45035 => "0111100111100000",
45036 => "0111100111100000",
45037 => "0111100111100000",
45038 => "0111100111100000",
45039 => "0111100111110000",
45040 => "0111100111110000",
45041 => "0111100111110000",
45042 => "0111100111110000",
45043 => "0111100111110000",
45044 => "0111100111110000",
45045 => "0111100111110000",
45046 => "0111100111110000",
45047 => "0111100111110000",
45048 => "0111100111110000",
45049 => "0111100111110000",
45050 => "0111100111110000",
45051 => "0111100111110000",
45052 => "0111100111110000",
45053 => "0111100111110000",
45054 => "0111100111110000",
45055 => "0111100111110000",
45056 => "0111100111110000",
45057 => "0111100111110000",
45058 => "0111100111110000",
45059 => "0111100111110000",
45060 => "0111100111110000",
45061 => "0111100111110000",
45062 => "0111100111110000",
45063 => "0111100111110000",
45064 => "0111100111110000",
45065 => "0111100111110000",
45066 => "0111100111110000",
45067 => "0111100111110000",
45068 => "0111100111110000",
45069 => "0111100111110000",
45070 => "0111100111110000",
45071 => "0111100111110000",
45072 => "0111100111110000",
45073 => "0111100111110000",
45074 => "0111100111110000",
45075 => "0111100111110000",
45076 => "0111100111110000",
45077 => "0111100111110000",
45078 => "0111100111110000",
45079 => "0111100111110000",
45080 => "0111100111110000",
45081 => "0111100111110000",
45082 => "0111100111110000",
45083 => "0111100111110000",
45084 => "0111101000000000",
45085 => "0111101000000000",
45086 => "0111101000000000",
45087 => "0111101000000000",
45088 => "0111101000000000",
45089 => "0111101000000000",
45090 => "0111101000000000",
45091 => "0111101000000000",
45092 => "0111101000000000",
45093 => "0111101000000000",
45094 => "0111101000000000",
45095 => "0111101000000000",
45096 => "0111101000000000",
45097 => "0111101000000000",
45098 => "0111101000000000",
45099 => "0111101000000000",
45100 => "0111101000000000",
45101 => "0111101000000000",
45102 => "0111101000000000",
45103 => "0111101000000000",
45104 => "0111101000000000",
45105 => "0111101000000000",
45106 => "0111101000000000",
45107 => "0111101000000000",
45108 => "0111101000000000",
45109 => "0111101000000000",
45110 => "0111101000000000",
45111 => "0111101000000000",
45112 => "0111101000000000",
45113 => "0111101000000000",
45114 => "0111101000000000",
45115 => "0111101000000000",
45116 => "0111101000000000",
45117 => "0111101000000000",
45118 => "0111101000000000",
45119 => "0111101000000000",
45120 => "0111101000000000",
45121 => "0111101000000000",
45122 => "0111101000000000",
45123 => "0111101000000000",
45124 => "0111101000000000",
45125 => "0111101000000000",
45126 => "0111101000000000",
45127 => "0111101000000000",
45128 => "0111101000010000",
45129 => "0111101000010000",
45130 => "0111101000010000",
45131 => "0111101000010000",
45132 => "0111101000010000",
45133 => "0111101000010000",
45134 => "0111101000010000",
45135 => "0111101000010000",
45136 => "0111101000010000",
45137 => "0111101000010000",
45138 => "0111101000010000",
45139 => "0111101000010000",
45140 => "0111101000010000",
45141 => "0111101000010000",
45142 => "0111101000010000",
45143 => "0111101000010000",
45144 => "0111101000010000",
45145 => "0111101000010000",
45146 => "0111101000010000",
45147 => "0111101000010000",
45148 => "0111101000010000",
45149 => "0111101000010000",
45150 => "0111101000010000",
45151 => "0111101000010000",
45152 => "0111101000010000",
45153 => "0111101000010000",
45154 => "0111101000010000",
45155 => "0111101000010000",
45156 => "0111101000010000",
45157 => "0111101000010000",
45158 => "0111101000010000",
45159 => "0111101000010000",
45160 => "0111101000010000",
45161 => "0111101000010000",
45162 => "0111101000010000",
45163 => "0111101000010000",
45164 => "0111101000010000",
45165 => "0111101000010000",
45166 => "0111101000010000",
45167 => "0111101000010000",
45168 => "0111101000010000",
45169 => "0111101000010000",
45170 => "0111101000010000",
45171 => "0111101000010000",
45172 => "0111101000010000",
45173 => "0111101000010000",
45174 => "0111101000100000",
45175 => "0111101000100000",
45176 => "0111101000100000",
45177 => "0111101000100000",
45178 => "0111101000100000",
45179 => "0111101000100000",
45180 => "0111101000100000",
45181 => "0111101000100000",
45182 => "0111101000100000",
45183 => "0111101000100000",
45184 => "0111101000100000",
45185 => "0111101000100000",
45186 => "0111101000100000",
45187 => "0111101000100000",
45188 => "0111101000100000",
45189 => "0111101000100000",
45190 => "0111101000100000",
45191 => "0111101000100000",
45192 => "0111101000100000",
45193 => "0111101000100000",
45194 => "0111101000100000",
45195 => "0111101000100000",
45196 => "0111101000100000",
45197 => "0111101000100000",
45198 => "0111101000100000",
45199 => "0111101000100000",
45200 => "0111101000100000",
45201 => "0111101000100000",
45202 => "0111101000100000",
45203 => "0111101000100000",
45204 => "0111101000100000",
45205 => "0111101000100000",
45206 => "0111101000100000",
45207 => "0111101000100000",
45208 => "0111101000100000",
45209 => "0111101000100000",
45210 => "0111101000100000",
45211 => "0111101000100000",
45212 => "0111101000100000",
45213 => "0111101000100000",
45214 => "0111101000100000",
45215 => "0111101000100000",
45216 => "0111101000100000",
45217 => "0111101000100000",
45218 => "0111101000100000",
45219 => "0111101000110000",
45220 => "0111101000110000",
45221 => "0111101000110000",
45222 => "0111101000110000",
45223 => "0111101000110000",
45224 => "0111101000110000",
45225 => "0111101000110000",
45226 => "0111101000110000",
45227 => "0111101000110000",
45228 => "0111101000110000",
45229 => "0111101000110000",
45230 => "0111101000110000",
45231 => "0111101000110000",
45232 => "0111101000110000",
45233 => "0111101000110000",
45234 => "0111101000110000",
45235 => "0111101000110000",
45236 => "0111101000110000",
45237 => "0111101000110000",
45238 => "0111101000110000",
45239 => "0111101000110000",
45240 => "0111101000110000",
45241 => "0111101000110000",
45242 => "0111101000110000",
45243 => "0111101000110000",
45244 => "0111101000110000",
45245 => "0111101000110000",
45246 => "0111101000110000",
45247 => "0111101000110000",
45248 => "0111101000110000",
45249 => "0111101000110000",
45250 => "0111101000110000",
45251 => "0111101000110000",
45252 => "0111101000110000",
45253 => "0111101000110000",
45254 => "0111101000110000",
45255 => "0111101000110000",
45256 => "0111101000110000",
45257 => "0111101000110000",
45258 => "0111101000110000",
45259 => "0111101000110000",
45260 => "0111101000110000",
45261 => "0111101000110000",
45262 => "0111101000110000",
45263 => "0111101000110000",
45264 => "0111101000110000",
45265 => "0111101001000000",
45266 => "0111101001000000",
45267 => "0111101001000000",
45268 => "0111101001000000",
45269 => "0111101001000000",
45270 => "0111101001000000",
45271 => "0111101001000000",
45272 => "0111101001000000",
45273 => "0111101001000000",
45274 => "0111101001000000",
45275 => "0111101001000000",
45276 => "0111101001000000",
45277 => "0111101001000000",
45278 => "0111101001000000",
45279 => "0111101001000000",
45280 => "0111101001000000",
45281 => "0111101001000000",
45282 => "0111101001000000",
45283 => "0111101001000000",
45284 => "0111101001000000",
45285 => "0111101001000000",
45286 => "0111101001000000",
45287 => "0111101001000000",
45288 => "0111101001000000",
45289 => "0111101001000000",
45290 => "0111101001000000",
45291 => "0111101001000000",
45292 => "0111101001000000",
45293 => "0111101001000000",
45294 => "0111101001000000",
45295 => "0111101001000000",
45296 => "0111101001000000",
45297 => "0111101001000000",
45298 => "0111101001000000",
45299 => "0111101001000000",
45300 => "0111101001000000",
45301 => "0111101001000000",
45302 => "0111101001000000",
45303 => "0111101001000000",
45304 => "0111101001000000",
45305 => "0111101001000000",
45306 => "0111101001000000",
45307 => "0111101001000000",
45308 => "0111101001000000",
45309 => "0111101001000000",
45310 => "0111101001000000",
45311 => "0111101001000000",
45312 => "0111101001010000",
45313 => "0111101001010000",
45314 => "0111101001010000",
45315 => "0111101001010000",
45316 => "0111101001010000",
45317 => "0111101001010000",
45318 => "0111101001010000",
45319 => "0111101001010000",
45320 => "0111101001010000",
45321 => "0111101001010000",
45322 => "0111101001010000",
45323 => "0111101001010000",
45324 => "0111101001010000",
45325 => "0111101001010000",
45326 => "0111101001010000",
45327 => "0111101001010000",
45328 => "0111101001010000",
45329 => "0111101001010000",
45330 => "0111101001010000",
45331 => "0111101001010000",
45332 => "0111101001010000",
45333 => "0111101001010000",
45334 => "0111101001010000",
45335 => "0111101001010000",
45336 => "0111101001010000",
45337 => "0111101001010000",
45338 => "0111101001010000",
45339 => "0111101001010000",
45340 => "0111101001010000",
45341 => "0111101001010000",
45342 => "0111101001010000",
45343 => "0111101001010000",
45344 => "0111101001010000",
45345 => "0111101001010000",
45346 => "0111101001010000",
45347 => "0111101001010000",
45348 => "0111101001010000",
45349 => "0111101001010000",
45350 => "0111101001010000",
45351 => "0111101001010000",
45352 => "0111101001010000",
45353 => "0111101001010000",
45354 => "0111101001010000",
45355 => "0111101001010000",
45356 => "0111101001010000",
45357 => "0111101001010000",
45358 => "0111101001010000",
45359 => "0111101001100000",
45360 => "0111101001100000",
45361 => "0111101001100000",
45362 => "0111101001100000",
45363 => "0111101001100000",
45364 => "0111101001100000",
45365 => "0111101001100000",
45366 => "0111101001100000",
45367 => "0111101001100000",
45368 => "0111101001100000",
45369 => "0111101001100000",
45370 => "0111101001100000",
45371 => "0111101001100000",
45372 => "0111101001100000",
45373 => "0111101001100000",
45374 => "0111101001100000",
45375 => "0111101001100000",
45376 => "0111101001100000",
45377 => "0111101001100000",
45378 => "0111101001100000",
45379 => "0111101001100000",
45380 => "0111101001100000",
45381 => "0111101001100000",
45382 => "0111101001100000",
45383 => "0111101001100000",
45384 => "0111101001100000",
45385 => "0111101001100000",
45386 => "0111101001100000",
45387 => "0111101001100000",
45388 => "0111101001100000",
45389 => "0111101001100000",
45390 => "0111101001100000",
45391 => "0111101001100000",
45392 => "0111101001100000",
45393 => "0111101001100000",
45394 => "0111101001100000",
45395 => "0111101001100000",
45396 => "0111101001100000",
45397 => "0111101001100000",
45398 => "0111101001100000",
45399 => "0111101001100000",
45400 => "0111101001100000",
45401 => "0111101001100000",
45402 => "0111101001100000",
45403 => "0111101001100000",
45404 => "0111101001100000",
45405 => "0111101001100000",
45406 => "0111101001100000",
45407 => "0111101001110000",
45408 => "0111101001110000",
45409 => "0111101001110000",
45410 => "0111101001110000",
45411 => "0111101001110000",
45412 => "0111101001110000",
45413 => "0111101001110000",
45414 => "0111101001110000",
45415 => "0111101001110000",
45416 => "0111101001110000",
45417 => "0111101001110000",
45418 => "0111101001110000",
45419 => "0111101001110000",
45420 => "0111101001110000",
45421 => "0111101001110000",
45422 => "0111101001110000",
45423 => "0111101001110000",
45424 => "0111101001110000",
45425 => "0111101001110000",
45426 => "0111101001110000",
45427 => "0111101001110000",
45428 => "0111101001110000",
45429 => "0111101001110000",
45430 => "0111101001110000",
45431 => "0111101001110000",
45432 => "0111101001110000",
45433 => "0111101001110000",
45434 => "0111101001110000",
45435 => "0111101001110000",
45436 => "0111101001110000",
45437 => "0111101001110000",
45438 => "0111101001110000",
45439 => "0111101001110000",
45440 => "0111101001110000",
45441 => "0111101001110000",
45442 => "0111101001110000",
45443 => "0111101001110000",
45444 => "0111101001110000",
45445 => "0111101001110000",
45446 => "0111101001110000",
45447 => "0111101001110000",
45448 => "0111101001110000",
45449 => "0111101001110000",
45450 => "0111101001110000",
45451 => "0111101001110000",
45452 => "0111101001110000",
45453 => "0111101001110000",
45454 => "0111101001110000",
45455 => "0111101010000000",
45456 => "0111101010000000",
45457 => "0111101010000000",
45458 => "0111101010000000",
45459 => "0111101010000000",
45460 => "0111101010000000",
45461 => "0111101010000000",
45462 => "0111101010000000",
45463 => "0111101010000000",
45464 => "0111101010000000",
45465 => "0111101010000000",
45466 => "0111101010000000",
45467 => "0111101010000000",
45468 => "0111101010000000",
45469 => "0111101010000000",
45470 => "0111101010000000",
45471 => "0111101010000000",
45472 => "0111101010000000",
45473 => "0111101010000000",
45474 => "0111101010000000",
45475 => "0111101010000000",
45476 => "0111101010000000",
45477 => "0111101010000000",
45478 => "0111101010000000",
45479 => "0111101010000000",
45480 => "0111101010000000",
45481 => "0111101010000000",
45482 => "0111101010000000",
45483 => "0111101010000000",
45484 => "0111101010000000",
45485 => "0111101010000000",
45486 => "0111101010000000",
45487 => "0111101010000000",
45488 => "0111101010000000",
45489 => "0111101010000000",
45490 => "0111101010000000",
45491 => "0111101010000000",
45492 => "0111101010000000",
45493 => "0111101010000000",
45494 => "0111101010000000",
45495 => "0111101010000000",
45496 => "0111101010000000",
45497 => "0111101010000000",
45498 => "0111101010000000",
45499 => "0111101010000000",
45500 => "0111101010000000",
45501 => "0111101010000000",
45502 => "0111101010000000",
45503 => "0111101010000000",
45504 => "0111101010010000",
45505 => "0111101010010000",
45506 => "0111101010010000",
45507 => "0111101010010000",
45508 => "0111101010010000",
45509 => "0111101010010000",
45510 => "0111101010010000",
45511 => "0111101010010000",
45512 => "0111101010010000",
45513 => "0111101010010000",
45514 => "0111101010010000",
45515 => "0111101010010000",
45516 => "0111101010010000",
45517 => "0111101010010000",
45518 => "0111101010010000",
45519 => "0111101010010000",
45520 => "0111101010010000",
45521 => "0111101010010000",
45522 => "0111101010010000",
45523 => "0111101010010000",
45524 => "0111101010010000",
45525 => "0111101010010000",
45526 => "0111101010010000",
45527 => "0111101010010000",
45528 => "0111101010010000",
45529 => "0111101010010000",
45530 => "0111101010010000",
45531 => "0111101010010000",
45532 => "0111101010010000",
45533 => "0111101010010000",
45534 => "0111101010010000",
45535 => "0111101010010000",
45536 => "0111101010010000",
45537 => "0111101010010000",
45538 => "0111101010010000",
45539 => "0111101010010000",
45540 => "0111101010010000",
45541 => "0111101010010000",
45542 => "0111101010010000",
45543 => "0111101010010000",
45544 => "0111101010010000",
45545 => "0111101010010000",
45546 => "0111101010010000",
45547 => "0111101010010000",
45548 => "0111101010010000",
45549 => "0111101010010000",
45550 => "0111101010010000",
45551 => "0111101010010000",
45552 => "0111101010010000",
45553 => "0111101010100000",
45554 => "0111101010100000",
45555 => "0111101010100000",
45556 => "0111101010100000",
45557 => "0111101010100000",
45558 => "0111101010100000",
45559 => "0111101010100000",
45560 => "0111101010100000",
45561 => "0111101010100000",
45562 => "0111101010100000",
45563 => "0111101010100000",
45564 => "0111101010100000",
45565 => "0111101010100000",
45566 => "0111101010100000",
45567 => "0111101010100000",
45568 => "0111101010100000",
45569 => "0111101010100000",
45570 => "0111101010100000",
45571 => "0111101010100000",
45572 => "0111101010100000",
45573 => "0111101010100000",
45574 => "0111101010100000",
45575 => "0111101010100000",
45576 => "0111101010100000",
45577 => "0111101010100000",
45578 => "0111101010100000",
45579 => "0111101010100000",
45580 => "0111101010100000",
45581 => "0111101010100000",
45582 => "0111101010100000",
45583 => "0111101010100000",
45584 => "0111101010100000",
45585 => "0111101010100000",
45586 => "0111101010100000",
45587 => "0111101010100000",
45588 => "0111101010100000",
45589 => "0111101010100000",
45590 => "0111101010100000",
45591 => "0111101010100000",
45592 => "0111101010100000",
45593 => "0111101010100000",
45594 => "0111101010100000",
45595 => "0111101010100000",
45596 => "0111101010100000",
45597 => "0111101010100000",
45598 => "0111101010100000",
45599 => "0111101010100000",
45600 => "0111101010100000",
45601 => "0111101010100000",
45602 => "0111101010110000",
45603 => "0111101010110000",
45604 => "0111101010110000",
45605 => "0111101010110000",
45606 => "0111101010110000",
45607 => "0111101010110000",
45608 => "0111101010110000",
45609 => "0111101010110000",
45610 => "0111101010110000",
45611 => "0111101010110000",
45612 => "0111101010110000",
45613 => "0111101010110000",
45614 => "0111101010110000",
45615 => "0111101010110000",
45616 => "0111101010110000",
45617 => "0111101010110000",
45618 => "0111101010110000",
45619 => "0111101010110000",
45620 => "0111101010110000",
45621 => "0111101010110000",
45622 => "0111101010110000",
45623 => "0111101010110000",
45624 => "0111101010110000",
45625 => "0111101010110000",
45626 => "0111101010110000",
45627 => "0111101010110000",
45628 => "0111101010110000",
45629 => "0111101010110000",
45630 => "0111101010110000",
45631 => "0111101010110000",
45632 => "0111101010110000",
45633 => "0111101010110000",
45634 => "0111101010110000",
45635 => "0111101010110000",
45636 => "0111101010110000",
45637 => "0111101010110000",
45638 => "0111101010110000",
45639 => "0111101010110000",
45640 => "0111101010110000",
45641 => "0111101010110000",
45642 => "0111101010110000",
45643 => "0111101010110000",
45644 => "0111101010110000",
45645 => "0111101010110000",
45646 => "0111101010110000",
45647 => "0111101010110000",
45648 => "0111101010110000",
45649 => "0111101010110000",
45650 => "0111101010110000",
45651 => "0111101010110000",
45652 => "0111101010110000",
45653 => "0111101011000000",
45654 => "0111101011000000",
45655 => "0111101011000000",
45656 => "0111101011000000",
45657 => "0111101011000000",
45658 => "0111101011000000",
45659 => "0111101011000000",
45660 => "0111101011000000",
45661 => "0111101011000000",
45662 => "0111101011000000",
45663 => "0111101011000000",
45664 => "0111101011000000",
45665 => "0111101011000000",
45666 => "0111101011000000",
45667 => "0111101011000000",
45668 => "0111101011000000",
45669 => "0111101011000000",
45670 => "0111101011000000",
45671 => "0111101011000000",
45672 => "0111101011000000",
45673 => "0111101011000000",
45674 => "0111101011000000",
45675 => "0111101011000000",
45676 => "0111101011000000",
45677 => "0111101011000000",
45678 => "0111101011000000",
45679 => "0111101011000000",
45680 => "0111101011000000",
45681 => "0111101011000000",
45682 => "0111101011000000",
45683 => "0111101011000000",
45684 => "0111101011000000",
45685 => "0111101011000000",
45686 => "0111101011000000",
45687 => "0111101011000000",
45688 => "0111101011000000",
45689 => "0111101011000000",
45690 => "0111101011000000",
45691 => "0111101011000000",
45692 => "0111101011000000",
45693 => "0111101011000000",
45694 => "0111101011000000",
45695 => "0111101011000000",
45696 => "0111101011000000",
45697 => "0111101011000000",
45698 => "0111101011000000",
45699 => "0111101011000000",
45700 => "0111101011000000",
45701 => "0111101011000000",
45702 => "0111101011000000",
45703 => "0111101011000000",
45704 => "0111101011010000",
45705 => "0111101011010000",
45706 => "0111101011010000",
45707 => "0111101011010000",
45708 => "0111101011010000",
45709 => "0111101011010000",
45710 => "0111101011010000",
45711 => "0111101011010000",
45712 => "0111101011010000",
45713 => "0111101011010000",
45714 => "0111101011010000",
45715 => "0111101011010000",
45716 => "0111101011010000",
45717 => "0111101011010000",
45718 => "0111101011010000",
45719 => "0111101011010000",
45720 => "0111101011010000",
45721 => "0111101011010000",
45722 => "0111101011010000",
45723 => "0111101011010000",
45724 => "0111101011010000",
45725 => "0111101011010000",
45726 => "0111101011010000",
45727 => "0111101011010000",
45728 => "0111101011010000",
45729 => "0111101011010000",
45730 => "0111101011010000",
45731 => "0111101011010000",
45732 => "0111101011010000",
45733 => "0111101011010000",
45734 => "0111101011010000",
45735 => "0111101011010000",
45736 => "0111101011010000",
45737 => "0111101011010000",
45738 => "0111101011010000",
45739 => "0111101011010000",
45740 => "0111101011010000",
45741 => "0111101011010000",
45742 => "0111101011010000",
45743 => "0111101011010000",
45744 => "0111101011010000",
45745 => "0111101011010000",
45746 => "0111101011010000",
45747 => "0111101011010000",
45748 => "0111101011010000",
45749 => "0111101011010000",
45750 => "0111101011010000",
45751 => "0111101011010000",
45752 => "0111101011010000",
45753 => "0111101011010000",
45754 => "0111101011010000",
45755 => "0111101011100000",
45756 => "0111101011100000",
45757 => "0111101011100000",
45758 => "0111101011100000",
45759 => "0111101011100000",
45760 => "0111101011100000",
45761 => "0111101011100000",
45762 => "0111101011100000",
45763 => "0111101011100000",
45764 => "0111101011100000",
45765 => "0111101011100000",
45766 => "0111101011100000",
45767 => "0111101011100000",
45768 => "0111101011100000",
45769 => "0111101011100000",
45770 => "0111101011100000",
45771 => "0111101011100000",
45772 => "0111101011100000",
45773 => "0111101011100000",
45774 => "0111101011100000",
45775 => "0111101011100000",
45776 => "0111101011100000",
45777 => "0111101011100000",
45778 => "0111101011100000",
45779 => "0111101011100000",
45780 => "0111101011100000",
45781 => "0111101011100000",
45782 => "0111101011100000",
45783 => "0111101011100000",
45784 => "0111101011100000",
45785 => "0111101011100000",
45786 => "0111101011100000",
45787 => "0111101011100000",
45788 => "0111101011100000",
45789 => "0111101011100000",
45790 => "0111101011100000",
45791 => "0111101011100000",
45792 => "0111101011100000",
45793 => "0111101011100000",
45794 => "0111101011100000",
45795 => "0111101011100000",
45796 => "0111101011100000",
45797 => "0111101011100000",
45798 => "0111101011100000",
45799 => "0111101011100000",
45800 => "0111101011100000",
45801 => "0111101011100000",
45802 => "0111101011100000",
45803 => "0111101011100000",
45804 => "0111101011100000",
45805 => "0111101011100000",
45806 => "0111101011100000",
45807 => "0111101011110000",
45808 => "0111101011110000",
45809 => "0111101011110000",
45810 => "0111101011110000",
45811 => "0111101011110000",
45812 => "0111101011110000",
45813 => "0111101011110000",
45814 => "0111101011110000",
45815 => "0111101011110000",
45816 => "0111101011110000",
45817 => "0111101011110000",
45818 => "0111101011110000",
45819 => "0111101011110000",
45820 => "0111101011110000",
45821 => "0111101011110000",
45822 => "0111101011110000",
45823 => "0111101011110000",
45824 => "0111101011110000",
45825 => "0111101011110000",
45826 => "0111101011110000",
45827 => "0111101011110000",
45828 => "0111101011110000",
45829 => "0111101011110000",
45830 => "0111101011110000",
45831 => "0111101011110000",
45832 => "0111101011110000",
45833 => "0111101011110000",
45834 => "0111101011110000",
45835 => "0111101011110000",
45836 => "0111101011110000",
45837 => "0111101011110000",
45838 => "0111101011110000",
45839 => "0111101011110000",
45840 => "0111101011110000",
45841 => "0111101011110000",
45842 => "0111101011110000",
45843 => "0111101011110000",
45844 => "0111101011110000",
45845 => "0111101011110000",
45846 => "0111101011110000",
45847 => "0111101011110000",
45848 => "0111101011110000",
45849 => "0111101011110000",
45850 => "0111101011110000",
45851 => "0111101011110000",
45852 => "0111101011110000",
45853 => "0111101011110000",
45854 => "0111101011110000",
45855 => "0111101011110000",
45856 => "0111101011110000",
45857 => "0111101011110000",
45858 => "0111101011110000",
45859 => "0111101011110000",
45860 => "0111101100000000",
45861 => "0111101100000000",
45862 => "0111101100000000",
45863 => "0111101100000000",
45864 => "0111101100000000",
45865 => "0111101100000000",
45866 => "0111101100000000",
45867 => "0111101100000000",
45868 => "0111101100000000",
45869 => "0111101100000000",
45870 => "0111101100000000",
45871 => "0111101100000000",
45872 => "0111101100000000",
45873 => "0111101100000000",
45874 => "0111101100000000",
45875 => "0111101100000000",
45876 => "0111101100000000",
45877 => "0111101100000000",
45878 => "0111101100000000",
45879 => "0111101100000000",
45880 => "0111101100000000",
45881 => "0111101100000000",
45882 => "0111101100000000",
45883 => "0111101100000000",
45884 => "0111101100000000",
45885 => "0111101100000000",
45886 => "0111101100000000",
45887 => "0111101100000000",
45888 => "0111101100000000",
45889 => "0111101100000000",
45890 => "0111101100000000",
45891 => "0111101100000000",
45892 => "0111101100000000",
45893 => "0111101100000000",
45894 => "0111101100000000",
45895 => "0111101100000000",
45896 => "0111101100000000",
45897 => "0111101100000000",
45898 => "0111101100000000",
45899 => "0111101100000000",
45900 => "0111101100000000",
45901 => "0111101100000000",
45902 => "0111101100000000",
45903 => "0111101100000000",
45904 => "0111101100000000",
45905 => "0111101100000000",
45906 => "0111101100000000",
45907 => "0111101100000000",
45908 => "0111101100000000",
45909 => "0111101100000000",
45910 => "0111101100000000",
45911 => "0111101100000000",
45912 => "0111101100000000",
45913 => "0111101100010000",
45914 => "0111101100010000",
45915 => "0111101100010000",
45916 => "0111101100010000",
45917 => "0111101100010000",
45918 => "0111101100010000",
45919 => "0111101100010000",
45920 => "0111101100010000",
45921 => "0111101100010000",
45922 => "0111101100010000",
45923 => "0111101100010000",
45924 => "0111101100010000",
45925 => "0111101100010000",
45926 => "0111101100010000",
45927 => "0111101100010000",
45928 => "0111101100010000",
45929 => "0111101100010000",
45930 => "0111101100010000",
45931 => "0111101100010000",
45932 => "0111101100010000",
45933 => "0111101100010000",
45934 => "0111101100010000",
45935 => "0111101100010000",
45936 => "0111101100010000",
45937 => "0111101100010000",
45938 => "0111101100010000",
45939 => "0111101100010000",
45940 => "0111101100010000",
45941 => "0111101100010000",
45942 => "0111101100010000",
45943 => "0111101100010000",
45944 => "0111101100010000",
45945 => "0111101100010000",
45946 => "0111101100010000",
45947 => "0111101100010000",
45948 => "0111101100010000",
45949 => "0111101100010000",
45950 => "0111101100010000",
45951 => "0111101100010000",
45952 => "0111101100010000",
45953 => "0111101100010000",
45954 => "0111101100010000",
45955 => "0111101100010000",
45956 => "0111101100010000",
45957 => "0111101100010000",
45958 => "0111101100010000",
45959 => "0111101100010000",
45960 => "0111101100010000",
45961 => "0111101100010000",
45962 => "0111101100010000",
45963 => "0111101100010000",
45964 => "0111101100010000",
45965 => "0111101100010000",
45966 => "0111101100010000",
45967 => "0111101100100000",
45968 => "0111101100100000",
45969 => "0111101100100000",
45970 => "0111101100100000",
45971 => "0111101100100000",
45972 => "0111101100100000",
45973 => "0111101100100000",
45974 => "0111101100100000",
45975 => "0111101100100000",
45976 => "0111101100100000",
45977 => "0111101100100000",
45978 => "0111101100100000",
45979 => "0111101100100000",
45980 => "0111101100100000",
45981 => "0111101100100000",
45982 => "0111101100100000",
45983 => "0111101100100000",
45984 => "0111101100100000",
45985 => "0111101100100000",
45986 => "0111101100100000",
45987 => "0111101100100000",
45988 => "0111101100100000",
45989 => "0111101100100000",
45990 => "0111101100100000",
45991 => "0111101100100000",
45992 => "0111101100100000",
45993 => "0111101100100000",
45994 => "0111101100100000",
45995 => "0111101100100000",
45996 => "0111101100100000",
45997 => "0111101100100000",
45998 => "0111101100100000",
45999 => "0111101100100000",
46000 => "0111101100100000",
46001 => "0111101100100000",
46002 => "0111101100100000",
46003 => "0111101100100000",
46004 => "0111101100100000",
46005 => "0111101100100000",
46006 => "0111101100100000",
46007 => "0111101100100000",
46008 => "0111101100100000",
46009 => "0111101100100000",
46010 => "0111101100100000",
46011 => "0111101100100000",
46012 => "0111101100100000",
46013 => "0111101100100000",
46014 => "0111101100100000",
46015 => "0111101100100000",
46016 => "0111101100100000",
46017 => "0111101100100000",
46018 => "0111101100100000",
46019 => "0111101100100000",
46020 => "0111101100100000",
46021 => "0111101100110000",
46022 => "0111101100110000",
46023 => "0111101100110000",
46024 => "0111101100110000",
46025 => "0111101100110000",
46026 => "0111101100110000",
46027 => "0111101100110000",
46028 => "0111101100110000",
46029 => "0111101100110000",
46030 => "0111101100110000",
46031 => "0111101100110000",
46032 => "0111101100110000",
46033 => "0111101100110000",
46034 => "0111101100110000",
46035 => "0111101100110000",
46036 => "0111101100110000",
46037 => "0111101100110000",
46038 => "0111101100110000",
46039 => "0111101100110000",
46040 => "0111101100110000",
46041 => "0111101100110000",
46042 => "0111101100110000",
46043 => "0111101100110000",
46044 => "0111101100110000",
46045 => "0111101100110000",
46046 => "0111101100110000",
46047 => "0111101100110000",
46048 => "0111101100110000",
46049 => "0111101100110000",
46050 => "0111101100110000",
46051 => "0111101100110000",
46052 => "0111101100110000",
46053 => "0111101100110000",
46054 => "0111101100110000",
46055 => "0111101100110000",
46056 => "0111101100110000",
46057 => "0111101100110000",
46058 => "0111101100110000",
46059 => "0111101100110000",
46060 => "0111101100110000",
46061 => "0111101100110000",
46062 => "0111101100110000",
46063 => "0111101100110000",
46064 => "0111101100110000",
46065 => "0111101100110000",
46066 => "0111101100110000",
46067 => "0111101100110000",
46068 => "0111101100110000",
46069 => "0111101100110000",
46070 => "0111101100110000",
46071 => "0111101100110000",
46072 => "0111101100110000",
46073 => "0111101100110000",
46074 => "0111101100110000",
46075 => "0111101100110000",
46076 => "0111101100110000",
46077 => "0111101101000000",
46078 => "0111101101000000",
46079 => "0111101101000000",
46080 => "0111101101000000",
46081 => "0111101101000000",
46082 => "0111101101000000",
46083 => "0111101101000000",
46084 => "0111101101000000",
46085 => "0111101101000000",
46086 => "0111101101000000",
46087 => "0111101101000000",
46088 => "0111101101000000",
46089 => "0111101101000000",
46090 => "0111101101000000",
46091 => "0111101101000000",
46092 => "0111101101000000",
46093 => "0111101101000000",
46094 => "0111101101000000",
46095 => "0111101101000000",
46096 => "0111101101000000",
46097 => "0111101101000000",
46098 => "0111101101000000",
46099 => "0111101101000000",
46100 => "0111101101000000",
46101 => "0111101101000000",
46102 => "0111101101000000",
46103 => "0111101101000000",
46104 => "0111101101000000",
46105 => "0111101101000000",
46106 => "0111101101000000",
46107 => "0111101101000000",
46108 => "0111101101000000",
46109 => "0111101101000000",
46110 => "0111101101000000",
46111 => "0111101101000000",
46112 => "0111101101000000",
46113 => "0111101101000000",
46114 => "0111101101000000",
46115 => "0111101101000000",
46116 => "0111101101000000",
46117 => "0111101101000000",
46118 => "0111101101000000",
46119 => "0111101101000000",
46120 => "0111101101000000",
46121 => "0111101101000000",
46122 => "0111101101000000",
46123 => "0111101101000000",
46124 => "0111101101000000",
46125 => "0111101101000000",
46126 => "0111101101000000",
46127 => "0111101101000000",
46128 => "0111101101000000",
46129 => "0111101101000000",
46130 => "0111101101000000",
46131 => "0111101101000000",
46132 => "0111101101000000",
46133 => "0111101101010000",
46134 => "0111101101010000",
46135 => "0111101101010000",
46136 => "0111101101010000",
46137 => "0111101101010000",
46138 => "0111101101010000",
46139 => "0111101101010000",
46140 => "0111101101010000",
46141 => "0111101101010000",
46142 => "0111101101010000",
46143 => "0111101101010000",
46144 => "0111101101010000",
46145 => "0111101101010000",
46146 => "0111101101010000",
46147 => "0111101101010000",
46148 => "0111101101010000",
46149 => "0111101101010000",
46150 => "0111101101010000",
46151 => "0111101101010000",
46152 => "0111101101010000",
46153 => "0111101101010000",
46154 => "0111101101010000",
46155 => "0111101101010000",
46156 => "0111101101010000",
46157 => "0111101101010000",
46158 => "0111101101010000",
46159 => "0111101101010000",
46160 => "0111101101010000",
46161 => "0111101101010000",
46162 => "0111101101010000",
46163 => "0111101101010000",
46164 => "0111101101010000",
46165 => "0111101101010000",
46166 => "0111101101010000",
46167 => "0111101101010000",
46168 => "0111101101010000",
46169 => "0111101101010000",
46170 => "0111101101010000",
46171 => "0111101101010000",
46172 => "0111101101010000",
46173 => "0111101101010000",
46174 => "0111101101010000",
46175 => "0111101101010000",
46176 => "0111101101010000",
46177 => "0111101101010000",
46178 => "0111101101010000",
46179 => "0111101101010000",
46180 => "0111101101010000",
46181 => "0111101101010000",
46182 => "0111101101010000",
46183 => "0111101101010000",
46184 => "0111101101010000",
46185 => "0111101101010000",
46186 => "0111101101010000",
46187 => "0111101101010000",
46188 => "0111101101010000",
46189 => "0111101101100000",
46190 => "0111101101100000",
46191 => "0111101101100000",
46192 => "0111101101100000",
46193 => "0111101101100000",
46194 => "0111101101100000",
46195 => "0111101101100000",
46196 => "0111101101100000",
46197 => "0111101101100000",
46198 => "0111101101100000",
46199 => "0111101101100000",
46200 => "0111101101100000",
46201 => "0111101101100000",
46202 => "0111101101100000",
46203 => "0111101101100000",
46204 => "0111101101100000",
46205 => "0111101101100000",
46206 => "0111101101100000",
46207 => "0111101101100000",
46208 => "0111101101100000",
46209 => "0111101101100000",
46210 => "0111101101100000",
46211 => "0111101101100000",
46212 => "0111101101100000",
46213 => "0111101101100000",
46214 => "0111101101100000",
46215 => "0111101101100000",
46216 => "0111101101100000",
46217 => "0111101101100000",
46218 => "0111101101100000",
46219 => "0111101101100000",
46220 => "0111101101100000",
46221 => "0111101101100000",
46222 => "0111101101100000",
46223 => "0111101101100000",
46224 => "0111101101100000",
46225 => "0111101101100000",
46226 => "0111101101100000",
46227 => "0111101101100000",
46228 => "0111101101100000",
46229 => "0111101101100000",
46230 => "0111101101100000",
46231 => "0111101101100000",
46232 => "0111101101100000",
46233 => "0111101101100000",
46234 => "0111101101100000",
46235 => "0111101101100000",
46236 => "0111101101100000",
46237 => "0111101101100000",
46238 => "0111101101100000",
46239 => "0111101101100000",
46240 => "0111101101100000",
46241 => "0111101101100000",
46242 => "0111101101100000",
46243 => "0111101101100000",
46244 => "0111101101100000",
46245 => "0111101101100000",
46246 => "0111101101100000",
46247 => "0111101101110000",
46248 => "0111101101110000",
46249 => "0111101101110000",
46250 => "0111101101110000",
46251 => "0111101101110000",
46252 => "0111101101110000",
46253 => "0111101101110000",
46254 => "0111101101110000",
46255 => "0111101101110000",
46256 => "0111101101110000",
46257 => "0111101101110000",
46258 => "0111101101110000",
46259 => "0111101101110000",
46260 => "0111101101110000",
46261 => "0111101101110000",
46262 => "0111101101110000",
46263 => "0111101101110000",
46264 => "0111101101110000",
46265 => "0111101101110000",
46266 => "0111101101110000",
46267 => "0111101101110000",
46268 => "0111101101110000",
46269 => "0111101101110000",
46270 => "0111101101110000",
46271 => "0111101101110000",
46272 => "0111101101110000",
46273 => "0111101101110000",
46274 => "0111101101110000",
46275 => "0111101101110000",
46276 => "0111101101110000",
46277 => "0111101101110000",
46278 => "0111101101110000",
46279 => "0111101101110000",
46280 => "0111101101110000",
46281 => "0111101101110000",
46282 => "0111101101110000",
46283 => "0111101101110000",
46284 => "0111101101110000",
46285 => "0111101101110000",
46286 => "0111101101110000",
46287 => "0111101101110000",
46288 => "0111101101110000",
46289 => "0111101101110000",
46290 => "0111101101110000",
46291 => "0111101101110000",
46292 => "0111101101110000",
46293 => "0111101101110000",
46294 => "0111101101110000",
46295 => "0111101101110000",
46296 => "0111101101110000",
46297 => "0111101101110000",
46298 => "0111101101110000",
46299 => "0111101101110000",
46300 => "0111101101110000",
46301 => "0111101101110000",
46302 => "0111101101110000",
46303 => "0111101101110000",
46304 => "0111101101110000",
46305 => "0111101110000000",
46306 => "0111101110000000",
46307 => "0111101110000000",
46308 => "0111101110000000",
46309 => "0111101110000000",
46310 => "0111101110000000",
46311 => "0111101110000000",
46312 => "0111101110000000",
46313 => "0111101110000000",
46314 => "0111101110000000",
46315 => "0111101110000000",
46316 => "0111101110000000",
46317 => "0111101110000000",
46318 => "0111101110000000",
46319 => "0111101110000000",
46320 => "0111101110000000",
46321 => "0111101110000000",
46322 => "0111101110000000",
46323 => "0111101110000000",
46324 => "0111101110000000",
46325 => "0111101110000000",
46326 => "0111101110000000",
46327 => "0111101110000000",
46328 => "0111101110000000",
46329 => "0111101110000000",
46330 => "0111101110000000",
46331 => "0111101110000000",
46332 => "0111101110000000",
46333 => "0111101110000000",
46334 => "0111101110000000",
46335 => "0111101110000000",
46336 => "0111101110000000",
46337 => "0111101110000000",
46338 => "0111101110000000",
46339 => "0111101110000000",
46340 => "0111101110000000",
46341 => "0111101110000000",
46342 => "0111101110000000",
46343 => "0111101110000000",
46344 => "0111101110000000",
46345 => "0111101110000000",
46346 => "0111101110000000",
46347 => "0111101110000000",
46348 => "0111101110000000",
46349 => "0111101110000000",
46350 => "0111101110000000",
46351 => "0111101110000000",
46352 => "0111101110000000",
46353 => "0111101110000000",
46354 => "0111101110000000",
46355 => "0111101110000000",
46356 => "0111101110000000",
46357 => "0111101110000000",
46358 => "0111101110000000",
46359 => "0111101110000000",
46360 => "0111101110000000",
46361 => "0111101110000000",
46362 => "0111101110000000",
46363 => "0111101110000000",
46364 => "0111101110010000",
46365 => "0111101110010000",
46366 => "0111101110010000",
46367 => "0111101110010000",
46368 => "0111101110010000",
46369 => "0111101110010000",
46370 => "0111101110010000",
46371 => "0111101110010000",
46372 => "0111101110010000",
46373 => "0111101110010000",
46374 => "0111101110010000",
46375 => "0111101110010000",
46376 => "0111101110010000",
46377 => "0111101110010000",
46378 => "0111101110010000",
46379 => "0111101110010000",
46380 => "0111101110010000",
46381 => "0111101110010000",
46382 => "0111101110010000",
46383 => "0111101110010000",
46384 => "0111101110010000",
46385 => "0111101110010000",
46386 => "0111101110010000",
46387 => "0111101110010000",
46388 => "0111101110010000",
46389 => "0111101110010000",
46390 => "0111101110010000",
46391 => "0111101110010000",
46392 => "0111101110010000",
46393 => "0111101110010000",
46394 => "0111101110010000",
46395 => "0111101110010000",
46396 => "0111101110010000",
46397 => "0111101110010000",
46398 => "0111101110010000",
46399 => "0111101110010000",
46400 => "0111101110010000",
46401 => "0111101110010000",
46402 => "0111101110010000",
46403 => "0111101110010000",
46404 => "0111101110010000",
46405 => "0111101110010000",
46406 => "0111101110010000",
46407 => "0111101110010000",
46408 => "0111101110010000",
46409 => "0111101110010000",
46410 => "0111101110010000",
46411 => "0111101110010000",
46412 => "0111101110010000",
46413 => "0111101110010000",
46414 => "0111101110010000",
46415 => "0111101110010000",
46416 => "0111101110010000",
46417 => "0111101110010000",
46418 => "0111101110010000",
46419 => "0111101110010000",
46420 => "0111101110010000",
46421 => "0111101110010000",
46422 => "0111101110010000",
46423 => "0111101110010000",
46424 => "0111101110100000",
46425 => "0111101110100000",
46426 => "0111101110100000",
46427 => "0111101110100000",
46428 => "0111101110100000",
46429 => "0111101110100000",
46430 => "0111101110100000",
46431 => "0111101110100000",
46432 => "0111101110100000",
46433 => "0111101110100000",
46434 => "0111101110100000",
46435 => "0111101110100000",
46436 => "0111101110100000",
46437 => "0111101110100000",
46438 => "0111101110100000",
46439 => "0111101110100000",
46440 => "0111101110100000",
46441 => "0111101110100000",
46442 => "0111101110100000",
46443 => "0111101110100000",
46444 => "0111101110100000",
46445 => "0111101110100000",
46446 => "0111101110100000",
46447 => "0111101110100000",
46448 => "0111101110100000",
46449 => "0111101110100000",
46450 => "0111101110100000",
46451 => "0111101110100000",
46452 => "0111101110100000",
46453 => "0111101110100000",
46454 => "0111101110100000",
46455 => "0111101110100000",
46456 => "0111101110100000",
46457 => "0111101110100000",
46458 => "0111101110100000",
46459 => "0111101110100000",
46460 => "0111101110100000",
46461 => "0111101110100000",
46462 => "0111101110100000",
46463 => "0111101110100000",
46464 => "0111101110100000",
46465 => "0111101110100000",
46466 => "0111101110100000",
46467 => "0111101110100000",
46468 => "0111101110100000",
46469 => "0111101110100000",
46470 => "0111101110100000",
46471 => "0111101110100000",
46472 => "0111101110100000",
46473 => "0111101110100000",
46474 => "0111101110100000",
46475 => "0111101110100000",
46476 => "0111101110100000",
46477 => "0111101110100000",
46478 => "0111101110100000",
46479 => "0111101110100000",
46480 => "0111101110100000",
46481 => "0111101110100000",
46482 => "0111101110100000",
46483 => "0111101110100000",
46484 => "0111101110110000",
46485 => "0111101110110000",
46486 => "0111101110110000",
46487 => "0111101110110000",
46488 => "0111101110110000",
46489 => "0111101110110000",
46490 => "0111101110110000",
46491 => "0111101110110000",
46492 => "0111101110110000",
46493 => "0111101110110000",
46494 => "0111101110110000",
46495 => "0111101110110000",
46496 => "0111101110110000",
46497 => "0111101110110000",
46498 => "0111101110110000",
46499 => "0111101110110000",
46500 => "0111101110110000",
46501 => "0111101110110000",
46502 => "0111101110110000",
46503 => "0111101110110000",
46504 => "0111101110110000",
46505 => "0111101110110000",
46506 => "0111101110110000",
46507 => "0111101110110000",
46508 => "0111101110110000",
46509 => "0111101110110000",
46510 => "0111101110110000",
46511 => "0111101110110000",
46512 => "0111101110110000",
46513 => "0111101110110000",
46514 => "0111101110110000",
46515 => "0111101110110000",
46516 => "0111101110110000",
46517 => "0111101110110000",
46518 => "0111101110110000",
46519 => "0111101110110000",
46520 => "0111101110110000",
46521 => "0111101110110000",
46522 => "0111101110110000",
46523 => "0111101110110000",
46524 => "0111101110110000",
46525 => "0111101110110000",
46526 => "0111101110110000",
46527 => "0111101110110000",
46528 => "0111101110110000",
46529 => "0111101110110000",
46530 => "0111101110110000",
46531 => "0111101110110000",
46532 => "0111101110110000",
46533 => "0111101110110000",
46534 => "0111101110110000",
46535 => "0111101110110000",
46536 => "0111101110110000",
46537 => "0111101110110000",
46538 => "0111101110110000",
46539 => "0111101110110000",
46540 => "0111101110110000",
46541 => "0111101110110000",
46542 => "0111101110110000",
46543 => "0111101110110000",
46544 => "0111101110110000",
46545 => "0111101110110000",
46546 => "0111101111000000",
46547 => "0111101111000000",
46548 => "0111101111000000",
46549 => "0111101111000000",
46550 => "0111101111000000",
46551 => "0111101111000000",
46552 => "0111101111000000",
46553 => "0111101111000000",
46554 => "0111101111000000",
46555 => "0111101111000000",
46556 => "0111101111000000",
46557 => "0111101111000000",
46558 => "0111101111000000",
46559 => "0111101111000000",
46560 => "0111101111000000",
46561 => "0111101111000000",
46562 => "0111101111000000",
46563 => "0111101111000000",
46564 => "0111101111000000",
46565 => "0111101111000000",
46566 => "0111101111000000",
46567 => "0111101111000000",
46568 => "0111101111000000",
46569 => "0111101111000000",
46570 => "0111101111000000",
46571 => "0111101111000000",
46572 => "0111101111000000",
46573 => "0111101111000000",
46574 => "0111101111000000",
46575 => "0111101111000000",
46576 => "0111101111000000",
46577 => "0111101111000000",
46578 => "0111101111000000",
46579 => "0111101111000000",
46580 => "0111101111000000",
46581 => "0111101111000000",
46582 => "0111101111000000",
46583 => "0111101111000000",
46584 => "0111101111000000",
46585 => "0111101111000000",
46586 => "0111101111000000",
46587 => "0111101111000000",
46588 => "0111101111000000",
46589 => "0111101111000000",
46590 => "0111101111000000",
46591 => "0111101111000000",
46592 => "0111101111000000",
46593 => "0111101111000000",
46594 => "0111101111000000",
46595 => "0111101111000000",
46596 => "0111101111000000",
46597 => "0111101111000000",
46598 => "0111101111000000",
46599 => "0111101111000000",
46600 => "0111101111000000",
46601 => "0111101111000000",
46602 => "0111101111000000",
46603 => "0111101111000000",
46604 => "0111101111000000",
46605 => "0111101111000000",
46606 => "0111101111000000",
46607 => "0111101111000000",
46608 => "0111101111010000",
46609 => "0111101111010000",
46610 => "0111101111010000",
46611 => "0111101111010000",
46612 => "0111101111010000",
46613 => "0111101111010000",
46614 => "0111101111010000",
46615 => "0111101111010000",
46616 => "0111101111010000",
46617 => "0111101111010000",
46618 => "0111101111010000",
46619 => "0111101111010000",
46620 => "0111101111010000",
46621 => "0111101111010000",
46622 => "0111101111010000",
46623 => "0111101111010000",
46624 => "0111101111010000",
46625 => "0111101111010000",
46626 => "0111101111010000",
46627 => "0111101111010000",
46628 => "0111101111010000",
46629 => "0111101111010000",
46630 => "0111101111010000",
46631 => "0111101111010000",
46632 => "0111101111010000",
46633 => "0111101111010000",
46634 => "0111101111010000",
46635 => "0111101111010000",
46636 => "0111101111010000",
46637 => "0111101111010000",
46638 => "0111101111010000",
46639 => "0111101111010000",
46640 => "0111101111010000",
46641 => "0111101111010000",
46642 => "0111101111010000",
46643 => "0111101111010000",
46644 => "0111101111010000",
46645 => "0111101111010000",
46646 => "0111101111010000",
46647 => "0111101111010000",
46648 => "0111101111010000",
46649 => "0111101111010000",
46650 => "0111101111010000",
46651 => "0111101111010000",
46652 => "0111101111010000",
46653 => "0111101111010000",
46654 => "0111101111010000",
46655 => "0111101111010000",
46656 => "0111101111010000",
46657 => "0111101111010000",
46658 => "0111101111010000",
46659 => "0111101111010000",
46660 => "0111101111010000",
46661 => "0111101111010000",
46662 => "0111101111010000",
46663 => "0111101111010000",
46664 => "0111101111010000",
46665 => "0111101111010000",
46666 => "0111101111010000",
46667 => "0111101111010000",
46668 => "0111101111010000",
46669 => "0111101111010000",
46670 => "0111101111010000",
46671 => "0111101111100000",
46672 => "0111101111100000",
46673 => "0111101111100000",
46674 => "0111101111100000",
46675 => "0111101111100000",
46676 => "0111101111100000",
46677 => "0111101111100000",
46678 => "0111101111100000",
46679 => "0111101111100000",
46680 => "0111101111100000",
46681 => "0111101111100000",
46682 => "0111101111100000",
46683 => "0111101111100000",
46684 => "0111101111100000",
46685 => "0111101111100000",
46686 => "0111101111100000",
46687 => "0111101111100000",
46688 => "0111101111100000",
46689 => "0111101111100000",
46690 => "0111101111100000",
46691 => "0111101111100000",
46692 => "0111101111100000",
46693 => "0111101111100000",
46694 => "0111101111100000",
46695 => "0111101111100000",
46696 => "0111101111100000",
46697 => "0111101111100000",
46698 => "0111101111100000",
46699 => "0111101111100000",
46700 => "0111101111100000",
46701 => "0111101111100000",
46702 => "0111101111100000",
46703 => "0111101111100000",
46704 => "0111101111100000",
46705 => "0111101111100000",
46706 => "0111101111100000",
46707 => "0111101111100000",
46708 => "0111101111100000",
46709 => "0111101111100000",
46710 => "0111101111100000",
46711 => "0111101111100000",
46712 => "0111101111100000",
46713 => "0111101111100000",
46714 => "0111101111100000",
46715 => "0111101111100000",
46716 => "0111101111100000",
46717 => "0111101111100000",
46718 => "0111101111100000",
46719 => "0111101111100000",
46720 => "0111101111100000",
46721 => "0111101111100000",
46722 => "0111101111100000",
46723 => "0111101111100000",
46724 => "0111101111100000",
46725 => "0111101111100000",
46726 => "0111101111100000",
46727 => "0111101111100000",
46728 => "0111101111100000",
46729 => "0111101111100000",
46730 => "0111101111100000",
46731 => "0111101111100000",
46732 => "0111101111100000",
46733 => "0111101111100000",
46734 => "0111101111100000",
46735 => "0111101111110000",
46736 => "0111101111110000",
46737 => "0111101111110000",
46738 => "0111101111110000",
46739 => "0111101111110000",
46740 => "0111101111110000",
46741 => "0111101111110000",
46742 => "0111101111110000",
46743 => "0111101111110000",
46744 => "0111101111110000",
46745 => "0111101111110000",
46746 => "0111101111110000",
46747 => "0111101111110000",
46748 => "0111101111110000",
46749 => "0111101111110000",
46750 => "0111101111110000",
46751 => "0111101111110000",
46752 => "0111101111110000",
46753 => "0111101111110000",
46754 => "0111101111110000",
46755 => "0111101111110000",
46756 => "0111101111110000",
46757 => "0111101111110000",
46758 => "0111101111110000",
46759 => "0111101111110000",
46760 => "0111101111110000",
46761 => "0111101111110000",
46762 => "0111101111110000",
46763 => "0111101111110000",
46764 => "0111101111110000",
46765 => "0111101111110000",
46766 => "0111101111110000",
46767 => "0111101111110000",
46768 => "0111101111110000",
46769 => "0111101111110000",
46770 => "0111101111110000",
46771 => "0111101111110000",
46772 => "0111101111110000",
46773 => "0111101111110000",
46774 => "0111101111110000",
46775 => "0111101111110000",
46776 => "0111101111110000",
46777 => "0111101111110000",
46778 => "0111101111110000",
46779 => "0111101111110000",
46780 => "0111101111110000",
46781 => "0111101111110000",
46782 => "0111101111110000",
46783 => "0111101111110000",
46784 => "0111101111110000",
46785 => "0111101111110000",
46786 => "0111101111110000",
46787 => "0111101111110000",
46788 => "0111101111110000",
46789 => "0111101111110000",
46790 => "0111101111110000",
46791 => "0111101111110000",
46792 => "0111101111110000",
46793 => "0111101111110000",
46794 => "0111101111110000",
46795 => "0111101111110000",
46796 => "0111101111110000",
46797 => "0111101111110000",
46798 => "0111101111110000",
46799 => "0111101111110000",
46800 => "0111110000000000",
46801 => "0111110000000000",
46802 => "0111110000000000",
46803 => "0111110000000000",
46804 => "0111110000000000",
46805 => "0111110000000000",
46806 => "0111110000000000",
46807 => "0111110000000000",
46808 => "0111110000000000",
46809 => "0111110000000000",
46810 => "0111110000000000",
46811 => "0111110000000000",
46812 => "0111110000000000",
46813 => "0111110000000000",
46814 => "0111110000000000",
46815 => "0111110000000000",
46816 => "0111110000000000",
46817 => "0111110000000000",
46818 => "0111110000000000",
46819 => "0111110000000000",
46820 => "0111110000000000",
46821 => "0111110000000000",
46822 => "0111110000000000",
46823 => "0111110000000000",
46824 => "0111110000000000",
46825 => "0111110000000000",
46826 => "0111110000000000",
46827 => "0111110000000000",
46828 => "0111110000000000",
46829 => "0111110000000000",
46830 => "0111110000000000",
46831 => "0111110000000000",
46832 => "0111110000000000",
46833 => "0111110000000000",
46834 => "0111110000000000",
46835 => "0111110000000000",
46836 => "0111110000000000",
46837 => "0111110000000000",
46838 => "0111110000000000",
46839 => "0111110000000000",
46840 => "0111110000000000",
46841 => "0111110000000000",
46842 => "0111110000000000",
46843 => "0111110000000000",
46844 => "0111110000000000",
46845 => "0111110000000000",
46846 => "0111110000000000",
46847 => "0111110000000000",
46848 => "0111110000000000",
46849 => "0111110000000000",
46850 => "0111110000000000",
46851 => "0111110000000000",
46852 => "0111110000000000",
46853 => "0111110000000000",
46854 => "0111110000000000",
46855 => "0111110000000000",
46856 => "0111110000000000",
46857 => "0111110000000000",
46858 => "0111110000000000",
46859 => "0111110000000000",
46860 => "0111110000000000",
46861 => "0111110000000000",
46862 => "0111110000000000",
46863 => "0111110000000000",
46864 => "0111110000000000",
46865 => "0111110000000000",
46866 => "0111110000000000",
46867 => "0111110000010000",
46868 => "0111110000010000",
46869 => "0111110000010000",
46870 => "0111110000010000",
46871 => "0111110000010000",
46872 => "0111110000010000",
46873 => "0111110000010000",
46874 => "0111110000010000",
46875 => "0111110000010000",
46876 => "0111110000010000",
46877 => "0111110000010000",
46878 => "0111110000010000",
46879 => "0111110000010000",
46880 => "0111110000010000",
46881 => "0111110000010000",
46882 => "0111110000010000",
46883 => "0111110000010000",
46884 => "0111110000010000",
46885 => "0111110000010000",
46886 => "0111110000010000",
46887 => "0111110000010000",
46888 => "0111110000010000",
46889 => "0111110000010000",
46890 => "0111110000010000",
46891 => "0111110000010000",
46892 => "0111110000010000",
46893 => "0111110000010000",
46894 => "0111110000010000",
46895 => "0111110000010000",
46896 => "0111110000010000",
46897 => "0111110000010000",
46898 => "0111110000010000",
46899 => "0111110000010000",
46900 => "0111110000010000",
46901 => "0111110000010000",
46902 => "0111110000010000",
46903 => "0111110000010000",
46904 => "0111110000010000",
46905 => "0111110000010000",
46906 => "0111110000010000",
46907 => "0111110000010000",
46908 => "0111110000010000",
46909 => "0111110000010000",
46910 => "0111110000010000",
46911 => "0111110000010000",
46912 => "0111110000010000",
46913 => "0111110000010000",
46914 => "0111110000010000",
46915 => "0111110000010000",
46916 => "0111110000010000",
46917 => "0111110000010000",
46918 => "0111110000010000",
46919 => "0111110000010000",
46920 => "0111110000010000",
46921 => "0111110000010000",
46922 => "0111110000010000",
46923 => "0111110000010000",
46924 => "0111110000010000",
46925 => "0111110000010000",
46926 => "0111110000010000",
46927 => "0111110000010000",
46928 => "0111110000010000",
46929 => "0111110000010000",
46930 => "0111110000010000",
46931 => "0111110000010000",
46932 => "0111110000010000",
46933 => "0111110000010000",
46934 => "0111110000100000",
46935 => "0111110000100000",
46936 => "0111110000100000",
46937 => "0111110000100000",
46938 => "0111110000100000",
46939 => "0111110000100000",
46940 => "0111110000100000",
46941 => "0111110000100000",
46942 => "0111110000100000",
46943 => "0111110000100000",
46944 => "0111110000100000",
46945 => "0111110000100000",
46946 => "0111110000100000",
46947 => "0111110000100000",
46948 => "0111110000100000",
46949 => "0111110000100000",
46950 => "0111110000100000",
46951 => "0111110000100000",
46952 => "0111110000100000",
46953 => "0111110000100000",
46954 => "0111110000100000",
46955 => "0111110000100000",
46956 => "0111110000100000",
46957 => "0111110000100000",
46958 => "0111110000100000",
46959 => "0111110000100000",
46960 => "0111110000100000",
46961 => "0111110000100000",
46962 => "0111110000100000",
46963 => "0111110000100000",
46964 => "0111110000100000",
46965 => "0111110000100000",
46966 => "0111110000100000",
46967 => "0111110000100000",
46968 => "0111110000100000",
46969 => "0111110000100000",
46970 => "0111110000100000",
46971 => "0111110000100000",
46972 => "0111110000100000",
46973 => "0111110000100000",
46974 => "0111110000100000",
46975 => "0111110000100000",
46976 => "0111110000100000",
46977 => "0111110000100000",
46978 => "0111110000100000",
46979 => "0111110000100000",
46980 => "0111110000100000",
46981 => "0111110000100000",
46982 => "0111110000100000",
46983 => "0111110000100000",
46984 => "0111110000100000",
46985 => "0111110000100000",
46986 => "0111110000100000",
46987 => "0111110000100000",
46988 => "0111110000100000",
46989 => "0111110000100000",
46990 => "0111110000100000",
46991 => "0111110000100000",
46992 => "0111110000100000",
46993 => "0111110000100000",
46994 => "0111110000100000",
46995 => "0111110000100000",
46996 => "0111110000100000",
46997 => "0111110000100000",
46998 => "0111110000100000",
46999 => "0111110000100000",
47000 => "0111110000100000",
47001 => "0111110000100000",
47002 => "0111110000110000",
47003 => "0111110000110000",
47004 => "0111110000110000",
47005 => "0111110000110000",
47006 => "0111110000110000",
47007 => "0111110000110000",
47008 => "0111110000110000",
47009 => "0111110000110000",
47010 => "0111110000110000",
47011 => "0111110000110000",
47012 => "0111110000110000",
47013 => "0111110000110000",
47014 => "0111110000110000",
47015 => "0111110000110000",
47016 => "0111110000110000",
47017 => "0111110000110000",
47018 => "0111110000110000",
47019 => "0111110000110000",
47020 => "0111110000110000",
47021 => "0111110000110000",
47022 => "0111110000110000",
47023 => "0111110000110000",
47024 => "0111110000110000",
47025 => "0111110000110000",
47026 => "0111110000110000",
47027 => "0111110000110000",
47028 => "0111110000110000",
47029 => "0111110000110000",
47030 => "0111110000110000",
47031 => "0111110000110000",
47032 => "0111110000110000",
47033 => "0111110000110000",
47034 => "0111110000110000",
47035 => "0111110000110000",
47036 => "0111110000110000",
47037 => "0111110000110000",
47038 => "0111110000110000",
47039 => "0111110000110000",
47040 => "0111110000110000",
47041 => "0111110000110000",
47042 => "0111110000110000",
47043 => "0111110000110000",
47044 => "0111110000110000",
47045 => "0111110000110000",
47046 => "0111110000110000",
47047 => "0111110000110000",
47048 => "0111110000110000",
47049 => "0111110000110000",
47050 => "0111110000110000",
47051 => "0111110000110000",
47052 => "0111110000110000",
47053 => "0111110000110000",
47054 => "0111110000110000",
47055 => "0111110000110000",
47056 => "0111110000110000",
47057 => "0111110000110000",
47058 => "0111110000110000",
47059 => "0111110000110000",
47060 => "0111110000110000",
47061 => "0111110000110000",
47062 => "0111110000110000",
47063 => "0111110000110000",
47064 => "0111110000110000",
47065 => "0111110000110000",
47066 => "0111110000110000",
47067 => "0111110000110000",
47068 => "0111110000110000",
47069 => "0111110000110000",
47070 => "0111110000110000",
47071 => "0111110001000000",
47072 => "0111110001000000",
47073 => "0111110001000000",
47074 => "0111110001000000",
47075 => "0111110001000000",
47076 => "0111110001000000",
47077 => "0111110001000000",
47078 => "0111110001000000",
47079 => "0111110001000000",
47080 => "0111110001000000",
47081 => "0111110001000000",
47082 => "0111110001000000",
47083 => "0111110001000000",
47084 => "0111110001000000",
47085 => "0111110001000000",
47086 => "0111110001000000",
47087 => "0111110001000000",
47088 => "0111110001000000",
47089 => "0111110001000000",
47090 => "0111110001000000",
47091 => "0111110001000000",
47092 => "0111110001000000",
47093 => "0111110001000000",
47094 => "0111110001000000",
47095 => "0111110001000000",
47096 => "0111110001000000",
47097 => "0111110001000000",
47098 => "0111110001000000",
47099 => "0111110001000000",
47100 => "0111110001000000",
47101 => "0111110001000000",
47102 => "0111110001000000",
47103 => "0111110001000000",
47104 => "0111110001000000",
47105 => "0111110001000000",
47106 => "0111110001000000",
47107 => "0111110001000000",
47108 => "0111110001000000",
47109 => "0111110001000000",
47110 => "0111110001000000",
47111 => "0111110001000000",
47112 => "0111110001000000",
47113 => "0111110001000000",
47114 => "0111110001000000",
47115 => "0111110001000000",
47116 => "0111110001000000",
47117 => "0111110001000000",
47118 => "0111110001000000",
47119 => "0111110001000000",
47120 => "0111110001000000",
47121 => "0111110001000000",
47122 => "0111110001000000",
47123 => "0111110001000000",
47124 => "0111110001000000",
47125 => "0111110001000000",
47126 => "0111110001000000",
47127 => "0111110001000000",
47128 => "0111110001000000",
47129 => "0111110001000000",
47130 => "0111110001000000",
47131 => "0111110001000000",
47132 => "0111110001000000",
47133 => "0111110001000000",
47134 => "0111110001000000",
47135 => "0111110001000000",
47136 => "0111110001000000",
47137 => "0111110001000000",
47138 => "0111110001000000",
47139 => "0111110001000000",
47140 => "0111110001000000",
47141 => "0111110001010000",
47142 => "0111110001010000",
47143 => "0111110001010000",
47144 => "0111110001010000",
47145 => "0111110001010000",
47146 => "0111110001010000",
47147 => "0111110001010000",
47148 => "0111110001010000",
47149 => "0111110001010000",
47150 => "0111110001010000",
47151 => "0111110001010000",
47152 => "0111110001010000",
47153 => "0111110001010000",
47154 => "0111110001010000",
47155 => "0111110001010000",
47156 => "0111110001010000",
47157 => "0111110001010000",
47158 => "0111110001010000",
47159 => "0111110001010000",
47160 => "0111110001010000",
47161 => "0111110001010000",
47162 => "0111110001010000",
47163 => "0111110001010000",
47164 => "0111110001010000",
47165 => "0111110001010000",
47166 => "0111110001010000",
47167 => "0111110001010000",
47168 => "0111110001010000",
47169 => "0111110001010000",
47170 => "0111110001010000",
47171 => "0111110001010000",
47172 => "0111110001010000",
47173 => "0111110001010000",
47174 => "0111110001010000",
47175 => "0111110001010000",
47176 => "0111110001010000",
47177 => "0111110001010000",
47178 => "0111110001010000",
47179 => "0111110001010000",
47180 => "0111110001010000",
47181 => "0111110001010000",
47182 => "0111110001010000",
47183 => "0111110001010000",
47184 => "0111110001010000",
47185 => "0111110001010000",
47186 => "0111110001010000",
47187 => "0111110001010000",
47188 => "0111110001010000",
47189 => "0111110001010000",
47190 => "0111110001010000",
47191 => "0111110001010000",
47192 => "0111110001010000",
47193 => "0111110001010000",
47194 => "0111110001010000",
47195 => "0111110001010000",
47196 => "0111110001010000",
47197 => "0111110001010000",
47198 => "0111110001010000",
47199 => "0111110001010000",
47200 => "0111110001010000",
47201 => "0111110001010000",
47202 => "0111110001010000",
47203 => "0111110001010000",
47204 => "0111110001010000",
47205 => "0111110001010000",
47206 => "0111110001010000",
47207 => "0111110001010000",
47208 => "0111110001010000",
47209 => "0111110001010000",
47210 => "0111110001010000",
47211 => "0111110001010000",
47212 => "0111110001010000",
47213 => "0111110001100000",
47214 => "0111110001100000",
47215 => "0111110001100000",
47216 => "0111110001100000",
47217 => "0111110001100000",
47218 => "0111110001100000",
47219 => "0111110001100000",
47220 => "0111110001100000",
47221 => "0111110001100000",
47222 => "0111110001100000",
47223 => "0111110001100000",
47224 => "0111110001100000",
47225 => "0111110001100000",
47226 => "0111110001100000",
47227 => "0111110001100000",
47228 => "0111110001100000",
47229 => "0111110001100000",
47230 => "0111110001100000",
47231 => "0111110001100000",
47232 => "0111110001100000",
47233 => "0111110001100000",
47234 => "0111110001100000",
47235 => "0111110001100000",
47236 => "0111110001100000",
47237 => "0111110001100000",
47238 => "0111110001100000",
47239 => "0111110001100000",
47240 => "0111110001100000",
47241 => "0111110001100000",
47242 => "0111110001100000",
47243 => "0111110001100000",
47244 => "0111110001100000",
47245 => "0111110001100000",
47246 => "0111110001100000",
47247 => "0111110001100000",
47248 => "0111110001100000",
47249 => "0111110001100000",
47250 => "0111110001100000",
47251 => "0111110001100000",
47252 => "0111110001100000",
47253 => "0111110001100000",
47254 => "0111110001100000",
47255 => "0111110001100000",
47256 => "0111110001100000",
47257 => "0111110001100000",
47258 => "0111110001100000",
47259 => "0111110001100000",
47260 => "0111110001100000",
47261 => "0111110001100000",
47262 => "0111110001100000",
47263 => "0111110001100000",
47264 => "0111110001100000",
47265 => "0111110001100000",
47266 => "0111110001100000",
47267 => "0111110001100000",
47268 => "0111110001100000",
47269 => "0111110001100000",
47270 => "0111110001100000",
47271 => "0111110001100000",
47272 => "0111110001100000",
47273 => "0111110001100000",
47274 => "0111110001100000",
47275 => "0111110001100000",
47276 => "0111110001100000",
47277 => "0111110001100000",
47278 => "0111110001100000",
47279 => "0111110001100000",
47280 => "0111110001100000",
47281 => "0111110001100000",
47282 => "0111110001100000",
47283 => "0111110001100000",
47284 => "0111110001100000",
47285 => "0111110001110000",
47286 => "0111110001110000",
47287 => "0111110001110000",
47288 => "0111110001110000",
47289 => "0111110001110000",
47290 => "0111110001110000",
47291 => "0111110001110000",
47292 => "0111110001110000",
47293 => "0111110001110000",
47294 => "0111110001110000",
47295 => "0111110001110000",
47296 => "0111110001110000",
47297 => "0111110001110000",
47298 => "0111110001110000",
47299 => "0111110001110000",
47300 => "0111110001110000",
47301 => "0111110001110000",
47302 => "0111110001110000",
47303 => "0111110001110000",
47304 => "0111110001110000",
47305 => "0111110001110000",
47306 => "0111110001110000",
47307 => "0111110001110000",
47308 => "0111110001110000",
47309 => "0111110001110000",
47310 => "0111110001110000",
47311 => "0111110001110000",
47312 => "0111110001110000",
47313 => "0111110001110000",
47314 => "0111110001110000",
47315 => "0111110001110000",
47316 => "0111110001110000",
47317 => "0111110001110000",
47318 => "0111110001110000",
47319 => "0111110001110000",
47320 => "0111110001110000",
47321 => "0111110001110000",
47322 => "0111110001110000",
47323 => "0111110001110000",
47324 => "0111110001110000",
47325 => "0111110001110000",
47326 => "0111110001110000",
47327 => "0111110001110000",
47328 => "0111110001110000",
47329 => "0111110001110000",
47330 => "0111110001110000",
47331 => "0111110001110000",
47332 => "0111110001110000",
47333 => "0111110001110000",
47334 => "0111110001110000",
47335 => "0111110001110000",
47336 => "0111110001110000",
47337 => "0111110001110000",
47338 => "0111110001110000",
47339 => "0111110001110000",
47340 => "0111110001110000",
47341 => "0111110001110000",
47342 => "0111110001110000",
47343 => "0111110001110000",
47344 => "0111110001110000",
47345 => "0111110001110000",
47346 => "0111110001110000",
47347 => "0111110001110000",
47348 => "0111110001110000",
47349 => "0111110001110000",
47350 => "0111110001110000",
47351 => "0111110001110000",
47352 => "0111110001110000",
47353 => "0111110001110000",
47354 => "0111110001110000",
47355 => "0111110001110000",
47356 => "0111110001110000",
47357 => "0111110001110000",
47358 => "0111110001110000",
47359 => "0111110010000000",
47360 => "0111110010000000",
47361 => "0111110010000000",
47362 => "0111110010000000",
47363 => "0111110010000000",
47364 => "0111110010000000",
47365 => "0111110010000000",
47366 => "0111110010000000",
47367 => "0111110010000000",
47368 => "0111110010000000",
47369 => "0111110010000000",
47370 => "0111110010000000",
47371 => "0111110010000000",
47372 => "0111110010000000",
47373 => "0111110010000000",
47374 => "0111110010000000",
47375 => "0111110010000000",
47376 => "0111110010000000",
47377 => "0111110010000000",
47378 => "0111110010000000",
47379 => "0111110010000000",
47380 => "0111110010000000",
47381 => "0111110010000000",
47382 => "0111110010000000",
47383 => "0111110010000000",
47384 => "0111110010000000",
47385 => "0111110010000000",
47386 => "0111110010000000",
47387 => "0111110010000000",
47388 => "0111110010000000",
47389 => "0111110010000000",
47390 => "0111110010000000",
47391 => "0111110010000000",
47392 => "0111110010000000",
47393 => "0111110010000000",
47394 => "0111110010000000",
47395 => "0111110010000000",
47396 => "0111110010000000",
47397 => "0111110010000000",
47398 => "0111110010000000",
47399 => "0111110010000000",
47400 => "0111110010000000",
47401 => "0111110010000000",
47402 => "0111110010000000",
47403 => "0111110010000000",
47404 => "0111110010000000",
47405 => "0111110010000000",
47406 => "0111110010000000",
47407 => "0111110010000000",
47408 => "0111110010000000",
47409 => "0111110010000000",
47410 => "0111110010000000",
47411 => "0111110010000000",
47412 => "0111110010000000",
47413 => "0111110010000000",
47414 => "0111110010000000",
47415 => "0111110010000000",
47416 => "0111110010000000",
47417 => "0111110010000000",
47418 => "0111110010000000",
47419 => "0111110010000000",
47420 => "0111110010000000",
47421 => "0111110010000000",
47422 => "0111110010000000",
47423 => "0111110010000000",
47424 => "0111110010000000",
47425 => "0111110010000000",
47426 => "0111110010000000",
47427 => "0111110010000000",
47428 => "0111110010000000",
47429 => "0111110010000000",
47430 => "0111110010000000",
47431 => "0111110010000000",
47432 => "0111110010000000",
47433 => "0111110010000000",
47434 => "0111110010000000",
47435 => "0111110010010000",
47436 => "0111110010010000",
47437 => "0111110010010000",
47438 => "0111110010010000",
47439 => "0111110010010000",
47440 => "0111110010010000",
47441 => "0111110010010000",
47442 => "0111110010010000",
47443 => "0111110010010000",
47444 => "0111110010010000",
47445 => "0111110010010000",
47446 => "0111110010010000",
47447 => "0111110010010000",
47448 => "0111110010010000",
47449 => "0111110010010000",
47450 => "0111110010010000",
47451 => "0111110010010000",
47452 => "0111110010010000",
47453 => "0111110010010000",
47454 => "0111110010010000",
47455 => "0111110010010000",
47456 => "0111110010010000",
47457 => "0111110010010000",
47458 => "0111110010010000",
47459 => "0111110010010000",
47460 => "0111110010010000",
47461 => "0111110010010000",
47462 => "0111110010010000",
47463 => "0111110010010000",
47464 => "0111110010010000",
47465 => "0111110010010000",
47466 => "0111110010010000",
47467 => "0111110010010000",
47468 => "0111110010010000",
47469 => "0111110010010000",
47470 => "0111110010010000",
47471 => "0111110010010000",
47472 => "0111110010010000",
47473 => "0111110010010000",
47474 => "0111110010010000",
47475 => "0111110010010000",
47476 => "0111110010010000",
47477 => "0111110010010000",
47478 => "0111110010010000",
47479 => "0111110010010000",
47480 => "0111110010010000",
47481 => "0111110010010000",
47482 => "0111110010010000",
47483 => "0111110010010000",
47484 => "0111110010010000",
47485 => "0111110010010000",
47486 => "0111110010010000",
47487 => "0111110010010000",
47488 => "0111110010010000",
47489 => "0111110010010000",
47490 => "0111110010010000",
47491 => "0111110010010000",
47492 => "0111110010010000",
47493 => "0111110010010000",
47494 => "0111110010010000",
47495 => "0111110010010000",
47496 => "0111110010010000",
47497 => "0111110010010000",
47498 => "0111110010010000",
47499 => "0111110010010000",
47500 => "0111110010010000",
47501 => "0111110010010000",
47502 => "0111110010010000",
47503 => "0111110010010000",
47504 => "0111110010010000",
47505 => "0111110010010000",
47506 => "0111110010010000",
47507 => "0111110010010000",
47508 => "0111110010010000",
47509 => "0111110010010000",
47510 => "0111110010010000",
47511 => "0111110010100000",
47512 => "0111110010100000",
47513 => "0111110010100000",
47514 => "0111110010100000",
47515 => "0111110010100000",
47516 => "0111110010100000",
47517 => "0111110010100000",
47518 => "0111110010100000",
47519 => "0111110010100000",
47520 => "0111110010100000",
47521 => "0111110010100000",
47522 => "0111110010100000",
47523 => "0111110010100000",
47524 => "0111110010100000",
47525 => "0111110010100000",
47526 => "0111110010100000",
47527 => "0111110010100000",
47528 => "0111110010100000",
47529 => "0111110010100000",
47530 => "0111110010100000",
47531 => "0111110010100000",
47532 => "0111110010100000",
47533 => "0111110010100000",
47534 => "0111110010100000",
47535 => "0111110010100000",
47536 => "0111110010100000",
47537 => "0111110010100000",
47538 => "0111110010100000",
47539 => "0111110010100000",
47540 => "0111110010100000",
47541 => "0111110010100000",
47542 => "0111110010100000",
47543 => "0111110010100000",
47544 => "0111110010100000",
47545 => "0111110010100000",
47546 => "0111110010100000",
47547 => "0111110010100000",
47548 => "0111110010100000",
47549 => "0111110010100000",
47550 => "0111110010100000",
47551 => "0111110010100000",
47552 => "0111110010100000",
47553 => "0111110010100000",
47554 => "0111110010100000",
47555 => "0111110010100000",
47556 => "0111110010100000",
47557 => "0111110010100000",
47558 => "0111110010100000",
47559 => "0111110010100000",
47560 => "0111110010100000",
47561 => "0111110010100000",
47562 => "0111110010100000",
47563 => "0111110010100000",
47564 => "0111110010100000",
47565 => "0111110010100000",
47566 => "0111110010100000",
47567 => "0111110010100000",
47568 => "0111110010100000",
47569 => "0111110010100000",
47570 => "0111110010100000",
47571 => "0111110010100000",
47572 => "0111110010100000",
47573 => "0111110010100000",
47574 => "0111110010100000",
47575 => "0111110010100000",
47576 => "0111110010100000",
47577 => "0111110010100000",
47578 => "0111110010100000",
47579 => "0111110010100000",
47580 => "0111110010100000",
47581 => "0111110010100000",
47582 => "0111110010100000",
47583 => "0111110010100000",
47584 => "0111110010100000",
47585 => "0111110010100000",
47586 => "0111110010100000",
47587 => "0111110010100000",
47588 => "0111110010100000",
47589 => "0111110010110000",
47590 => "0111110010110000",
47591 => "0111110010110000",
47592 => "0111110010110000",
47593 => "0111110010110000",
47594 => "0111110010110000",
47595 => "0111110010110000",
47596 => "0111110010110000",
47597 => "0111110010110000",
47598 => "0111110010110000",
47599 => "0111110010110000",
47600 => "0111110010110000",
47601 => "0111110010110000",
47602 => "0111110010110000",
47603 => "0111110010110000",
47604 => "0111110010110000",
47605 => "0111110010110000",
47606 => "0111110010110000",
47607 => "0111110010110000",
47608 => "0111110010110000",
47609 => "0111110010110000",
47610 => "0111110010110000",
47611 => "0111110010110000",
47612 => "0111110010110000",
47613 => "0111110010110000",
47614 => "0111110010110000",
47615 => "0111110010110000",
47616 => "0111110010110000",
47617 => "0111110010110000",
47618 => "0111110010110000",
47619 => "0111110010110000",
47620 => "0111110010110000",
47621 => "0111110010110000",
47622 => "0111110010110000",
47623 => "0111110010110000",
47624 => "0111110010110000",
47625 => "0111110010110000",
47626 => "0111110010110000",
47627 => "0111110010110000",
47628 => "0111110010110000",
47629 => "0111110010110000",
47630 => "0111110010110000",
47631 => "0111110010110000",
47632 => "0111110010110000",
47633 => "0111110010110000",
47634 => "0111110010110000",
47635 => "0111110010110000",
47636 => "0111110010110000",
47637 => "0111110010110000",
47638 => "0111110010110000",
47639 => "0111110010110000",
47640 => "0111110010110000",
47641 => "0111110010110000",
47642 => "0111110010110000",
47643 => "0111110010110000",
47644 => "0111110010110000",
47645 => "0111110010110000",
47646 => "0111110010110000",
47647 => "0111110010110000",
47648 => "0111110010110000",
47649 => "0111110010110000",
47650 => "0111110010110000",
47651 => "0111110010110000",
47652 => "0111110010110000",
47653 => "0111110010110000",
47654 => "0111110010110000",
47655 => "0111110010110000",
47656 => "0111110010110000",
47657 => "0111110010110000",
47658 => "0111110010110000",
47659 => "0111110010110000",
47660 => "0111110010110000",
47661 => "0111110010110000",
47662 => "0111110010110000",
47663 => "0111110010110000",
47664 => "0111110010110000",
47665 => "0111110010110000",
47666 => "0111110010110000",
47667 => "0111110010110000",
47668 => "0111110011000000",
47669 => "0111110011000000",
47670 => "0111110011000000",
47671 => "0111110011000000",
47672 => "0111110011000000",
47673 => "0111110011000000",
47674 => "0111110011000000",
47675 => "0111110011000000",
47676 => "0111110011000000",
47677 => "0111110011000000",
47678 => "0111110011000000",
47679 => "0111110011000000",
47680 => "0111110011000000",
47681 => "0111110011000000",
47682 => "0111110011000000",
47683 => "0111110011000000",
47684 => "0111110011000000",
47685 => "0111110011000000",
47686 => "0111110011000000",
47687 => "0111110011000000",
47688 => "0111110011000000",
47689 => "0111110011000000",
47690 => "0111110011000000",
47691 => "0111110011000000",
47692 => "0111110011000000",
47693 => "0111110011000000",
47694 => "0111110011000000",
47695 => "0111110011000000",
47696 => "0111110011000000",
47697 => "0111110011000000",
47698 => "0111110011000000",
47699 => "0111110011000000",
47700 => "0111110011000000",
47701 => "0111110011000000",
47702 => "0111110011000000",
47703 => "0111110011000000",
47704 => "0111110011000000",
47705 => "0111110011000000",
47706 => "0111110011000000",
47707 => "0111110011000000",
47708 => "0111110011000000",
47709 => "0111110011000000",
47710 => "0111110011000000",
47711 => "0111110011000000",
47712 => "0111110011000000",
47713 => "0111110011000000",
47714 => "0111110011000000",
47715 => "0111110011000000",
47716 => "0111110011000000",
47717 => "0111110011000000",
47718 => "0111110011000000",
47719 => "0111110011000000",
47720 => "0111110011000000",
47721 => "0111110011000000",
47722 => "0111110011000000",
47723 => "0111110011000000",
47724 => "0111110011000000",
47725 => "0111110011000000",
47726 => "0111110011000000",
47727 => "0111110011000000",
47728 => "0111110011000000",
47729 => "0111110011000000",
47730 => "0111110011000000",
47731 => "0111110011000000",
47732 => "0111110011000000",
47733 => "0111110011000000",
47734 => "0111110011000000",
47735 => "0111110011000000",
47736 => "0111110011000000",
47737 => "0111110011000000",
47738 => "0111110011000000",
47739 => "0111110011000000",
47740 => "0111110011000000",
47741 => "0111110011000000",
47742 => "0111110011000000",
47743 => "0111110011000000",
47744 => "0111110011000000",
47745 => "0111110011000000",
47746 => "0111110011000000",
47747 => "0111110011000000",
47748 => "0111110011000000",
47749 => "0111110011010000",
47750 => "0111110011010000",
47751 => "0111110011010000",
47752 => "0111110011010000",
47753 => "0111110011010000",
47754 => "0111110011010000",
47755 => "0111110011010000",
47756 => "0111110011010000",
47757 => "0111110011010000",
47758 => "0111110011010000",
47759 => "0111110011010000",
47760 => "0111110011010000",
47761 => "0111110011010000",
47762 => "0111110011010000",
47763 => "0111110011010000",
47764 => "0111110011010000",
47765 => "0111110011010000",
47766 => "0111110011010000",
47767 => "0111110011010000",
47768 => "0111110011010000",
47769 => "0111110011010000",
47770 => "0111110011010000",
47771 => "0111110011010000",
47772 => "0111110011010000",
47773 => "0111110011010000",
47774 => "0111110011010000",
47775 => "0111110011010000",
47776 => "0111110011010000",
47777 => "0111110011010000",
47778 => "0111110011010000",
47779 => "0111110011010000",
47780 => "0111110011010000",
47781 => "0111110011010000",
47782 => "0111110011010000",
47783 => "0111110011010000",
47784 => "0111110011010000",
47785 => "0111110011010000",
47786 => "0111110011010000",
47787 => "0111110011010000",
47788 => "0111110011010000",
47789 => "0111110011010000",
47790 => "0111110011010000",
47791 => "0111110011010000",
47792 => "0111110011010000",
47793 => "0111110011010000",
47794 => "0111110011010000",
47795 => "0111110011010000",
47796 => "0111110011010000",
47797 => "0111110011010000",
47798 => "0111110011010000",
47799 => "0111110011010000",
47800 => "0111110011010000",
47801 => "0111110011010000",
47802 => "0111110011010000",
47803 => "0111110011010000",
47804 => "0111110011010000",
47805 => "0111110011010000",
47806 => "0111110011010000",
47807 => "0111110011010000",
47808 => "0111110011010000",
47809 => "0111110011010000",
47810 => "0111110011010000",
47811 => "0111110011010000",
47812 => "0111110011010000",
47813 => "0111110011010000",
47814 => "0111110011010000",
47815 => "0111110011010000",
47816 => "0111110011010000",
47817 => "0111110011010000",
47818 => "0111110011010000",
47819 => "0111110011010000",
47820 => "0111110011010000",
47821 => "0111110011010000",
47822 => "0111110011010000",
47823 => "0111110011010000",
47824 => "0111110011010000",
47825 => "0111110011010000",
47826 => "0111110011010000",
47827 => "0111110011010000",
47828 => "0111110011010000",
47829 => "0111110011010000",
47830 => "0111110011010000",
47831 => "0111110011010000",
47832 => "0111110011100000",
47833 => "0111110011100000",
47834 => "0111110011100000",
47835 => "0111110011100000",
47836 => "0111110011100000",
47837 => "0111110011100000",
47838 => "0111110011100000",
47839 => "0111110011100000",
47840 => "0111110011100000",
47841 => "0111110011100000",
47842 => "0111110011100000",
47843 => "0111110011100000",
47844 => "0111110011100000",
47845 => "0111110011100000",
47846 => "0111110011100000",
47847 => "0111110011100000",
47848 => "0111110011100000",
47849 => "0111110011100000",
47850 => "0111110011100000",
47851 => "0111110011100000",
47852 => "0111110011100000",
47853 => "0111110011100000",
47854 => "0111110011100000",
47855 => "0111110011100000",
47856 => "0111110011100000",
47857 => "0111110011100000",
47858 => "0111110011100000",
47859 => "0111110011100000",
47860 => "0111110011100000",
47861 => "0111110011100000",
47862 => "0111110011100000",
47863 => "0111110011100000",
47864 => "0111110011100000",
47865 => "0111110011100000",
47866 => "0111110011100000",
47867 => "0111110011100000",
47868 => "0111110011100000",
47869 => "0111110011100000",
47870 => "0111110011100000",
47871 => "0111110011100000",
47872 => "0111110011100000",
47873 => "0111110011100000",
47874 => "0111110011100000",
47875 => "0111110011100000",
47876 => "0111110011100000",
47877 => "0111110011100000",
47878 => "0111110011100000",
47879 => "0111110011100000",
47880 => "0111110011100000",
47881 => "0111110011100000",
47882 => "0111110011100000",
47883 => "0111110011100000",
47884 => "0111110011100000",
47885 => "0111110011100000",
47886 => "0111110011100000",
47887 => "0111110011100000",
47888 => "0111110011100000",
47889 => "0111110011100000",
47890 => "0111110011100000",
47891 => "0111110011100000",
47892 => "0111110011100000",
47893 => "0111110011100000",
47894 => "0111110011100000",
47895 => "0111110011100000",
47896 => "0111110011100000",
47897 => "0111110011100000",
47898 => "0111110011100000",
47899 => "0111110011100000",
47900 => "0111110011100000",
47901 => "0111110011100000",
47902 => "0111110011100000",
47903 => "0111110011100000",
47904 => "0111110011100000",
47905 => "0111110011100000",
47906 => "0111110011100000",
47907 => "0111110011100000",
47908 => "0111110011100000",
47909 => "0111110011100000",
47910 => "0111110011100000",
47911 => "0111110011100000",
47912 => "0111110011100000",
47913 => "0111110011100000",
47914 => "0111110011100000",
47915 => "0111110011100000",
47916 => "0111110011110000",
47917 => "0111110011110000",
47918 => "0111110011110000",
47919 => "0111110011110000",
47920 => "0111110011110000",
47921 => "0111110011110000",
47922 => "0111110011110000",
47923 => "0111110011110000",
47924 => "0111110011110000",
47925 => "0111110011110000",
47926 => "0111110011110000",
47927 => "0111110011110000",
47928 => "0111110011110000",
47929 => "0111110011110000",
47930 => "0111110011110000",
47931 => "0111110011110000",
47932 => "0111110011110000",
47933 => "0111110011110000",
47934 => "0111110011110000",
47935 => "0111110011110000",
47936 => "0111110011110000",
47937 => "0111110011110000",
47938 => "0111110011110000",
47939 => "0111110011110000",
47940 => "0111110011110000",
47941 => "0111110011110000",
47942 => "0111110011110000",
47943 => "0111110011110000",
47944 => "0111110011110000",
47945 => "0111110011110000",
47946 => "0111110011110000",
47947 => "0111110011110000",
47948 => "0111110011110000",
47949 => "0111110011110000",
47950 => "0111110011110000",
47951 => "0111110011110000",
47952 => "0111110011110000",
47953 => "0111110011110000",
47954 => "0111110011110000",
47955 => "0111110011110000",
47956 => "0111110011110000",
47957 => "0111110011110000",
47958 => "0111110011110000",
47959 => "0111110011110000",
47960 => "0111110011110000",
47961 => "0111110011110000",
47962 => "0111110011110000",
47963 => "0111110011110000",
47964 => "0111110011110000",
47965 => "0111110011110000",
47966 => "0111110011110000",
47967 => "0111110011110000",
47968 => "0111110011110000",
47969 => "0111110011110000",
47970 => "0111110011110000",
47971 => "0111110011110000",
47972 => "0111110011110000",
47973 => "0111110011110000",
47974 => "0111110011110000",
47975 => "0111110011110000",
47976 => "0111110011110000",
47977 => "0111110011110000",
47978 => "0111110011110000",
47979 => "0111110011110000",
47980 => "0111110011110000",
47981 => "0111110011110000",
47982 => "0111110011110000",
47983 => "0111110011110000",
47984 => "0111110011110000",
47985 => "0111110011110000",
47986 => "0111110011110000",
47987 => "0111110011110000",
47988 => "0111110011110000",
47989 => "0111110011110000",
47990 => "0111110011110000",
47991 => "0111110011110000",
47992 => "0111110011110000",
47993 => "0111110011110000",
47994 => "0111110011110000",
47995 => "0111110011110000",
47996 => "0111110011110000",
47997 => "0111110011110000",
47998 => "0111110011110000",
47999 => "0111110011110000",
48000 => "0111110011110000",
48001 => "0111110100000000",
48002 => "0111110100000000",
48003 => "0111110100000000",
48004 => "0111110100000000",
48005 => "0111110100000000",
48006 => "0111110100000000",
48007 => "0111110100000000",
48008 => "0111110100000000",
48009 => "0111110100000000",
48010 => "0111110100000000",
48011 => "0111110100000000",
48012 => "0111110100000000",
48013 => "0111110100000000",
48014 => "0111110100000000",
48015 => "0111110100000000",
48016 => "0111110100000000",
48017 => "0111110100000000",
48018 => "0111110100000000",
48019 => "0111110100000000",
48020 => "0111110100000000",
48021 => "0111110100000000",
48022 => "0111110100000000",
48023 => "0111110100000000",
48024 => "0111110100000000",
48025 => "0111110100000000",
48026 => "0111110100000000",
48027 => "0111110100000000",
48028 => "0111110100000000",
48029 => "0111110100000000",
48030 => "0111110100000000",
48031 => "0111110100000000",
48032 => "0111110100000000",
48033 => "0111110100000000",
48034 => "0111110100000000",
48035 => "0111110100000000",
48036 => "0111110100000000",
48037 => "0111110100000000",
48038 => "0111110100000000",
48039 => "0111110100000000",
48040 => "0111110100000000",
48041 => "0111110100000000",
48042 => "0111110100000000",
48043 => "0111110100000000",
48044 => "0111110100000000",
48045 => "0111110100000000",
48046 => "0111110100000000",
48047 => "0111110100000000",
48048 => "0111110100000000",
48049 => "0111110100000000",
48050 => "0111110100000000",
48051 => "0111110100000000",
48052 => "0111110100000000",
48053 => "0111110100000000",
48054 => "0111110100000000",
48055 => "0111110100000000",
48056 => "0111110100000000",
48057 => "0111110100000000",
48058 => "0111110100000000",
48059 => "0111110100000000",
48060 => "0111110100000000",
48061 => "0111110100000000",
48062 => "0111110100000000",
48063 => "0111110100000000",
48064 => "0111110100000000",
48065 => "0111110100000000",
48066 => "0111110100000000",
48067 => "0111110100000000",
48068 => "0111110100000000",
48069 => "0111110100000000",
48070 => "0111110100000000",
48071 => "0111110100000000",
48072 => "0111110100000000",
48073 => "0111110100000000",
48074 => "0111110100000000",
48075 => "0111110100000000",
48076 => "0111110100000000",
48077 => "0111110100000000",
48078 => "0111110100000000",
48079 => "0111110100000000",
48080 => "0111110100000000",
48081 => "0111110100000000",
48082 => "0111110100000000",
48083 => "0111110100000000",
48084 => "0111110100000000",
48085 => "0111110100000000",
48086 => "0111110100000000",
48087 => "0111110100000000",
48088 => "0111110100000000",
48089 => "0111110100010000",
48090 => "0111110100010000",
48091 => "0111110100010000",
48092 => "0111110100010000",
48093 => "0111110100010000",
48094 => "0111110100010000",
48095 => "0111110100010000",
48096 => "0111110100010000",
48097 => "0111110100010000",
48098 => "0111110100010000",
48099 => "0111110100010000",
48100 => "0111110100010000",
48101 => "0111110100010000",
48102 => "0111110100010000",
48103 => "0111110100010000",
48104 => "0111110100010000",
48105 => "0111110100010000",
48106 => "0111110100010000",
48107 => "0111110100010000",
48108 => "0111110100010000",
48109 => "0111110100010000",
48110 => "0111110100010000",
48111 => "0111110100010000",
48112 => "0111110100010000",
48113 => "0111110100010000",
48114 => "0111110100010000",
48115 => "0111110100010000",
48116 => "0111110100010000",
48117 => "0111110100010000",
48118 => "0111110100010000",
48119 => "0111110100010000",
48120 => "0111110100010000",
48121 => "0111110100010000",
48122 => "0111110100010000",
48123 => "0111110100010000",
48124 => "0111110100010000",
48125 => "0111110100010000",
48126 => "0111110100010000",
48127 => "0111110100010000",
48128 => "0111110100010000",
48129 => "0111110100010000",
48130 => "0111110100010000",
48131 => "0111110100010000",
48132 => "0111110100010000",
48133 => "0111110100010000",
48134 => "0111110100010000",
48135 => "0111110100010000",
48136 => "0111110100010000",
48137 => "0111110100010000",
48138 => "0111110100010000",
48139 => "0111110100010000",
48140 => "0111110100010000",
48141 => "0111110100010000",
48142 => "0111110100010000",
48143 => "0111110100010000",
48144 => "0111110100010000",
48145 => "0111110100010000",
48146 => "0111110100010000",
48147 => "0111110100010000",
48148 => "0111110100010000",
48149 => "0111110100010000",
48150 => "0111110100010000",
48151 => "0111110100010000",
48152 => "0111110100010000",
48153 => "0111110100010000",
48154 => "0111110100010000",
48155 => "0111110100010000",
48156 => "0111110100010000",
48157 => "0111110100010000",
48158 => "0111110100010000",
48159 => "0111110100010000",
48160 => "0111110100010000",
48161 => "0111110100010000",
48162 => "0111110100010000",
48163 => "0111110100010000",
48164 => "0111110100010000",
48165 => "0111110100010000",
48166 => "0111110100010000",
48167 => "0111110100010000",
48168 => "0111110100010000",
48169 => "0111110100010000",
48170 => "0111110100010000",
48171 => "0111110100010000",
48172 => "0111110100010000",
48173 => "0111110100010000",
48174 => "0111110100010000",
48175 => "0111110100010000",
48176 => "0111110100010000",
48177 => "0111110100010000",
48178 => "0111110100100000",
48179 => "0111110100100000",
48180 => "0111110100100000",
48181 => "0111110100100000",
48182 => "0111110100100000",
48183 => "0111110100100000",
48184 => "0111110100100000",
48185 => "0111110100100000",
48186 => "0111110100100000",
48187 => "0111110100100000",
48188 => "0111110100100000",
48189 => "0111110100100000",
48190 => "0111110100100000",
48191 => "0111110100100000",
48192 => "0111110100100000",
48193 => "0111110100100000",
48194 => "0111110100100000",
48195 => "0111110100100000",
48196 => "0111110100100000",
48197 => "0111110100100000",
48198 => "0111110100100000",
48199 => "0111110100100000",
48200 => "0111110100100000",
48201 => "0111110100100000",
48202 => "0111110100100000",
48203 => "0111110100100000",
48204 => "0111110100100000",
48205 => "0111110100100000",
48206 => "0111110100100000",
48207 => "0111110100100000",
48208 => "0111110100100000",
48209 => "0111110100100000",
48210 => "0111110100100000",
48211 => "0111110100100000",
48212 => "0111110100100000",
48213 => "0111110100100000",
48214 => "0111110100100000",
48215 => "0111110100100000",
48216 => "0111110100100000",
48217 => "0111110100100000",
48218 => "0111110100100000",
48219 => "0111110100100000",
48220 => "0111110100100000",
48221 => "0111110100100000",
48222 => "0111110100100000",
48223 => "0111110100100000",
48224 => "0111110100100000",
48225 => "0111110100100000",
48226 => "0111110100100000",
48227 => "0111110100100000",
48228 => "0111110100100000",
48229 => "0111110100100000",
48230 => "0111110100100000",
48231 => "0111110100100000",
48232 => "0111110100100000",
48233 => "0111110100100000",
48234 => "0111110100100000",
48235 => "0111110100100000",
48236 => "0111110100100000",
48237 => "0111110100100000",
48238 => "0111110100100000",
48239 => "0111110100100000",
48240 => "0111110100100000",
48241 => "0111110100100000",
48242 => "0111110100100000",
48243 => "0111110100100000",
48244 => "0111110100100000",
48245 => "0111110100100000",
48246 => "0111110100100000",
48247 => "0111110100100000",
48248 => "0111110100100000",
48249 => "0111110100100000",
48250 => "0111110100100000",
48251 => "0111110100100000",
48252 => "0111110100100000",
48253 => "0111110100100000",
48254 => "0111110100100000",
48255 => "0111110100100000",
48256 => "0111110100100000",
48257 => "0111110100100000",
48258 => "0111110100100000",
48259 => "0111110100100000",
48260 => "0111110100100000",
48261 => "0111110100100000",
48262 => "0111110100100000",
48263 => "0111110100100000",
48264 => "0111110100100000",
48265 => "0111110100100000",
48266 => "0111110100100000",
48267 => "0111110100100000",
48268 => "0111110100100000",
48269 => "0111110100110000",
48270 => "0111110100110000",
48271 => "0111110100110000",
48272 => "0111110100110000",
48273 => "0111110100110000",
48274 => "0111110100110000",
48275 => "0111110100110000",
48276 => "0111110100110000",
48277 => "0111110100110000",
48278 => "0111110100110000",
48279 => "0111110100110000",
48280 => "0111110100110000",
48281 => "0111110100110000",
48282 => "0111110100110000",
48283 => "0111110100110000",
48284 => "0111110100110000",
48285 => "0111110100110000",
48286 => "0111110100110000",
48287 => "0111110100110000",
48288 => "0111110100110000",
48289 => "0111110100110000",
48290 => "0111110100110000",
48291 => "0111110100110000",
48292 => "0111110100110000",
48293 => "0111110100110000",
48294 => "0111110100110000",
48295 => "0111110100110000",
48296 => "0111110100110000",
48297 => "0111110100110000",
48298 => "0111110100110000",
48299 => "0111110100110000",
48300 => "0111110100110000",
48301 => "0111110100110000",
48302 => "0111110100110000",
48303 => "0111110100110000",
48304 => "0111110100110000",
48305 => "0111110100110000",
48306 => "0111110100110000",
48307 => "0111110100110000",
48308 => "0111110100110000",
48309 => "0111110100110000",
48310 => "0111110100110000",
48311 => "0111110100110000",
48312 => "0111110100110000",
48313 => "0111110100110000",
48314 => "0111110100110000",
48315 => "0111110100110000",
48316 => "0111110100110000",
48317 => "0111110100110000",
48318 => "0111110100110000",
48319 => "0111110100110000",
48320 => "0111110100110000",
48321 => "0111110100110000",
48322 => "0111110100110000",
48323 => "0111110100110000",
48324 => "0111110100110000",
48325 => "0111110100110000",
48326 => "0111110100110000",
48327 => "0111110100110000",
48328 => "0111110100110000",
48329 => "0111110100110000",
48330 => "0111110100110000",
48331 => "0111110100110000",
48332 => "0111110100110000",
48333 => "0111110100110000",
48334 => "0111110100110000",
48335 => "0111110100110000",
48336 => "0111110100110000",
48337 => "0111110100110000",
48338 => "0111110100110000",
48339 => "0111110100110000",
48340 => "0111110100110000",
48341 => "0111110100110000",
48342 => "0111110100110000",
48343 => "0111110100110000",
48344 => "0111110100110000",
48345 => "0111110100110000",
48346 => "0111110100110000",
48347 => "0111110100110000",
48348 => "0111110100110000",
48349 => "0111110100110000",
48350 => "0111110100110000",
48351 => "0111110100110000",
48352 => "0111110100110000",
48353 => "0111110100110000",
48354 => "0111110100110000",
48355 => "0111110100110000",
48356 => "0111110100110000",
48357 => "0111110100110000",
48358 => "0111110100110000",
48359 => "0111110100110000",
48360 => "0111110100110000",
48361 => "0111110100110000",
48362 => "0111110101000000",
48363 => "0111110101000000",
48364 => "0111110101000000",
48365 => "0111110101000000",
48366 => "0111110101000000",
48367 => "0111110101000000",
48368 => "0111110101000000",
48369 => "0111110101000000",
48370 => "0111110101000000",
48371 => "0111110101000000",
48372 => "0111110101000000",
48373 => "0111110101000000",
48374 => "0111110101000000",
48375 => "0111110101000000",
48376 => "0111110101000000",
48377 => "0111110101000000",
48378 => "0111110101000000",
48379 => "0111110101000000",
48380 => "0111110101000000",
48381 => "0111110101000000",
48382 => "0111110101000000",
48383 => "0111110101000000",
48384 => "0111110101000000",
48385 => "0111110101000000",
48386 => "0111110101000000",
48387 => "0111110101000000",
48388 => "0111110101000000",
48389 => "0111110101000000",
48390 => "0111110101000000",
48391 => "0111110101000000",
48392 => "0111110101000000",
48393 => "0111110101000000",
48394 => "0111110101000000",
48395 => "0111110101000000",
48396 => "0111110101000000",
48397 => "0111110101000000",
48398 => "0111110101000000",
48399 => "0111110101000000",
48400 => "0111110101000000",
48401 => "0111110101000000",
48402 => "0111110101000000",
48403 => "0111110101000000",
48404 => "0111110101000000",
48405 => "0111110101000000",
48406 => "0111110101000000",
48407 => "0111110101000000",
48408 => "0111110101000000",
48409 => "0111110101000000",
48410 => "0111110101000000",
48411 => "0111110101000000",
48412 => "0111110101000000",
48413 => "0111110101000000",
48414 => "0111110101000000",
48415 => "0111110101000000",
48416 => "0111110101000000",
48417 => "0111110101000000",
48418 => "0111110101000000",
48419 => "0111110101000000",
48420 => "0111110101000000",
48421 => "0111110101000000",
48422 => "0111110101000000",
48423 => "0111110101000000",
48424 => "0111110101000000",
48425 => "0111110101000000",
48426 => "0111110101000000",
48427 => "0111110101000000",
48428 => "0111110101000000",
48429 => "0111110101000000",
48430 => "0111110101000000",
48431 => "0111110101000000",
48432 => "0111110101000000",
48433 => "0111110101000000",
48434 => "0111110101000000",
48435 => "0111110101000000",
48436 => "0111110101000000",
48437 => "0111110101000000",
48438 => "0111110101000000",
48439 => "0111110101000000",
48440 => "0111110101000000",
48441 => "0111110101000000",
48442 => "0111110101000000",
48443 => "0111110101000000",
48444 => "0111110101000000",
48445 => "0111110101000000",
48446 => "0111110101000000",
48447 => "0111110101000000",
48448 => "0111110101000000",
48449 => "0111110101000000",
48450 => "0111110101000000",
48451 => "0111110101000000",
48452 => "0111110101000000",
48453 => "0111110101000000",
48454 => "0111110101000000",
48455 => "0111110101000000",
48456 => "0111110101000000",
48457 => "0111110101010000",
48458 => "0111110101010000",
48459 => "0111110101010000",
48460 => "0111110101010000",
48461 => "0111110101010000",
48462 => "0111110101010000",
48463 => "0111110101010000",
48464 => "0111110101010000",
48465 => "0111110101010000",
48466 => "0111110101010000",
48467 => "0111110101010000",
48468 => "0111110101010000",
48469 => "0111110101010000",
48470 => "0111110101010000",
48471 => "0111110101010000",
48472 => "0111110101010000",
48473 => "0111110101010000",
48474 => "0111110101010000",
48475 => "0111110101010000",
48476 => "0111110101010000",
48477 => "0111110101010000",
48478 => "0111110101010000",
48479 => "0111110101010000",
48480 => "0111110101010000",
48481 => "0111110101010000",
48482 => "0111110101010000",
48483 => "0111110101010000",
48484 => "0111110101010000",
48485 => "0111110101010000",
48486 => "0111110101010000",
48487 => "0111110101010000",
48488 => "0111110101010000",
48489 => "0111110101010000",
48490 => "0111110101010000",
48491 => "0111110101010000",
48492 => "0111110101010000",
48493 => "0111110101010000",
48494 => "0111110101010000",
48495 => "0111110101010000",
48496 => "0111110101010000",
48497 => "0111110101010000",
48498 => "0111110101010000",
48499 => "0111110101010000",
48500 => "0111110101010000",
48501 => "0111110101010000",
48502 => "0111110101010000",
48503 => "0111110101010000",
48504 => "0111110101010000",
48505 => "0111110101010000",
48506 => "0111110101010000",
48507 => "0111110101010000",
48508 => "0111110101010000",
48509 => "0111110101010000",
48510 => "0111110101010000",
48511 => "0111110101010000",
48512 => "0111110101010000",
48513 => "0111110101010000",
48514 => "0111110101010000",
48515 => "0111110101010000",
48516 => "0111110101010000",
48517 => "0111110101010000",
48518 => "0111110101010000",
48519 => "0111110101010000",
48520 => "0111110101010000",
48521 => "0111110101010000",
48522 => "0111110101010000",
48523 => "0111110101010000",
48524 => "0111110101010000",
48525 => "0111110101010000",
48526 => "0111110101010000",
48527 => "0111110101010000",
48528 => "0111110101010000",
48529 => "0111110101010000",
48530 => "0111110101010000",
48531 => "0111110101010000",
48532 => "0111110101010000",
48533 => "0111110101010000",
48534 => "0111110101010000",
48535 => "0111110101010000",
48536 => "0111110101010000",
48537 => "0111110101010000",
48538 => "0111110101010000",
48539 => "0111110101010000",
48540 => "0111110101010000",
48541 => "0111110101010000",
48542 => "0111110101010000",
48543 => "0111110101010000",
48544 => "0111110101010000",
48545 => "0111110101010000",
48546 => "0111110101010000",
48547 => "0111110101010000",
48548 => "0111110101010000",
48549 => "0111110101010000",
48550 => "0111110101010000",
48551 => "0111110101010000",
48552 => "0111110101010000",
48553 => "0111110101010000",
48554 => "0111110101100000",
48555 => "0111110101100000",
48556 => "0111110101100000",
48557 => "0111110101100000",
48558 => "0111110101100000",
48559 => "0111110101100000",
48560 => "0111110101100000",
48561 => "0111110101100000",
48562 => "0111110101100000",
48563 => "0111110101100000",
48564 => "0111110101100000",
48565 => "0111110101100000",
48566 => "0111110101100000",
48567 => "0111110101100000",
48568 => "0111110101100000",
48569 => "0111110101100000",
48570 => "0111110101100000",
48571 => "0111110101100000",
48572 => "0111110101100000",
48573 => "0111110101100000",
48574 => "0111110101100000",
48575 => "0111110101100000",
48576 => "0111110101100000",
48577 => "0111110101100000",
48578 => "0111110101100000",
48579 => "0111110101100000",
48580 => "0111110101100000",
48581 => "0111110101100000",
48582 => "0111110101100000",
48583 => "0111110101100000",
48584 => "0111110101100000",
48585 => "0111110101100000",
48586 => "0111110101100000",
48587 => "0111110101100000",
48588 => "0111110101100000",
48589 => "0111110101100000",
48590 => "0111110101100000",
48591 => "0111110101100000",
48592 => "0111110101100000",
48593 => "0111110101100000",
48594 => "0111110101100000",
48595 => "0111110101100000",
48596 => "0111110101100000",
48597 => "0111110101100000",
48598 => "0111110101100000",
48599 => "0111110101100000",
48600 => "0111110101100000",
48601 => "0111110101100000",
48602 => "0111110101100000",
48603 => "0111110101100000",
48604 => "0111110101100000",
48605 => "0111110101100000",
48606 => "0111110101100000",
48607 => "0111110101100000",
48608 => "0111110101100000",
48609 => "0111110101100000",
48610 => "0111110101100000",
48611 => "0111110101100000",
48612 => "0111110101100000",
48613 => "0111110101100000",
48614 => "0111110101100000",
48615 => "0111110101100000",
48616 => "0111110101100000",
48617 => "0111110101100000",
48618 => "0111110101100000",
48619 => "0111110101100000",
48620 => "0111110101100000",
48621 => "0111110101100000",
48622 => "0111110101100000",
48623 => "0111110101100000",
48624 => "0111110101100000",
48625 => "0111110101100000",
48626 => "0111110101100000",
48627 => "0111110101100000",
48628 => "0111110101100000",
48629 => "0111110101100000",
48630 => "0111110101100000",
48631 => "0111110101100000",
48632 => "0111110101100000",
48633 => "0111110101100000",
48634 => "0111110101100000",
48635 => "0111110101100000",
48636 => "0111110101100000",
48637 => "0111110101100000",
48638 => "0111110101100000",
48639 => "0111110101100000",
48640 => "0111110101100000",
48641 => "0111110101100000",
48642 => "0111110101100000",
48643 => "0111110101100000",
48644 => "0111110101100000",
48645 => "0111110101100000",
48646 => "0111110101100000",
48647 => "0111110101100000",
48648 => "0111110101100000",
48649 => "0111110101100000",
48650 => "0111110101100000",
48651 => "0111110101100000",
48652 => "0111110101100000",
48653 => "0111110101100000",
48654 => "0111110101110000",
48655 => "0111110101110000",
48656 => "0111110101110000",
48657 => "0111110101110000",
48658 => "0111110101110000",
48659 => "0111110101110000",
48660 => "0111110101110000",
48661 => "0111110101110000",
48662 => "0111110101110000",
48663 => "0111110101110000",
48664 => "0111110101110000",
48665 => "0111110101110000",
48666 => "0111110101110000",
48667 => "0111110101110000",
48668 => "0111110101110000",
48669 => "0111110101110000",
48670 => "0111110101110000",
48671 => "0111110101110000",
48672 => "0111110101110000",
48673 => "0111110101110000",
48674 => "0111110101110000",
48675 => "0111110101110000",
48676 => "0111110101110000",
48677 => "0111110101110000",
48678 => "0111110101110000",
48679 => "0111110101110000",
48680 => "0111110101110000",
48681 => "0111110101110000",
48682 => "0111110101110000",
48683 => "0111110101110000",
48684 => "0111110101110000",
48685 => "0111110101110000",
48686 => "0111110101110000",
48687 => "0111110101110000",
48688 => "0111110101110000",
48689 => "0111110101110000",
48690 => "0111110101110000",
48691 => "0111110101110000",
48692 => "0111110101110000",
48693 => "0111110101110000",
48694 => "0111110101110000",
48695 => "0111110101110000",
48696 => "0111110101110000",
48697 => "0111110101110000",
48698 => "0111110101110000",
48699 => "0111110101110000",
48700 => "0111110101110000",
48701 => "0111110101110000",
48702 => "0111110101110000",
48703 => "0111110101110000",
48704 => "0111110101110000",
48705 => "0111110101110000",
48706 => "0111110101110000",
48707 => "0111110101110000",
48708 => "0111110101110000",
48709 => "0111110101110000",
48710 => "0111110101110000",
48711 => "0111110101110000",
48712 => "0111110101110000",
48713 => "0111110101110000",
48714 => "0111110101110000",
48715 => "0111110101110000",
48716 => "0111110101110000",
48717 => "0111110101110000",
48718 => "0111110101110000",
48719 => "0111110101110000",
48720 => "0111110101110000",
48721 => "0111110101110000",
48722 => "0111110101110000",
48723 => "0111110101110000",
48724 => "0111110101110000",
48725 => "0111110101110000",
48726 => "0111110101110000",
48727 => "0111110101110000",
48728 => "0111110101110000",
48729 => "0111110101110000",
48730 => "0111110101110000",
48731 => "0111110101110000",
48732 => "0111110101110000",
48733 => "0111110101110000",
48734 => "0111110101110000",
48735 => "0111110101110000",
48736 => "0111110101110000",
48737 => "0111110101110000",
48738 => "0111110101110000",
48739 => "0111110101110000",
48740 => "0111110101110000",
48741 => "0111110101110000",
48742 => "0111110101110000",
48743 => "0111110101110000",
48744 => "0111110101110000",
48745 => "0111110101110000",
48746 => "0111110101110000",
48747 => "0111110101110000",
48748 => "0111110101110000",
48749 => "0111110101110000",
48750 => "0111110101110000",
48751 => "0111110101110000",
48752 => "0111110101110000",
48753 => "0111110101110000",
48754 => "0111110101110000",
48755 => "0111110101110000",
48756 => "0111110110000000",
48757 => "0111110110000000",
48758 => "0111110110000000",
48759 => "0111110110000000",
48760 => "0111110110000000",
48761 => "0111110110000000",
48762 => "0111110110000000",
48763 => "0111110110000000",
48764 => "0111110110000000",
48765 => "0111110110000000",
48766 => "0111110110000000",
48767 => "0111110110000000",
48768 => "0111110110000000",
48769 => "0111110110000000",
48770 => "0111110110000000",
48771 => "0111110110000000",
48772 => "0111110110000000",
48773 => "0111110110000000",
48774 => "0111110110000000",
48775 => "0111110110000000",
48776 => "0111110110000000",
48777 => "0111110110000000",
48778 => "0111110110000000",
48779 => "0111110110000000",
48780 => "0111110110000000",
48781 => "0111110110000000",
48782 => "0111110110000000",
48783 => "0111110110000000",
48784 => "0111110110000000",
48785 => "0111110110000000",
48786 => "0111110110000000",
48787 => "0111110110000000",
48788 => "0111110110000000",
48789 => "0111110110000000",
48790 => "0111110110000000",
48791 => "0111110110000000",
48792 => "0111110110000000",
48793 => "0111110110000000",
48794 => "0111110110000000",
48795 => "0111110110000000",
48796 => "0111110110000000",
48797 => "0111110110000000",
48798 => "0111110110000000",
48799 => "0111110110000000",
48800 => "0111110110000000",
48801 => "0111110110000000",
48802 => "0111110110000000",
48803 => "0111110110000000",
48804 => "0111110110000000",
48805 => "0111110110000000",
48806 => "0111110110000000",
48807 => "0111110110000000",
48808 => "0111110110000000",
48809 => "0111110110000000",
48810 => "0111110110000000",
48811 => "0111110110000000",
48812 => "0111110110000000",
48813 => "0111110110000000",
48814 => "0111110110000000",
48815 => "0111110110000000",
48816 => "0111110110000000",
48817 => "0111110110000000",
48818 => "0111110110000000",
48819 => "0111110110000000",
48820 => "0111110110000000",
48821 => "0111110110000000",
48822 => "0111110110000000",
48823 => "0111110110000000",
48824 => "0111110110000000",
48825 => "0111110110000000",
48826 => "0111110110000000",
48827 => "0111110110000000",
48828 => "0111110110000000",
48829 => "0111110110000000",
48830 => "0111110110000000",
48831 => "0111110110000000",
48832 => "0111110110000000",
48833 => "0111110110000000",
48834 => "0111110110000000",
48835 => "0111110110000000",
48836 => "0111110110000000",
48837 => "0111110110000000",
48838 => "0111110110000000",
48839 => "0111110110000000",
48840 => "0111110110000000",
48841 => "0111110110000000",
48842 => "0111110110000000",
48843 => "0111110110000000",
48844 => "0111110110000000",
48845 => "0111110110000000",
48846 => "0111110110000000",
48847 => "0111110110000000",
48848 => "0111110110000000",
48849 => "0111110110000000",
48850 => "0111110110000000",
48851 => "0111110110000000",
48852 => "0111110110000000",
48853 => "0111110110000000",
48854 => "0111110110000000",
48855 => "0111110110000000",
48856 => "0111110110000000",
48857 => "0111110110000000",
48858 => "0111110110000000",
48859 => "0111110110000000",
48860 => "0111110110010000",
48861 => "0111110110010000",
48862 => "0111110110010000",
48863 => "0111110110010000",
48864 => "0111110110010000",
48865 => "0111110110010000",
48866 => "0111110110010000",
48867 => "0111110110010000",
48868 => "0111110110010000",
48869 => "0111110110010000",
48870 => "0111110110010000",
48871 => "0111110110010000",
48872 => "0111110110010000",
48873 => "0111110110010000",
48874 => "0111110110010000",
48875 => "0111110110010000",
48876 => "0111110110010000",
48877 => "0111110110010000",
48878 => "0111110110010000",
48879 => "0111110110010000",
48880 => "0111110110010000",
48881 => "0111110110010000",
48882 => "0111110110010000",
48883 => "0111110110010000",
48884 => "0111110110010000",
48885 => "0111110110010000",
48886 => "0111110110010000",
48887 => "0111110110010000",
48888 => "0111110110010000",
48889 => "0111110110010000",
48890 => "0111110110010000",
48891 => "0111110110010000",
48892 => "0111110110010000",
48893 => "0111110110010000",
48894 => "0111110110010000",
48895 => "0111110110010000",
48896 => "0111110110010000",
48897 => "0111110110010000",
48898 => "0111110110010000",
48899 => "0111110110010000",
48900 => "0111110110010000",
48901 => "0111110110010000",
48902 => "0111110110010000",
48903 => "0111110110010000",
48904 => "0111110110010000",
48905 => "0111110110010000",
48906 => "0111110110010000",
48907 => "0111110110010000",
48908 => "0111110110010000",
48909 => "0111110110010000",
48910 => "0111110110010000",
48911 => "0111110110010000",
48912 => "0111110110010000",
48913 => "0111110110010000",
48914 => "0111110110010000",
48915 => "0111110110010000",
48916 => "0111110110010000",
48917 => "0111110110010000",
48918 => "0111110110010000",
48919 => "0111110110010000",
48920 => "0111110110010000",
48921 => "0111110110010000",
48922 => "0111110110010000",
48923 => "0111110110010000",
48924 => "0111110110010000",
48925 => "0111110110010000",
48926 => "0111110110010000",
48927 => "0111110110010000",
48928 => "0111110110010000",
48929 => "0111110110010000",
48930 => "0111110110010000",
48931 => "0111110110010000",
48932 => "0111110110010000",
48933 => "0111110110010000",
48934 => "0111110110010000",
48935 => "0111110110010000",
48936 => "0111110110010000",
48937 => "0111110110010000",
48938 => "0111110110010000",
48939 => "0111110110010000",
48940 => "0111110110010000",
48941 => "0111110110010000",
48942 => "0111110110010000",
48943 => "0111110110010000",
48944 => "0111110110010000",
48945 => "0111110110010000",
48946 => "0111110110010000",
48947 => "0111110110010000",
48948 => "0111110110010000",
48949 => "0111110110010000",
48950 => "0111110110010000",
48951 => "0111110110010000",
48952 => "0111110110010000",
48953 => "0111110110010000",
48954 => "0111110110010000",
48955 => "0111110110010000",
48956 => "0111110110010000",
48957 => "0111110110010000",
48958 => "0111110110010000",
48959 => "0111110110010000",
48960 => "0111110110010000",
48961 => "0111110110010000",
48962 => "0111110110010000",
48963 => "0111110110010000",
48964 => "0111110110010000",
48965 => "0111110110010000",
48966 => "0111110110010000",
48967 => "0111110110100000",
48968 => "0111110110100000",
48969 => "0111110110100000",
48970 => "0111110110100000",
48971 => "0111110110100000",
48972 => "0111110110100000",
48973 => "0111110110100000",
48974 => "0111110110100000",
48975 => "0111110110100000",
48976 => "0111110110100000",
48977 => "0111110110100000",
48978 => "0111110110100000",
48979 => "0111110110100000",
48980 => "0111110110100000",
48981 => "0111110110100000",
48982 => "0111110110100000",
48983 => "0111110110100000",
48984 => "0111110110100000",
48985 => "0111110110100000",
48986 => "0111110110100000",
48987 => "0111110110100000",
48988 => "0111110110100000",
48989 => "0111110110100000",
48990 => "0111110110100000",
48991 => "0111110110100000",
48992 => "0111110110100000",
48993 => "0111110110100000",
48994 => "0111110110100000",
48995 => "0111110110100000",
48996 => "0111110110100000",
48997 => "0111110110100000",
48998 => "0111110110100000",
48999 => "0111110110100000",
49000 => "0111110110100000",
49001 => "0111110110100000",
49002 => "0111110110100000",
49003 => "0111110110100000",
49004 => "0111110110100000",
49005 => "0111110110100000",
49006 => "0111110110100000",
49007 => "0111110110100000",
49008 => "0111110110100000",
49009 => "0111110110100000",
49010 => "0111110110100000",
49011 => "0111110110100000",
49012 => "0111110110100000",
49013 => "0111110110100000",
49014 => "0111110110100000",
49015 => "0111110110100000",
49016 => "0111110110100000",
49017 => "0111110110100000",
49018 => "0111110110100000",
49019 => "0111110110100000",
49020 => "0111110110100000",
49021 => "0111110110100000",
49022 => "0111110110100000",
49023 => "0111110110100000",
49024 => "0111110110100000",
49025 => "0111110110100000",
49026 => "0111110110100000",
49027 => "0111110110100000",
49028 => "0111110110100000",
49029 => "0111110110100000",
49030 => "0111110110100000",
49031 => "0111110110100000",
49032 => "0111110110100000",
49033 => "0111110110100000",
49034 => "0111110110100000",
49035 => "0111110110100000",
49036 => "0111110110100000",
49037 => "0111110110100000",
49038 => "0111110110100000",
49039 => "0111110110100000",
49040 => "0111110110100000",
49041 => "0111110110100000",
49042 => "0111110110100000",
49043 => "0111110110100000",
49044 => "0111110110100000",
49045 => "0111110110100000",
49046 => "0111110110100000",
49047 => "0111110110100000",
49048 => "0111110110100000",
49049 => "0111110110100000",
49050 => "0111110110100000",
49051 => "0111110110100000",
49052 => "0111110110100000",
49053 => "0111110110100000",
49054 => "0111110110100000",
49055 => "0111110110100000",
49056 => "0111110110100000",
49057 => "0111110110100000",
49058 => "0111110110100000",
49059 => "0111110110100000",
49060 => "0111110110100000",
49061 => "0111110110100000",
49062 => "0111110110100000",
49063 => "0111110110100000",
49064 => "0111110110100000",
49065 => "0111110110100000",
49066 => "0111110110100000",
49067 => "0111110110100000",
49068 => "0111110110100000",
49069 => "0111110110100000",
49070 => "0111110110100000",
49071 => "0111110110100000",
49072 => "0111110110100000",
49073 => "0111110110100000",
49074 => "0111110110100000",
49075 => "0111110110100000",
49076 => "0111110110100000",
49077 => "0111110110110000",
49078 => "0111110110110000",
49079 => "0111110110110000",
49080 => "0111110110110000",
49081 => "0111110110110000",
49082 => "0111110110110000",
49083 => "0111110110110000",
49084 => "0111110110110000",
49085 => "0111110110110000",
49086 => "0111110110110000",
49087 => "0111110110110000",
49088 => "0111110110110000",
49089 => "0111110110110000",
49090 => "0111110110110000",
49091 => "0111110110110000",
49092 => "0111110110110000",
49093 => "0111110110110000",
49094 => "0111110110110000",
49095 => "0111110110110000",
49096 => "0111110110110000",
49097 => "0111110110110000",
49098 => "0111110110110000",
49099 => "0111110110110000",
49100 => "0111110110110000",
49101 => "0111110110110000",
49102 => "0111110110110000",
49103 => "0111110110110000",
49104 => "0111110110110000",
49105 => "0111110110110000",
49106 => "0111110110110000",
49107 => "0111110110110000",
49108 => "0111110110110000",
49109 => "0111110110110000",
49110 => "0111110110110000",
49111 => "0111110110110000",
49112 => "0111110110110000",
49113 => "0111110110110000",
49114 => "0111110110110000",
49115 => "0111110110110000",
49116 => "0111110110110000",
49117 => "0111110110110000",
49118 => "0111110110110000",
49119 => "0111110110110000",
49120 => "0111110110110000",
49121 => "0111110110110000",
49122 => "0111110110110000",
49123 => "0111110110110000",
49124 => "0111110110110000",
49125 => "0111110110110000",
49126 => "0111110110110000",
49127 => "0111110110110000",
49128 => "0111110110110000",
49129 => "0111110110110000",
49130 => "0111110110110000",
49131 => "0111110110110000",
49132 => "0111110110110000",
49133 => "0111110110110000",
49134 => "0111110110110000",
49135 => "0111110110110000",
49136 => "0111110110110000",
49137 => "0111110110110000",
49138 => "0111110110110000",
49139 => "0111110110110000",
49140 => "0111110110110000",
49141 => "0111110110110000",
49142 => "0111110110110000",
49143 => "0111110110110000",
49144 => "0111110110110000",
49145 => "0111110110110000",
49146 => "0111110110110000",
49147 => "0111110110110000",
49148 => "0111110110110000",
49149 => "0111110110110000",
49150 => "0111110110110000",
49151 => "0111110110110000",
49152 => "0111110110110000",
49153 => "0111110110110000",
49154 => "0111110110110000",
49155 => "0111110110110000",
49156 => "0111110110110000",
49157 => "0111110110110000",
49158 => "0111110110110000",
49159 => "0111110110110000",
49160 => "0111110110110000",
49161 => "0111110110110000",
49162 => "0111110110110000",
49163 => "0111110110110000",
49164 => "0111110110110000",
49165 => "0111110110110000",
49166 => "0111110110110000",
49167 => "0111110110110000",
49168 => "0111110110110000",
49169 => "0111110110110000",
49170 => "0111110110110000",
49171 => "0111110110110000",
49172 => "0111110110110000",
49173 => "0111110110110000",
49174 => "0111110110110000",
49175 => "0111110110110000",
49176 => "0111110110110000",
49177 => "0111110110110000",
49178 => "0111110110110000",
49179 => "0111110110110000",
49180 => "0111110110110000",
49181 => "0111110110110000",
49182 => "0111110110110000",
49183 => "0111110110110000",
49184 => "0111110110110000",
49185 => "0111110110110000",
49186 => "0111110110110000",
49187 => "0111110110110000",
49188 => "0111110110110000",
49189 => "0111110110110000",
49190 => "0111110111000000",
49191 => "0111110111000000",
49192 => "0111110111000000",
49193 => "0111110111000000",
49194 => "0111110111000000",
49195 => "0111110111000000",
49196 => "0111110111000000",
49197 => "0111110111000000",
49198 => "0111110111000000",
49199 => "0111110111000000",
49200 => "0111110111000000",
49201 => "0111110111000000",
49202 => "0111110111000000",
49203 => "0111110111000000",
49204 => "0111110111000000",
49205 => "0111110111000000",
49206 => "0111110111000000",
49207 => "0111110111000000",
49208 => "0111110111000000",
49209 => "0111110111000000",
49210 => "0111110111000000",
49211 => "0111110111000000",
49212 => "0111110111000000",
49213 => "0111110111000000",
49214 => "0111110111000000",
49215 => "0111110111000000",
49216 => "0111110111000000",
49217 => "0111110111000000",
49218 => "0111110111000000",
49219 => "0111110111000000",
49220 => "0111110111000000",
49221 => "0111110111000000",
49222 => "0111110111000000",
49223 => "0111110111000000",
49224 => "0111110111000000",
49225 => "0111110111000000",
49226 => "0111110111000000",
49227 => "0111110111000000",
49228 => "0111110111000000",
49229 => "0111110111000000",
49230 => "0111110111000000",
49231 => "0111110111000000",
49232 => "0111110111000000",
49233 => "0111110111000000",
49234 => "0111110111000000",
49235 => "0111110111000000",
49236 => "0111110111000000",
49237 => "0111110111000000",
49238 => "0111110111000000",
49239 => "0111110111000000",
49240 => "0111110111000000",
49241 => "0111110111000000",
49242 => "0111110111000000",
49243 => "0111110111000000",
49244 => "0111110111000000",
49245 => "0111110111000000",
49246 => "0111110111000000",
49247 => "0111110111000000",
49248 => "0111110111000000",
49249 => "0111110111000000",
49250 => "0111110111000000",
49251 => "0111110111000000",
49252 => "0111110111000000",
49253 => "0111110111000000",
49254 => "0111110111000000",
49255 => "0111110111000000",
49256 => "0111110111000000",
49257 => "0111110111000000",
49258 => "0111110111000000",
49259 => "0111110111000000",
49260 => "0111110111000000",
49261 => "0111110111000000",
49262 => "0111110111000000",
49263 => "0111110111000000",
49264 => "0111110111000000",
49265 => "0111110111000000",
49266 => "0111110111000000",
49267 => "0111110111000000",
49268 => "0111110111000000",
49269 => "0111110111000000",
49270 => "0111110111000000",
49271 => "0111110111000000",
49272 => "0111110111000000",
49273 => "0111110111000000",
49274 => "0111110111000000",
49275 => "0111110111000000",
49276 => "0111110111000000",
49277 => "0111110111000000",
49278 => "0111110111000000",
49279 => "0111110111000000",
49280 => "0111110111000000",
49281 => "0111110111000000",
49282 => "0111110111000000",
49283 => "0111110111000000",
49284 => "0111110111000000",
49285 => "0111110111000000",
49286 => "0111110111000000",
49287 => "0111110111000000",
49288 => "0111110111000000",
49289 => "0111110111000000",
49290 => "0111110111000000",
49291 => "0111110111000000",
49292 => "0111110111000000",
49293 => "0111110111000000",
49294 => "0111110111000000",
49295 => "0111110111000000",
49296 => "0111110111000000",
49297 => "0111110111000000",
49298 => "0111110111000000",
49299 => "0111110111000000",
49300 => "0111110111000000",
49301 => "0111110111000000",
49302 => "0111110111000000",
49303 => "0111110111000000",
49304 => "0111110111000000",
49305 => "0111110111000000",
49306 => "0111110111010000",
49307 => "0111110111010000",
49308 => "0111110111010000",
49309 => "0111110111010000",
49310 => "0111110111010000",
49311 => "0111110111010000",
49312 => "0111110111010000",
49313 => "0111110111010000",
49314 => "0111110111010000",
49315 => "0111110111010000",
49316 => "0111110111010000",
49317 => "0111110111010000",
49318 => "0111110111010000",
49319 => "0111110111010000",
49320 => "0111110111010000",
49321 => "0111110111010000",
49322 => "0111110111010000",
49323 => "0111110111010000",
49324 => "0111110111010000",
49325 => "0111110111010000",
49326 => "0111110111010000",
49327 => "0111110111010000",
49328 => "0111110111010000",
49329 => "0111110111010000",
49330 => "0111110111010000",
49331 => "0111110111010000",
49332 => "0111110111010000",
49333 => "0111110111010000",
49334 => "0111110111010000",
49335 => "0111110111010000",
49336 => "0111110111010000",
49337 => "0111110111010000",
49338 => "0111110111010000",
49339 => "0111110111010000",
49340 => "0111110111010000",
49341 => "0111110111010000",
49342 => "0111110111010000",
49343 => "0111110111010000",
49344 => "0111110111010000",
49345 => "0111110111010000",
49346 => "0111110111010000",
49347 => "0111110111010000",
49348 => "0111110111010000",
49349 => "0111110111010000",
49350 => "0111110111010000",
49351 => "0111110111010000",
49352 => "0111110111010000",
49353 => "0111110111010000",
49354 => "0111110111010000",
49355 => "0111110111010000",
49356 => "0111110111010000",
49357 => "0111110111010000",
49358 => "0111110111010000",
49359 => "0111110111010000",
49360 => "0111110111010000",
49361 => "0111110111010000",
49362 => "0111110111010000",
49363 => "0111110111010000",
49364 => "0111110111010000",
49365 => "0111110111010000",
49366 => "0111110111010000",
49367 => "0111110111010000",
49368 => "0111110111010000",
49369 => "0111110111010000",
49370 => "0111110111010000",
49371 => "0111110111010000",
49372 => "0111110111010000",
49373 => "0111110111010000",
49374 => "0111110111010000",
49375 => "0111110111010000",
49376 => "0111110111010000",
49377 => "0111110111010000",
49378 => "0111110111010000",
49379 => "0111110111010000",
49380 => "0111110111010000",
49381 => "0111110111010000",
49382 => "0111110111010000",
49383 => "0111110111010000",
49384 => "0111110111010000",
49385 => "0111110111010000",
49386 => "0111110111010000",
49387 => "0111110111010000",
49388 => "0111110111010000",
49389 => "0111110111010000",
49390 => "0111110111010000",
49391 => "0111110111010000",
49392 => "0111110111010000",
49393 => "0111110111010000",
49394 => "0111110111010000",
49395 => "0111110111010000",
49396 => "0111110111010000",
49397 => "0111110111010000",
49398 => "0111110111010000",
49399 => "0111110111010000",
49400 => "0111110111010000",
49401 => "0111110111010000",
49402 => "0111110111010000",
49403 => "0111110111010000",
49404 => "0111110111010000",
49405 => "0111110111010000",
49406 => "0111110111010000",
49407 => "0111110111010000",
49408 => "0111110111010000",
49409 => "0111110111010000",
49410 => "0111110111010000",
49411 => "0111110111010000",
49412 => "0111110111010000",
49413 => "0111110111010000",
49414 => "0111110111010000",
49415 => "0111110111010000",
49416 => "0111110111010000",
49417 => "0111110111010000",
49418 => "0111110111010000",
49419 => "0111110111010000",
49420 => "0111110111010000",
49421 => "0111110111010000",
49422 => "0111110111010000",
49423 => "0111110111010000",
49424 => "0111110111010000",
49425 => "0111110111100000",
49426 => "0111110111100000",
49427 => "0111110111100000",
49428 => "0111110111100000",
49429 => "0111110111100000",
49430 => "0111110111100000",
49431 => "0111110111100000",
49432 => "0111110111100000",
49433 => "0111110111100000",
49434 => "0111110111100000",
49435 => "0111110111100000",
49436 => "0111110111100000",
49437 => "0111110111100000",
49438 => "0111110111100000",
49439 => "0111110111100000",
49440 => "0111110111100000",
49441 => "0111110111100000",
49442 => "0111110111100000",
49443 => "0111110111100000",
49444 => "0111110111100000",
49445 => "0111110111100000",
49446 => "0111110111100000",
49447 => "0111110111100000",
49448 => "0111110111100000",
49449 => "0111110111100000",
49450 => "0111110111100000",
49451 => "0111110111100000",
49452 => "0111110111100000",
49453 => "0111110111100000",
49454 => "0111110111100000",
49455 => "0111110111100000",
49456 => "0111110111100000",
49457 => "0111110111100000",
49458 => "0111110111100000",
49459 => "0111110111100000",
49460 => "0111110111100000",
49461 => "0111110111100000",
49462 => "0111110111100000",
49463 => "0111110111100000",
49464 => "0111110111100000",
49465 => "0111110111100000",
49466 => "0111110111100000",
49467 => "0111110111100000",
49468 => "0111110111100000",
49469 => "0111110111100000",
49470 => "0111110111100000",
49471 => "0111110111100000",
49472 => "0111110111100000",
49473 => "0111110111100000",
49474 => "0111110111100000",
49475 => "0111110111100000",
49476 => "0111110111100000",
49477 => "0111110111100000",
49478 => "0111110111100000",
49479 => "0111110111100000",
49480 => "0111110111100000",
49481 => "0111110111100000",
49482 => "0111110111100000",
49483 => "0111110111100000",
49484 => "0111110111100000",
49485 => "0111110111100000",
49486 => "0111110111100000",
49487 => "0111110111100000",
49488 => "0111110111100000",
49489 => "0111110111100000",
49490 => "0111110111100000",
49491 => "0111110111100000",
49492 => "0111110111100000",
49493 => "0111110111100000",
49494 => "0111110111100000",
49495 => "0111110111100000",
49496 => "0111110111100000",
49497 => "0111110111100000",
49498 => "0111110111100000",
49499 => "0111110111100000",
49500 => "0111110111100000",
49501 => "0111110111100000",
49502 => "0111110111100000",
49503 => "0111110111100000",
49504 => "0111110111100000",
49505 => "0111110111100000",
49506 => "0111110111100000",
49507 => "0111110111100000",
49508 => "0111110111100000",
49509 => "0111110111100000",
49510 => "0111110111100000",
49511 => "0111110111100000",
49512 => "0111110111100000",
49513 => "0111110111100000",
49514 => "0111110111100000",
49515 => "0111110111100000",
49516 => "0111110111100000",
49517 => "0111110111100000",
49518 => "0111110111100000",
49519 => "0111110111100000",
49520 => "0111110111100000",
49521 => "0111110111100000",
49522 => "0111110111100000",
49523 => "0111110111100000",
49524 => "0111110111100000",
49525 => "0111110111100000",
49526 => "0111110111100000",
49527 => "0111110111100000",
49528 => "0111110111100000",
49529 => "0111110111100000",
49530 => "0111110111100000",
49531 => "0111110111100000",
49532 => "0111110111100000",
49533 => "0111110111100000",
49534 => "0111110111100000",
49535 => "0111110111100000",
49536 => "0111110111100000",
49537 => "0111110111100000",
49538 => "0111110111100000",
49539 => "0111110111100000",
49540 => "0111110111100000",
49541 => "0111110111100000",
49542 => "0111110111100000",
49543 => "0111110111100000",
49544 => "0111110111100000",
49545 => "0111110111100000",
49546 => "0111110111100000",
49547 => "0111110111110000",
49548 => "0111110111110000",
49549 => "0111110111110000",
49550 => "0111110111110000",
49551 => "0111110111110000",
49552 => "0111110111110000",
49553 => "0111110111110000",
49554 => "0111110111110000",
49555 => "0111110111110000",
49556 => "0111110111110000",
49557 => "0111110111110000",
49558 => "0111110111110000",
49559 => "0111110111110000",
49560 => "0111110111110000",
49561 => "0111110111110000",
49562 => "0111110111110000",
49563 => "0111110111110000",
49564 => "0111110111110000",
49565 => "0111110111110000",
49566 => "0111110111110000",
49567 => "0111110111110000",
49568 => "0111110111110000",
49569 => "0111110111110000",
49570 => "0111110111110000",
49571 => "0111110111110000",
49572 => "0111110111110000",
49573 => "0111110111110000",
49574 => "0111110111110000",
49575 => "0111110111110000",
49576 => "0111110111110000",
49577 => "0111110111110000",
49578 => "0111110111110000",
49579 => "0111110111110000",
49580 => "0111110111110000",
49581 => "0111110111110000",
49582 => "0111110111110000",
49583 => "0111110111110000",
49584 => "0111110111110000",
49585 => "0111110111110000",
49586 => "0111110111110000",
49587 => "0111110111110000",
49588 => "0111110111110000",
49589 => "0111110111110000",
49590 => "0111110111110000",
49591 => "0111110111110000",
49592 => "0111110111110000",
49593 => "0111110111110000",
49594 => "0111110111110000",
49595 => "0111110111110000",
49596 => "0111110111110000",
49597 => "0111110111110000",
49598 => "0111110111110000",
49599 => "0111110111110000",
49600 => "0111110111110000",
49601 => "0111110111110000",
49602 => "0111110111110000",
49603 => "0111110111110000",
49604 => "0111110111110000",
49605 => "0111110111110000",
49606 => "0111110111110000",
49607 => "0111110111110000",
49608 => "0111110111110000",
49609 => "0111110111110000",
49610 => "0111110111110000",
49611 => "0111110111110000",
49612 => "0111110111110000",
49613 => "0111110111110000",
49614 => "0111110111110000",
49615 => "0111110111110000",
49616 => "0111110111110000",
49617 => "0111110111110000",
49618 => "0111110111110000",
49619 => "0111110111110000",
49620 => "0111110111110000",
49621 => "0111110111110000",
49622 => "0111110111110000",
49623 => "0111110111110000",
49624 => "0111110111110000",
49625 => "0111110111110000",
49626 => "0111110111110000",
49627 => "0111110111110000",
49628 => "0111110111110000",
49629 => "0111110111110000",
49630 => "0111110111110000",
49631 => "0111110111110000",
49632 => "0111110111110000",
49633 => "0111110111110000",
49634 => "0111110111110000",
49635 => "0111110111110000",
49636 => "0111110111110000",
49637 => "0111110111110000",
49638 => "0111110111110000",
49639 => "0111110111110000",
49640 => "0111110111110000",
49641 => "0111110111110000",
49642 => "0111110111110000",
49643 => "0111110111110000",
49644 => "0111110111110000",
49645 => "0111110111110000",
49646 => "0111110111110000",
49647 => "0111110111110000",
49648 => "0111110111110000",
49649 => "0111110111110000",
49650 => "0111110111110000",
49651 => "0111110111110000",
49652 => "0111110111110000",
49653 => "0111110111110000",
49654 => "0111110111110000",
49655 => "0111110111110000",
49656 => "0111110111110000",
49657 => "0111110111110000",
49658 => "0111110111110000",
49659 => "0111110111110000",
49660 => "0111110111110000",
49661 => "0111110111110000",
49662 => "0111110111110000",
49663 => "0111110111110000",
49664 => "0111110111110000",
49665 => "0111110111110000",
49666 => "0111110111110000",
49667 => "0111110111110000",
49668 => "0111110111110000",
49669 => "0111110111110000",
49670 => "0111110111110000",
49671 => "0111110111110000",
49672 => "0111110111110000",
49673 => "0111110111110000",
49674 => "0111111000000000",
49675 => "0111111000000000",
49676 => "0111111000000000",
49677 => "0111111000000000",
49678 => "0111111000000000",
49679 => "0111111000000000",
49680 => "0111111000000000",
49681 => "0111111000000000",
49682 => "0111111000000000",
49683 => "0111111000000000",
49684 => "0111111000000000",
49685 => "0111111000000000",
49686 => "0111111000000000",
49687 => "0111111000000000",
49688 => "0111111000000000",
49689 => "0111111000000000",
49690 => "0111111000000000",
49691 => "0111111000000000",
49692 => "0111111000000000",
49693 => "0111111000000000",
49694 => "0111111000000000",
49695 => "0111111000000000",
49696 => "0111111000000000",
49697 => "0111111000000000",
49698 => "0111111000000000",
49699 => "0111111000000000",
49700 => "0111111000000000",
49701 => "0111111000000000",
49702 => "0111111000000000",
49703 => "0111111000000000",
49704 => "0111111000000000",
49705 => "0111111000000000",
49706 => "0111111000000000",
49707 => "0111111000000000",
49708 => "0111111000000000",
49709 => "0111111000000000",
49710 => "0111111000000000",
49711 => "0111111000000000",
49712 => "0111111000000000",
49713 => "0111111000000000",
49714 => "0111111000000000",
49715 => "0111111000000000",
49716 => "0111111000000000",
49717 => "0111111000000000",
49718 => "0111111000000000",
49719 => "0111111000000000",
49720 => "0111111000000000",
49721 => "0111111000000000",
49722 => "0111111000000000",
49723 => "0111111000000000",
49724 => "0111111000000000",
49725 => "0111111000000000",
49726 => "0111111000000000",
49727 => "0111111000000000",
49728 => "0111111000000000",
49729 => "0111111000000000",
49730 => "0111111000000000",
49731 => "0111111000000000",
49732 => "0111111000000000",
49733 => "0111111000000000",
49734 => "0111111000000000",
49735 => "0111111000000000",
49736 => "0111111000000000",
49737 => "0111111000000000",
49738 => "0111111000000000",
49739 => "0111111000000000",
49740 => "0111111000000000",
49741 => "0111111000000000",
49742 => "0111111000000000",
49743 => "0111111000000000",
49744 => "0111111000000000",
49745 => "0111111000000000",
49746 => "0111111000000000",
49747 => "0111111000000000",
49748 => "0111111000000000",
49749 => "0111111000000000",
49750 => "0111111000000000",
49751 => "0111111000000000",
49752 => "0111111000000000",
49753 => "0111111000000000",
49754 => "0111111000000000",
49755 => "0111111000000000",
49756 => "0111111000000000",
49757 => "0111111000000000",
49758 => "0111111000000000",
49759 => "0111111000000000",
49760 => "0111111000000000",
49761 => "0111111000000000",
49762 => "0111111000000000",
49763 => "0111111000000000",
49764 => "0111111000000000",
49765 => "0111111000000000",
49766 => "0111111000000000",
49767 => "0111111000000000",
49768 => "0111111000000000",
49769 => "0111111000000000",
49770 => "0111111000000000",
49771 => "0111111000000000",
49772 => "0111111000000000",
49773 => "0111111000000000",
49774 => "0111111000000000",
49775 => "0111111000000000",
49776 => "0111111000000000",
49777 => "0111111000000000",
49778 => "0111111000000000",
49779 => "0111111000000000",
49780 => "0111111000000000",
49781 => "0111111000000000",
49782 => "0111111000000000",
49783 => "0111111000000000",
49784 => "0111111000000000",
49785 => "0111111000000000",
49786 => "0111111000000000",
49787 => "0111111000000000",
49788 => "0111111000000000",
49789 => "0111111000000000",
49790 => "0111111000000000",
49791 => "0111111000000000",
49792 => "0111111000000000",
49793 => "0111111000000000",
49794 => "0111111000000000",
49795 => "0111111000000000",
49796 => "0111111000000000",
49797 => "0111111000000000",
49798 => "0111111000000000",
49799 => "0111111000000000",
49800 => "0111111000000000",
49801 => "0111111000000000",
49802 => "0111111000000000",
49803 => "0111111000000000",
49804 => "0111111000010000",
49805 => "0111111000010000",
49806 => "0111111000010000",
49807 => "0111111000010000",
49808 => "0111111000010000",
49809 => "0111111000010000",
49810 => "0111111000010000",
49811 => "0111111000010000",
49812 => "0111111000010000",
49813 => "0111111000010000",
49814 => "0111111000010000",
49815 => "0111111000010000",
49816 => "0111111000010000",
49817 => "0111111000010000",
49818 => "0111111000010000",
49819 => "0111111000010000",
49820 => "0111111000010000",
49821 => "0111111000010000",
49822 => "0111111000010000",
49823 => "0111111000010000",
49824 => "0111111000010000",
49825 => "0111111000010000",
49826 => "0111111000010000",
49827 => "0111111000010000",
49828 => "0111111000010000",
49829 => "0111111000010000",
49830 => "0111111000010000",
49831 => "0111111000010000",
49832 => "0111111000010000",
49833 => "0111111000010000",
49834 => "0111111000010000",
49835 => "0111111000010000",
49836 => "0111111000010000",
49837 => "0111111000010000",
49838 => "0111111000010000",
49839 => "0111111000010000",
49840 => "0111111000010000",
49841 => "0111111000010000",
49842 => "0111111000010000",
49843 => "0111111000010000",
49844 => "0111111000010000",
49845 => "0111111000010000",
49846 => "0111111000010000",
49847 => "0111111000010000",
49848 => "0111111000010000",
49849 => "0111111000010000",
49850 => "0111111000010000",
49851 => "0111111000010000",
49852 => "0111111000010000",
49853 => "0111111000010000",
49854 => "0111111000010000",
49855 => "0111111000010000",
49856 => "0111111000010000",
49857 => "0111111000010000",
49858 => "0111111000010000",
49859 => "0111111000010000",
49860 => "0111111000010000",
49861 => "0111111000010000",
49862 => "0111111000010000",
49863 => "0111111000010000",
49864 => "0111111000010000",
49865 => "0111111000010000",
49866 => "0111111000010000",
49867 => "0111111000010000",
49868 => "0111111000010000",
49869 => "0111111000010000",
49870 => "0111111000010000",
49871 => "0111111000010000",
49872 => "0111111000010000",
49873 => "0111111000010000",
49874 => "0111111000010000",
49875 => "0111111000010000",
49876 => "0111111000010000",
49877 => "0111111000010000",
49878 => "0111111000010000",
49879 => "0111111000010000",
49880 => "0111111000010000",
49881 => "0111111000010000",
49882 => "0111111000010000",
49883 => "0111111000010000",
49884 => "0111111000010000",
49885 => "0111111000010000",
49886 => "0111111000010000",
49887 => "0111111000010000",
49888 => "0111111000010000",
49889 => "0111111000010000",
49890 => "0111111000010000",
49891 => "0111111000010000",
49892 => "0111111000010000",
49893 => "0111111000010000",
49894 => "0111111000010000",
49895 => "0111111000010000",
49896 => "0111111000010000",
49897 => "0111111000010000",
49898 => "0111111000010000",
49899 => "0111111000010000",
49900 => "0111111000010000",
49901 => "0111111000010000",
49902 => "0111111000010000",
49903 => "0111111000010000",
49904 => "0111111000010000",
49905 => "0111111000010000",
49906 => "0111111000010000",
49907 => "0111111000010000",
49908 => "0111111000010000",
49909 => "0111111000010000",
49910 => "0111111000010000",
49911 => "0111111000010000",
49912 => "0111111000010000",
49913 => "0111111000010000",
49914 => "0111111000010000",
49915 => "0111111000010000",
49916 => "0111111000010000",
49917 => "0111111000010000",
49918 => "0111111000010000",
49919 => "0111111000010000",
49920 => "0111111000010000",
49921 => "0111111000010000",
49922 => "0111111000010000",
49923 => "0111111000010000",
49924 => "0111111000010000",
49925 => "0111111000010000",
49926 => "0111111000010000",
49927 => "0111111000010000",
49928 => "0111111000010000",
49929 => "0111111000010000",
49930 => "0111111000010000",
49931 => "0111111000010000",
49932 => "0111111000010000",
49933 => "0111111000010000",
49934 => "0111111000010000",
49935 => "0111111000010000",
49936 => "0111111000010000",
49937 => "0111111000010000",
49938 => "0111111000100000",
49939 => "0111111000100000",
49940 => "0111111000100000",
49941 => "0111111000100000",
49942 => "0111111000100000",
49943 => "0111111000100000",
49944 => "0111111000100000",
49945 => "0111111000100000",
49946 => "0111111000100000",
49947 => "0111111000100000",
49948 => "0111111000100000",
49949 => "0111111000100000",
49950 => "0111111000100000",
49951 => "0111111000100000",
49952 => "0111111000100000",
49953 => "0111111000100000",
49954 => "0111111000100000",
49955 => "0111111000100000",
49956 => "0111111000100000",
49957 => "0111111000100000",
49958 => "0111111000100000",
49959 => "0111111000100000",
49960 => "0111111000100000",
49961 => "0111111000100000",
49962 => "0111111000100000",
49963 => "0111111000100000",
49964 => "0111111000100000",
49965 => "0111111000100000",
49966 => "0111111000100000",
49967 => "0111111000100000",
49968 => "0111111000100000",
49969 => "0111111000100000",
49970 => "0111111000100000",
49971 => "0111111000100000",
49972 => "0111111000100000",
49973 => "0111111000100000",
49974 => "0111111000100000",
49975 => "0111111000100000",
49976 => "0111111000100000",
49977 => "0111111000100000",
49978 => "0111111000100000",
49979 => "0111111000100000",
49980 => "0111111000100000",
49981 => "0111111000100000",
49982 => "0111111000100000",
49983 => "0111111000100000",
49984 => "0111111000100000",
49985 => "0111111000100000",
49986 => "0111111000100000",
49987 => "0111111000100000",
49988 => "0111111000100000",
49989 => "0111111000100000",
49990 => "0111111000100000",
49991 => "0111111000100000",
49992 => "0111111000100000",
49993 => "0111111000100000",
49994 => "0111111000100000",
49995 => "0111111000100000",
49996 => "0111111000100000",
49997 => "0111111000100000",
49998 => "0111111000100000",
49999 => "0111111000100000",
50000 => "0111111000100000",
50001 => "0111111000100000",
50002 => "0111111000100000",
50003 => "0111111000100000",
50004 => "0111111000100000",
50005 => "0111111000100000",
50006 => "0111111000100000",
50007 => "0111111000100000",
50008 => "0111111000100000",
50009 => "0111111000100000",
50010 => "0111111000100000",
50011 => "0111111000100000",
50012 => "0111111000100000",
50013 => "0111111000100000",
50014 => "0111111000100000",
50015 => "0111111000100000",
50016 => "0111111000100000",
50017 => "0111111000100000",
50018 => "0111111000100000",
50019 => "0111111000100000",
50020 => "0111111000100000",
50021 => "0111111000100000",
50022 => "0111111000100000",
50023 => "0111111000100000",
50024 => "0111111000100000",
50025 => "0111111000100000",
50026 => "0111111000100000",
50027 => "0111111000100000",
50028 => "0111111000100000",
50029 => "0111111000100000",
50030 => "0111111000100000",
50031 => "0111111000100000",
50032 => "0111111000100000",
50033 => "0111111000100000",
50034 => "0111111000100000",
50035 => "0111111000100000",
50036 => "0111111000100000",
50037 => "0111111000100000",
50038 => "0111111000100000",
50039 => "0111111000100000",
50040 => "0111111000100000",
50041 => "0111111000100000",
50042 => "0111111000100000",
50043 => "0111111000100000",
50044 => "0111111000100000",
50045 => "0111111000100000",
50046 => "0111111000100000",
50047 => "0111111000100000",
50048 => "0111111000100000",
50049 => "0111111000100000",
50050 => "0111111000100000",
50051 => "0111111000100000",
50052 => "0111111000100000",
50053 => "0111111000100000",
50054 => "0111111000100000",
50055 => "0111111000100000",
50056 => "0111111000100000",
50057 => "0111111000100000",
50058 => "0111111000100000",
50059 => "0111111000100000",
50060 => "0111111000100000",
50061 => "0111111000100000",
50062 => "0111111000100000",
50063 => "0111111000100000",
50064 => "0111111000100000",
50065 => "0111111000100000",
50066 => "0111111000100000",
50067 => "0111111000100000",
50068 => "0111111000100000",
50069 => "0111111000100000",
50070 => "0111111000100000",
50071 => "0111111000100000",
50072 => "0111111000100000",
50073 => "0111111000100000",
50074 => "0111111000100000",
50075 => "0111111000100000",
50076 => "0111111000110000",
50077 => "0111111000110000",
50078 => "0111111000110000",
50079 => "0111111000110000",
50080 => "0111111000110000",
50081 => "0111111000110000",
50082 => "0111111000110000",
50083 => "0111111000110000",
50084 => "0111111000110000",
50085 => "0111111000110000",
50086 => "0111111000110000",
50087 => "0111111000110000",
50088 => "0111111000110000",
50089 => "0111111000110000",
50090 => "0111111000110000",
50091 => "0111111000110000",
50092 => "0111111000110000",
50093 => "0111111000110000",
50094 => "0111111000110000",
50095 => "0111111000110000",
50096 => "0111111000110000",
50097 => "0111111000110000",
50098 => "0111111000110000",
50099 => "0111111000110000",
50100 => "0111111000110000",
50101 => "0111111000110000",
50102 => "0111111000110000",
50103 => "0111111000110000",
50104 => "0111111000110000",
50105 => "0111111000110000",
50106 => "0111111000110000",
50107 => "0111111000110000",
50108 => "0111111000110000",
50109 => "0111111000110000",
50110 => "0111111000110000",
50111 => "0111111000110000",
50112 => "0111111000110000",
50113 => "0111111000110000",
50114 => "0111111000110000",
50115 => "0111111000110000",
50116 => "0111111000110000",
50117 => "0111111000110000",
50118 => "0111111000110000",
50119 => "0111111000110000",
50120 => "0111111000110000",
50121 => "0111111000110000",
50122 => "0111111000110000",
50123 => "0111111000110000",
50124 => "0111111000110000",
50125 => "0111111000110000",
50126 => "0111111000110000",
50127 => "0111111000110000",
50128 => "0111111000110000",
50129 => "0111111000110000",
50130 => "0111111000110000",
50131 => "0111111000110000",
50132 => "0111111000110000",
50133 => "0111111000110000",
50134 => "0111111000110000",
50135 => "0111111000110000",
50136 => "0111111000110000",
50137 => "0111111000110000",
50138 => "0111111000110000",
50139 => "0111111000110000",
50140 => "0111111000110000",
50141 => "0111111000110000",
50142 => "0111111000110000",
50143 => "0111111000110000",
50144 => "0111111000110000",
50145 => "0111111000110000",
50146 => "0111111000110000",
50147 => "0111111000110000",
50148 => "0111111000110000",
50149 => "0111111000110000",
50150 => "0111111000110000",
50151 => "0111111000110000",
50152 => "0111111000110000",
50153 => "0111111000110000",
50154 => "0111111000110000",
50155 => "0111111000110000",
50156 => "0111111000110000",
50157 => "0111111000110000",
50158 => "0111111000110000",
50159 => "0111111000110000",
50160 => "0111111000110000",
50161 => "0111111000110000",
50162 => "0111111000110000",
50163 => "0111111000110000",
50164 => "0111111000110000",
50165 => "0111111000110000",
50166 => "0111111000110000",
50167 => "0111111000110000",
50168 => "0111111000110000",
50169 => "0111111000110000",
50170 => "0111111000110000",
50171 => "0111111000110000",
50172 => "0111111000110000",
50173 => "0111111000110000",
50174 => "0111111000110000",
50175 => "0111111000110000",
50176 => "0111111000110000",
50177 => "0111111000110000",
50178 => "0111111000110000",
50179 => "0111111000110000",
50180 => "0111111000110000",
50181 => "0111111000110000",
50182 => "0111111000110000",
50183 => "0111111000110000",
50184 => "0111111000110000",
50185 => "0111111000110000",
50186 => "0111111000110000",
50187 => "0111111000110000",
50188 => "0111111000110000",
50189 => "0111111000110000",
50190 => "0111111000110000",
50191 => "0111111000110000",
50192 => "0111111000110000",
50193 => "0111111000110000",
50194 => "0111111000110000",
50195 => "0111111000110000",
50196 => "0111111000110000",
50197 => "0111111000110000",
50198 => "0111111000110000",
50199 => "0111111000110000",
50200 => "0111111000110000",
50201 => "0111111000110000",
50202 => "0111111000110000",
50203 => "0111111000110000",
50204 => "0111111000110000",
50205 => "0111111000110000",
50206 => "0111111000110000",
50207 => "0111111000110000",
50208 => "0111111000110000",
50209 => "0111111000110000",
50210 => "0111111000110000",
50211 => "0111111000110000",
50212 => "0111111000110000",
50213 => "0111111000110000",
50214 => "0111111000110000",
50215 => "0111111000110000",
50216 => "0111111000110000",
50217 => "0111111000110000",
50218 => "0111111000110000",
50219 => "0111111000110000",
50220 => "0111111001000000",
50221 => "0111111001000000",
50222 => "0111111001000000",
50223 => "0111111001000000",
50224 => "0111111001000000",
50225 => "0111111001000000",
50226 => "0111111001000000",
50227 => "0111111001000000",
50228 => "0111111001000000",
50229 => "0111111001000000",
50230 => "0111111001000000",
50231 => "0111111001000000",
50232 => "0111111001000000",
50233 => "0111111001000000",
50234 => "0111111001000000",
50235 => "0111111001000000",
50236 => "0111111001000000",
50237 => "0111111001000000",
50238 => "0111111001000000",
50239 => "0111111001000000",
50240 => "0111111001000000",
50241 => "0111111001000000",
50242 => "0111111001000000",
50243 => "0111111001000000",
50244 => "0111111001000000",
50245 => "0111111001000000",
50246 => "0111111001000000",
50247 => "0111111001000000",
50248 => "0111111001000000",
50249 => "0111111001000000",
50250 => "0111111001000000",
50251 => "0111111001000000",
50252 => "0111111001000000",
50253 => "0111111001000000",
50254 => "0111111001000000",
50255 => "0111111001000000",
50256 => "0111111001000000",
50257 => "0111111001000000",
50258 => "0111111001000000",
50259 => "0111111001000000",
50260 => "0111111001000000",
50261 => "0111111001000000",
50262 => "0111111001000000",
50263 => "0111111001000000",
50264 => "0111111001000000",
50265 => "0111111001000000",
50266 => "0111111001000000",
50267 => "0111111001000000",
50268 => "0111111001000000",
50269 => "0111111001000000",
50270 => "0111111001000000",
50271 => "0111111001000000",
50272 => "0111111001000000",
50273 => "0111111001000000",
50274 => "0111111001000000",
50275 => "0111111001000000",
50276 => "0111111001000000",
50277 => "0111111001000000",
50278 => "0111111001000000",
50279 => "0111111001000000",
50280 => "0111111001000000",
50281 => "0111111001000000",
50282 => "0111111001000000",
50283 => "0111111001000000",
50284 => "0111111001000000",
50285 => "0111111001000000",
50286 => "0111111001000000",
50287 => "0111111001000000",
50288 => "0111111001000000",
50289 => "0111111001000000",
50290 => "0111111001000000",
50291 => "0111111001000000",
50292 => "0111111001000000",
50293 => "0111111001000000",
50294 => "0111111001000000",
50295 => "0111111001000000",
50296 => "0111111001000000",
50297 => "0111111001000000",
50298 => "0111111001000000",
50299 => "0111111001000000",
50300 => "0111111001000000",
50301 => "0111111001000000",
50302 => "0111111001000000",
50303 => "0111111001000000",
50304 => "0111111001000000",
50305 => "0111111001000000",
50306 => "0111111001000000",
50307 => "0111111001000000",
50308 => "0111111001000000",
50309 => "0111111001000000",
50310 => "0111111001000000",
50311 => "0111111001000000",
50312 => "0111111001000000",
50313 => "0111111001000000",
50314 => "0111111001000000",
50315 => "0111111001000000",
50316 => "0111111001000000",
50317 => "0111111001000000",
50318 => "0111111001000000",
50319 => "0111111001000000",
50320 => "0111111001000000",
50321 => "0111111001000000",
50322 => "0111111001000000",
50323 => "0111111001000000",
50324 => "0111111001000000",
50325 => "0111111001000000",
50326 => "0111111001000000",
50327 => "0111111001000000",
50328 => "0111111001000000",
50329 => "0111111001000000",
50330 => "0111111001000000",
50331 => "0111111001000000",
50332 => "0111111001000000",
50333 => "0111111001000000",
50334 => "0111111001000000",
50335 => "0111111001000000",
50336 => "0111111001000000",
50337 => "0111111001000000",
50338 => "0111111001000000",
50339 => "0111111001000000",
50340 => "0111111001000000",
50341 => "0111111001000000",
50342 => "0111111001000000",
50343 => "0111111001000000",
50344 => "0111111001000000",
50345 => "0111111001000000",
50346 => "0111111001000000",
50347 => "0111111001000000",
50348 => "0111111001000000",
50349 => "0111111001000000",
50350 => "0111111001000000",
50351 => "0111111001000000",
50352 => "0111111001000000",
50353 => "0111111001000000",
50354 => "0111111001000000",
50355 => "0111111001000000",
50356 => "0111111001000000",
50357 => "0111111001000000",
50358 => "0111111001000000",
50359 => "0111111001000000",
50360 => "0111111001000000",
50361 => "0111111001000000",
50362 => "0111111001000000",
50363 => "0111111001000000",
50364 => "0111111001000000",
50365 => "0111111001000000",
50366 => "0111111001000000",
50367 => "0111111001000000",
50368 => "0111111001010000",
50369 => "0111111001010000",
50370 => "0111111001010000",
50371 => "0111111001010000",
50372 => "0111111001010000",
50373 => "0111111001010000",
50374 => "0111111001010000",
50375 => "0111111001010000",
50376 => "0111111001010000",
50377 => "0111111001010000",
50378 => "0111111001010000",
50379 => "0111111001010000",
50380 => "0111111001010000",
50381 => "0111111001010000",
50382 => "0111111001010000",
50383 => "0111111001010000",
50384 => "0111111001010000",
50385 => "0111111001010000",
50386 => "0111111001010000",
50387 => "0111111001010000",
50388 => "0111111001010000",
50389 => "0111111001010000",
50390 => "0111111001010000",
50391 => "0111111001010000",
50392 => "0111111001010000",
50393 => "0111111001010000",
50394 => "0111111001010000",
50395 => "0111111001010000",
50396 => "0111111001010000",
50397 => "0111111001010000",
50398 => "0111111001010000",
50399 => "0111111001010000",
50400 => "0111111001010000",
50401 => "0111111001010000",
50402 => "0111111001010000",
50403 => "0111111001010000",
50404 => "0111111001010000",
50405 => "0111111001010000",
50406 => "0111111001010000",
50407 => "0111111001010000",
50408 => "0111111001010000",
50409 => "0111111001010000",
50410 => "0111111001010000",
50411 => "0111111001010000",
50412 => "0111111001010000",
50413 => "0111111001010000",
50414 => "0111111001010000",
50415 => "0111111001010000",
50416 => "0111111001010000",
50417 => "0111111001010000",
50418 => "0111111001010000",
50419 => "0111111001010000",
50420 => "0111111001010000",
50421 => "0111111001010000",
50422 => "0111111001010000",
50423 => "0111111001010000",
50424 => "0111111001010000",
50425 => "0111111001010000",
50426 => "0111111001010000",
50427 => "0111111001010000",
50428 => "0111111001010000",
50429 => "0111111001010000",
50430 => "0111111001010000",
50431 => "0111111001010000",
50432 => "0111111001010000",
50433 => "0111111001010000",
50434 => "0111111001010000",
50435 => "0111111001010000",
50436 => "0111111001010000",
50437 => "0111111001010000",
50438 => "0111111001010000",
50439 => "0111111001010000",
50440 => "0111111001010000",
50441 => "0111111001010000",
50442 => "0111111001010000",
50443 => "0111111001010000",
50444 => "0111111001010000",
50445 => "0111111001010000",
50446 => "0111111001010000",
50447 => "0111111001010000",
50448 => "0111111001010000",
50449 => "0111111001010000",
50450 => "0111111001010000",
50451 => "0111111001010000",
50452 => "0111111001010000",
50453 => "0111111001010000",
50454 => "0111111001010000",
50455 => "0111111001010000",
50456 => "0111111001010000",
50457 => "0111111001010000",
50458 => "0111111001010000",
50459 => "0111111001010000",
50460 => "0111111001010000",
50461 => "0111111001010000",
50462 => "0111111001010000",
50463 => "0111111001010000",
50464 => "0111111001010000",
50465 => "0111111001010000",
50466 => "0111111001010000",
50467 => "0111111001010000",
50468 => "0111111001010000",
50469 => "0111111001010000",
50470 => "0111111001010000",
50471 => "0111111001010000",
50472 => "0111111001010000",
50473 => "0111111001010000",
50474 => "0111111001010000",
50475 => "0111111001010000",
50476 => "0111111001010000",
50477 => "0111111001010000",
50478 => "0111111001010000",
50479 => "0111111001010000",
50480 => "0111111001010000",
50481 => "0111111001010000",
50482 => "0111111001010000",
50483 => "0111111001010000",
50484 => "0111111001010000",
50485 => "0111111001010000",
50486 => "0111111001010000",
50487 => "0111111001010000",
50488 => "0111111001010000",
50489 => "0111111001010000",
50490 => "0111111001010000",
50491 => "0111111001010000",
50492 => "0111111001010000",
50493 => "0111111001010000",
50494 => "0111111001010000",
50495 => "0111111001010000",
50496 => "0111111001010000",
50497 => "0111111001010000",
50498 => "0111111001010000",
50499 => "0111111001010000",
50500 => "0111111001010000",
50501 => "0111111001010000",
50502 => "0111111001010000",
50503 => "0111111001010000",
50504 => "0111111001010000",
50505 => "0111111001010000",
50506 => "0111111001010000",
50507 => "0111111001010000",
50508 => "0111111001010000",
50509 => "0111111001010000",
50510 => "0111111001010000",
50511 => "0111111001010000",
50512 => "0111111001010000",
50513 => "0111111001010000",
50514 => "0111111001010000",
50515 => "0111111001010000",
50516 => "0111111001010000",
50517 => "0111111001010000",
50518 => "0111111001010000",
50519 => "0111111001010000",
50520 => "0111111001010000",
50521 => "0111111001010000",
50522 => "0111111001100000",
50523 => "0111111001100000",
50524 => "0111111001100000",
50525 => "0111111001100000",
50526 => "0111111001100000",
50527 => "0111111001100000",
50528 => "0111111001100000",
50529 => "0111111001100000",
50530 => "0111111001100000",
50531 => "0111111001100000",
50532 => "0111111001100000",
50533 => "0111111001100000",
50534 => "0111111001100000",
50535 => "0111111001100000",
50536 => "0111111001100000",
50537 => "0111111001100000",
50538 => "0111111001100000",
50539 => "0111111001100000",
50540 => "0111111001100000",
50541 => "0111111001100000",
50542 => "0111111001100000",
50543 => "0111111001100000",
50544 => "0111111001100000",
50545 => "0111111001100000",
50546 => "0111111001100000",
50547 => "0111111001100000",
50548 => "0111111001100000",
50549 => "0111111001100000",
50550 => "0111111001100000",
50551 => "0111111001100000",
50552 => "0111111001100000",
50553 => "0111111001100000",
50554 => "0111111001100000",
50555 => "0111111001100000",
50556 => "0111111001100000",
50557 => "0111111001100000",
50558 => "0111111001100000",
50559 => "0111111001100000",
50560 => "0111111001100000",
50561 => "0111111001100000",
50562 => "0111111001100000",
50563 => "0111111001100000",
50564 => "0111111001100000",
50565 => "0111111001100000",
50566 => "0111111001100000",
50567 => "0111111001100000",
50568 => "0111111001100000",
50569 => "0111111001100000",
50570 => "0111111001100000",
50571 => "0111111001100000",
50572 => "0111111001100000",
50573 => "0111111001100000",
50574 => "0111111001100000",
50575 => "0111111001100000",
50576 => "0111111001100000",
50577 => "0111111001100000",
50578 => "0111111001100000",
50579 => "0111111001100000",
50580 => "0111111001100000",
50581 => "0111111001100000",
50582 => "0111111001100000",
50583 => "0111111001100000",
50584 => "0111111001100000",
50585 => "0111111001100000",
50586 => "0111111001100000",
50587 => "0111111001100000",
50588 => "0111111001100000",
50589 => "0111111001100000",
50590 => "0111111001100000",
50591 => "0111111001100000",
50592 => "0111111001100000",
50593 => "0111111001100000",
50594 => "0111111001100000",
50595 => "0111111001100000",
50596 => "0111111001100000",
50597 => "0111111001100000",
50598 => "0111111001100000",
50599 => "0111111001100000",
50600 => "0111111001100000",
50601 => "0111111001100000",
50602 => "0111111001100000",
50603 => "0111111001100000",
50604 => "0111111001100000",
50605 => "0111111001100000",
50606 => "0111111001100000",
50607 => "0111111001100000",
50608 => "0111111001100000",
50609 => "0111111001100000",
50610 => "0111111001100000",
50611 => "0111111001100000",
50612 => "0111111001100000",
50613 => "0111111001100000",
50614 => "0111111001100000",
50615 => "0111111001100000",
50616 => "0111111001100000",
50617 => "0111111001100000",
50618 => "0111111001100000",
50619 => "0111111001100000",
50620 => "0111111001100000",
50621 => "0111111001100000",
50622 => "0111111001100000",
50623 => "0111111001100000",
50624 => "0111111001100000",
50625 => "0111111001100000",
50626 => "0111111001100000",
50627 => "0111111001100000",
50628 => "0111111001100000",
50629 => "0111111001100000",
50630 => "0111111001100000",
50631 => "0111111001100000",
50632 => "0111111001100000",
50633 => "0111111001100000",
50634 => "0111111001100000",
50635 => "0111111001100000",
50636 => "0111111001100000",
50637 => "0111111001100000",
50638 => "0111111001100000",
50639 => "0111111001100000",
50640 => "0111111001100000",
50641 => "0111111001100000",
50642 => "0111111001100000",
50643 => "0111111001100000",
50644 => "0111111001100000",
50645 => "0111111001100000",
50646 => "0111111001100000",
50647 => "0111111001100000",
50648 => "0111111001100000",
50649 => "0111111001100000",
50650 => "0111111001100000",
50651 => "0111111001100000",
50652 => "0111111001100000",
50653 => "0111111001100000",
50654 => "0111111001100000",
50655 => "0111111001100000",
50656 => "0111111001100000",
50657 => "0111111001100000",
50658 => "0111111001100000",
50659 => "0111111001100000",
50660 => "0111111001100000",
50661 => "0111111001100000",
50662 => "0111111001100000",
50663 => "0111111001100000",
50664 => "0111111001100000",
50665 => "0111111001100000",
50666 => "0111111001100000",
50667 => "0111111001100000",
50668 => "0111111001100000",
50669 => "0111111001100000",
50670 => "0111111001100000",
50671 => "0111111001100000",
50672 => "0111111001100000",
50673 => "0111111001100000",
50674 => "0111111001100000",
50675 => "0111111001100000",
50676 => "0111111001100000",
50677 => "0111111001100000",
50678 => "0111111001100000",
50679 => "0111111001100000",
50680 => "0111111001100000",
50681 => "0111111001110000",
50682 => "0111111001110000",
50683 => "0111111001110000",
50684 => "0111111001110000",
50685 => "0111111001110000",
50686 => "0111111001110000",
50687 => "0111111001110000",
50688 => "0111111001110000",
50689 => "0111111001110000",
50690 => "0111111001110000",
50691 => "0111111001110000",
50692 => "0111111001110000",
50693 => "0111111001110000",
50694 => "0111111001110000",
50695 => "0111111001110000",
50696 => "0111111001110000",
50697 => "0111111001110000",
50698 => "0111111001110000",
50699 => "0111111001110000",
50700 => "0111111001110000",
50701 => "0111111001110000",
50702 => "0111111001110000",
50703 => "0111111001110000",
50704 => "0111111001110000",
50705 => "0111111001110000",
50706 => "0111111001110000",
50707 => "0111111001110000",
50708 => "0111111001110000",
50709 => "0111111001110000",
50710 => "0111111001110000",
50711 => "0111111001110000",
50712 => "0111111001110000",
50713 => "0111111001110000",
50714 => "0111111001110000",
50715 => "0111111001110000",
50716 => "0111111001110000",
50717 => "0111111001110000",
50718 => "0111111001110000",
50719 => "0111111001110000",
50720 => "0111111001110000",
50721 => "0111111001110000",
50722 => "0111111001110000",
50723 => "0111111001110000",
50724 => "0111111001110000",
50725 => "0111111001110000",
50726 => "0111111001110000",
50727 => "0111111001110000",
50728 => "0111111001110000",
50729 => "0111111001110000",
50730 => "0111111001110000",
50731 => "0111111001110000",
50732 => "0111111001110000",
50733 => "0111111001110000",
50734 => "0111111001110000",
50735 => "0111111001110000",
50736 => "0111111001110000",
50737 => "0111111001110000",
50738 => "0111111001110000",
50739 => "0111111001110000",
50740 => "0111111001110000",
50741 => "0111111001110000",
50742 => "0111111001110000",
50743 => "0111111001110000",
50744 => "0111111001110000",
50745 => "0111111001110000",
50746 => "0111111001110000",
50747 => "0111111001110000",
50748 => "0111111001110000",
50749 => "0111111001110000",
50750 => "0111111001110000",
50751 => "0111111001110000",
50752 => "0111111001110000",
50753 => "0111111001110000",
50754 => "0111111001110000",
50755 => "0111111001110000",
50756 => "0111111001110000",
50757 => "0111111001110000",
50758 => "0111111001110000",
50759 => "0111111001110000",
50760 => "0111111001110000",
50761 => "0111111001110000",
50762 => "0111111001110000",
50763 => "0111111001110000",
50764 => "0111111001110000",
50765 => "0111111001110000",
50766 => "0111111001110000",
50767 => "0111111001110000",
50768 => "0111111001110000",
50769 => "0111111001110000",
50770 => "0111111001110000",
50771 => "0111111001110000",
50772 => "0111111001110000",
50773 => "0111111001110000",
50774 => "0111111001110000",
50775 => "0111111001110000",
50776 => "0111111001110000",
50777 => "0111111001110000",
50778 => "0111111001110000",
50779 => "0111111001110000",
50780 => "0111111001110000",
50781 => "0111111001110000",
50782 => "0111111001110000",
50783 => "0111111001110000",
50784 => "0111111001110000",
50785 => "0111111001110000",
50786 => "0111111001110000",
50787 => "0111111001110000",
50788 => "0111111001110000",
50789 => "0111111001110000",
50790 => "0111111001110000",
50791 => "0111111001110000",
50792 => "0111111001110000",
50793 => "0111111001110000",
50794 => "0111111001110000",
50795 => "0111111001110000",
50796 => "0111111001110000",
50797 => "0111111001110000",
50798 => "0111111001110000",
50799 => "0111111001110000",
50800 => "0111111001110000",
50801 => "0111111001110000",
50802 => "0111111001110000",
50803 => "0111111001110000",
50804 => "0111111001110000",
50805 => "0111111001110000",
50806 => "0111111001110000",
50807 => "0111111001110000",
50808 => "0111111001110000",
50809 => "0111111001110000",
50810 => "0111111001110000",
50811 => "0111111001110000",
50812 => "0111111001110000",
50813 => "0111111001110000",
50814 => "0111111001110000",
50815 => "0111111001110000",
50816 => "0111111001110000",
50817 => "0111111001110000",
50818 => "0111111001110000",
50819 => "0111111001110000",
50820 => "0111111001110000",
50821 => "0111111001110000",
50822 => "0111111001110000",
50823 => "0111111001110000",
50824 => "0111111001110000",
50825 => "0111111001110000",
50826 => "0111111001110000",
50827 => "0111111001110000",
50828 => "0111111001110000",
50829 => "0111111001110000",
50830 => "0111111001110000",
50831 => "0111111001110000",
50832 => "0111111001110000",
50833 => "0111111001110000",
50834 => "0111111001110000",
50835 => "0111111001110000",
50836 => "0111111001110000",
50837 => "0111111001110000",
50838 => "0111111001110000",
50839 => "0111111001110000",
50840 => "0111111001110000",
50841 => "0111111001110000",
50842 => "0111111001110000",
50843 => "0111111001110000",
50844 => "0111111001110000",
50845 => "0111111001110000",
50846 => "0111111001110000",
50847 => "0111111010000000",
50848 => "0111111010000000",
50849 => "0111111010000000",
50850 => "0111111010000000",
50851 => "0111111010000000",
50852 => "0111111010000000",
50853 => "0111111010000000",
50854 => "0111111010000000",
50855 => "0111111010000000",
50856 => "0111111010000000",
50857 => "0111111010000000",
50858 => "0111111010000000",
50859 => "0111111010000000",
50860 => "0111111010000000",
50861 => "0111111010000000",
50862 => "0111111010000000",
50863 => "0111111010000000",
50864 => "0111111010000000",
50865 => "0111111010000000",
50866 => "0111111010000000",
50867 => "0111111010000000",
50868 => "0111111010000000",
50869 => "0111111010000000",
50870 => "0111111010000000",
50871 => "0111111010000000",
50872 => "0111111010000000",
50873 => "0111111010000000",
50874 => "0111111010000000",
50875 => "0111111010000000",
50876 => "0111111010000000",
50877 => "0111111010000000",
50878 => "0111111010000000",
50879 => "0111111010000000",
50880 => "0111111010000000",
50881 => "0111111010000000",
50882 => "0111111010000000",
50883 => "0111111010000000",
50884 => "0111111010000000",
50885 => "0111111010000000",
50886 => "0111111010000000",
50887 => "0111111010000000",
50888 => "0111111010000000",
50889 => "0111111010000000",
50890 => "0111111010000000",
50891 => "0111111010000000",
50892 => "0111111010000000",
50893 => "0111111010000000",
50894 => "0111111010000000",
50895 => "0111111010000000",
50896 => "0111111010000000",
50897 => "0111111010000000",
50898 => "0111111010000000",
50899 => "0111111010000000",
50900 => "0111111010000000",
50901 => "0111111010000000",
50902 => "0111111010000000",
50903 => "0111111010000000",
50904 => "0111111010000000",
50905 => "0111111010000000",
50906 => "0111111010000000",
50907 => "0111111010000000",
50908 => "0111111010000000",
50909 => "0111111010000000",
50910 => "0111111010000000",
50911 => "0111111010000000",
50912 => "0111111010000000",
50913 => "0111111010000000",
50914 => "0111111010000000",
50915 => "0111111010000000",
50916 => "0111111010000000",
50917 => "0111111010000000",
50918 => "0111111010000000",
50919 => "0111111010000000",
50920 => "0111111010000000",
50921 => "0111111010000000",
50922 => "0111111010000000",
50923 => "0111111010000000",
50924 => "0111111010000000",
50925 => "0111111010000000",
50926 => "0111111010000000",
50927 => "0111111010000000",
50928 => "0111111010000000",
50929 => "0111111010000000",
50930 => "0111111010000000",
50931 => "0111111010000000",
50932 => "0111111010000000",
50933 => "0111111010000000",
50934 => "0111111010000000",
50935 => "0111111010000000",
50936 => "0111111010000000",
50937 => "0111111010000000",
50938 => "0111111010000000",
50939 => "0111111010000000",
50940 => "0111111010000000",
50941 => "0111111010000000",
50942 => "0111111010000000",
50943 => "0111111010000000",
50944 => "0111111010000000",
50945 => "0111111010000000",
50946 => "0111111010000000",
50947 => "0111111010000000",
50948 => "0111111010000000",
50949 => "0111111010000000",
50950 => "0111111010000000",
50951 => "0111111010000000",
50952 => "0111111010000000",
50953 => "0111111010000000",
50954 => "0111111010000000",
50955 => "0111111010000000",
50956 => "0111111010000000",
50957 => "0111111010000000",
50958 => "0111111010000000",
50959 => "0111111010000000",
50960 => "0111111010000000",
50961 => "0111111010000000",
50962 => "0111111010000000",
50963 => "0111111010000000",
50964 => "0111111010000000",
50965 => "0111111010000000",
50966 => "0111111010000000",
50967 => "0111111010000000",
50968 => "0111111010000000",
50969 => "0111111010000000",
50970 => "0111111010000000",
50971 => "0111111010000000",
50972 => "0111111010000000",
50973 => "0111111010000000",
50974 => "0111111010000000",
50975 => "0111111010000000",
50976 => "0111111010000000",
50977 => "0111111010000000",
50978 => "0111111010000000",
50979 => "0111111010000000",
50980 => "0111111010000000",
50981 => "0111111010000000",
50982 => "0111111010000000",
50983 => "0111111010000000",
50984 => "0111111010000000",
50985 => "0111111010000000",
50986 => "0111111010000000",
50987 => "0111111010000000",
50988 => "0111111010000000",
50989 => "0111111010000000",
50990 => "0111111010000000",
50991 => "0111111010000000",
50992 => "0111111010000000",
50993 => "0111111010000000",
50994 => "0111111010000000",
50995 => "0111111010000000",
50996 => "0111111010000000",
50997 => "0111111010000000",
50998 => "0111111010000000",
50999 => "0111111010000000",
51000 => "0111111010000000",
51001 => "0111111010000000",
51002 => "0111111010000000",
51003 => "0111111010000000",
51004 => "0111111010000000",
51005 => "0111111010000000",
51006 => "0111111010000000",
51007 => "0111111010000000",
51008 => "0111111010000000",
51009 => "0111111010000000",
51010 => "0111111010000000",
51011 => "0111111010000000",
51012 => "0111111010000000",
51013 => "0111111010000000",
51014 => "0111111010000000",
51015 => "0111111010000000",
51016 => "0111111010000000",
51017 => "0111111010000000",
51018 => "0111111010000000",
51019 => "0111111010000000",
51020 => "0111111010010000",
51021 => "0111111010010000",
51022 => "0111111010010000",
51023 => "0111111010010000",
51024 => "0111111010010000",
51025 => "0111111010010000",
51026 => "0111111010010000",
51027 => "0111111010010000",
51028 => "0111111010010000",
51029 => "0111111010010000",
51030 => "0111111010010000",
51031 => "0111111010010000",
51032 => "0111111010010000",
51033 => "0111111010010000",
51034 => "0111111010010000",
51035 => "0111111010010000",
51036 => "0111111010010000",
51037 => "0111111010010000",
51038 => "0111111010010000",
51039 => "0111111010010000",
51040 => "0111111010010000",
51041 => "0111111010010000",
51042 => "0111111010010000",
51043 => "0111111010010000",
51044 => "0111111010010000",
51045 => "0111111010010000",
51046 => "0111111010010000",
51047 => "0111111010010000",
51048 => "0111111010010000",
51049 => "0111111010010000",
51050 => "0111111010010000",
51051 => "0111111010010000",
51052 => "0111111010010000",
51053 => "0111111010010000",
51054 => "0111111010010000",
51055 => "0111111010010000",
51056 => "0111111010010000",
51057 => "0111111010010000",
51058 => "0111111010010000",
51059 => "0111111010010000",
51060 => "0111111010010000",
51061 => "0111111010010000",
51062 => "0111111010010000",
51063 => "0111111010010000",
51064 => "0111111010010000",
51065 => "0111111010010000",
51066 => "0111111010010000",
51067 => "0111111010010000",
51068 => "0111111010010000",
51069 => "0111111010010000",
51070 => "0111111010010000",
51071 => "0111111010010000",
51072 => "0111111010010000",
51073 => "0111111010010000",
51074 => "0111111010010000",
51075 => "0111111010010000",
51076 => "0111111010010000",
51077 => "0111111010010000",
51078 => "0111111010010000",
51079 => "0111111010010000",
51080 => "0111111010010000",
51081 => "0111111010010000",
51082 => "0111111010010000",
51083 => "0111111010010000",
51084 => "0111111010010000",
51085 => "0111111010010000",
51086 => "0111111010010000",
51087 => "0111111010010000",
51088 => "0111111010010000",
51089 => "0111111010010000",
51090 => "0111111010010000",
51091 => "0111111010010000",
51092 => "0111111010010000",
51093 => "0111111010010000",
51094 => "0111111010010000",
51095 => "0111111010010000",
51096 => "0111111010010000",
51097 => "0111111010010000",
51098 => "0111111010010000",
51099 => "0111111010010000",
51100 => "0111111010010000",
51101 => "0111111010010000",
51102 => "0111111010010000",
51103 => "0111111010010000",
51104 => "0111111010010000",
51105 => "0111111010010000",
51106 => "0111111010010000",
51107 => "0111111010010000",
51108 => "0111111010010000",
51109 => "0111111010010000",
51110 => "0111111010010000",
51111 => "0111111010010000",
51112 => "0111111010010000",
51113 => "0111111010010000",
51114 => "0111111010010000",
51115 => "0111111010010000",
51116 => "0111111010010000",
51117 => "0111111010010000",
51118 => "0111111010010000",
51119 => "0111111010010000",
51120 => "0111111010010000",
51121 => "0111111010010000",
51122 => "0111111010010000",
51123 => "0111111010010000",
51124 => "0111111010010000",
51125 => "0111111010010000",
51126 => "0111111010010000",
51127 => "0111111010010000",
51128 => "0111111010010000",
51129 => "0111111010010000",
51130 => "0111111010010000",
51131 => "0111111010010000",
51132 => "0111111010010000",
51133 => "0111111010010000",
51134 => "0111111010010000",
51135 => "0111111010010000",
51136 => "0111111010010000",
51137 => "0111111010010000",
51138 => "0111111010010000",
51139 => "0111111010010000",
51140 => "0111111010010000",
51141 => "0111111010010000",
51142 => "0111111010010000",
51143 => "0111111010010000",
51144 => "0111111010010000",
51145 => "0111111010010000",
51146 => "0111111010010000",
51147 => "0111111010010000",
51148 => "0111111010010000",
51149 => "0111111010010000",
51150 => "0111111010010000",
51151 => "0111111010010000",
51152 => "0111111010010000",
51153 => "0111111010010000",
51154 => "0111111010010000",
51155 => "0111111010010000",
51156 => "0111111010010000",
51157 => "0111111010010000",
51158 => "0111111010010000",
51159 => "0111111010010000",
51160 => "0111111010010000",
51161 => "0111111010010000",
51162 => "0111111010010000",
51163 => "0111111010010000",
51164 => "0111111010010000",
51165 => "0111111010010000",
51166 => "0111111010010000",
51167 => "0111111010010000",
51168 => "0111111010010000",
51169 => "0111111010010000",
51170 => "0111111010010000",
51171 => "0111111010010000",
51172 => "0111111010010000",
51173 => "0111111010010000",
51174 => "0111111010010000",
51175 => "0111111010010000",
51176 => "0111111010010000",
51177 => "0111111010010000",
51178 => "0111111010010000",
51179 => "0111111010010000",
51180 => "0111111010010000",
51181 => "0111111010010000",
51182 => "0111111010010000",
51183 => "0111111010010000",
51184 => "0111111010010000",
51185 => "0111111010010000",
51186 => "0111111010010000",
51187 => "0111111010010000",
51188 => "0111111010010000",
51189 => "0111111010010000",
51190 => "0111111010010000",
51191 => "0111111010010000",
51192 => "0111111010010000",
51193 => "0111111010010000",
51194 => "0111111010010000",
51195 => "0111111010010000",
51196 => "0111111010010000",
51197 => "0111111010010000",
51198 => "0111111010010000",
51199 => "0111111010010000",
51200 => "0111111010100000",
51201 => "0111111010100000",
51202 => "0111111010100000",
51203 => "0111111010100000",
51204 => "0111111010100000",
51205 => "0111111010100000",
51206 => "0111111010100000",
51207 => "0111111010100000",
51208 => "0111111010100000",
51209 => "0111111010100000",
51210 => "0111111010100000",
51211 => "0111111010100000",
51212 => "0111111010100000",
51213 => "0111111010100000",
51214 => "0111111010100000",
51215 => "0111111010100000",
51216 => "0111111010100000",
51217 => "0111111010100000",
51218 => "0111111010100000",
51219 => "0111111010100000",
51220 => "0111111010100000",
51221 => "0111111010100000",
51222 => "0111111010100000",
51223 => "0111111010100000",
51224 => "0111111010100000",
51225 => "0111111010100000",
51226 => "0111111010100000",
51227 => "0111111010100000",
51228 => "0111111010100000",
51229 => "0111111010100000",
51230 => "0111111010100000",
51231 => "0111111010100000",
51232 => "0111111010100000",
51233 => "0111111010100000",
51234 => "0111111010100000",
51235 => "0111111010100000",
51236 => "0111111010100000",
51237 => "0111111010100000",
51238 => "0111111010100000",
51239 => "0111111010100000",
51240 => "0111111010100000",
51241 => "0111111010100000",
51242 => "0111111010100000",
51243 => "0111111010100000",
51244 => "0111111010100000",
51245 => "0111111010100000",
51246 => "0111111010100000",
51247 => "0111111010100000",
51248 => "0111111010100000",
51249 => "0111111010100000",
51250 => "0111111010100000",
51251 => "0111111010100000",
51252 => "0111111010100000",
51253 => "0111111010100000",
51254 => "0111111010100000",
51255 => "0111111010100000",
51256 => "0111111010100000",
51257 => "0111111010100000",
51258 => "0111111010100000",
51259 => "0111111010100000",
51260 => "0111111010100000",
51261 => "0111111010100000",
51262 => "0111111010100000",
51263 => "0111111010100000",
51264 => "0111111010100000",
51265 => "0111111010100000",
51266 => "0111111010100000",
51267 => "0111111010100000",
51268 => "0111111010100000",
51269 => "0111111010100000",
51270 => "0111111010100000",
51271 => "0111111010100000",
51272 => "0111111010100000",
51273 => "0111111010100000",
51274 => "0111111010100000",
51275 => "0111111010100000",
51276 => "0111111010100000",
51277 => "0111111010100000",
51278 => "0111111010100000",
51279 => "0111111010100000",
51280 => "0111111010100000",
51281 => "0111111010100000",
51282 => "0111111010100000",
51283 => "0111111010100000",
51284 => "0111111010100000",
51285 => "0111111010100000",
51286 => "0111111010100000",
51287 => "0111111010100000",
51288 => "0111111010100000",
51289 => "0111111010100000",
51290 => "0111111010100000",
51291 => "0111111010100000",
51292 => "0111111010100000",
51293 => "0111111010100000",
51294 => "0111111010100000",
51295 => "0111111010100000",
51296 => "0111111010100000",
51297 => "0111111010100000",
51298 => "0111111010100000",
51299 => "0111111010100000",
51300 => "0111111010100000",
51301 => "0111111010100000",
51302 => "0111111010100000",
51303 => "0111111010100000",
51304 => "0111111010100000",
51305 => "0111111010100000",
51306 => "0111111010100000",
51307 => "0111111010100000",
51308 => "0111111010100000",
51309 => "0111111010100000",
51310 => "0111111010100000",
51311 => "0111111010100000",
51312 => "0111111010100000",
51313 => "0111111010100000",
51314 => "0111111010100000",
51315 => "0111111010100000",
51316 => "0111111010100000",
51317 => "0111111010100000",
51318 => "0111111010100000",
51319 => "0111111010100000",
51320 => "0111111010100000",
51321 => "0111111010100000",
51322 => "0111111010100000",
51323 => "0111111010100000",
51324 => "0111111010100000",
51325 => "0111111010100000",
51326 => "0111111010100000",
51327 => "0111111010100000",
51328 => "0111111010100000",
51329 => "0111111010100000",
51330 => "0111111010100000",
51331 => "0111111010100000",
51332 => "0111111010100000",
51333 => "0111111010100000",
51334 => "0111111010100000",
51335 => "0111111010100000",
51336 => "0111111010100000",
51337 => "0111111010100000",
51338 => "0111111010100000",
51339 => "0111111010100000",
51340 => "0111111010100000",
51341 => "0111111010100000",
51342 => "0111111010100000",
51343 => "0111111010100000",
51344 => "0111111010100000",
51345 => "0111111010100000",
51346 => "0111111010100000",
51347 => "0111111010100000",
51348 => "0111111010100000",
51349 => "0111111010100000",
51350 => "0111111010100000",
51351 => "0111111010100000",
51352 => "0111111010100000",
51353 => "0111111010100000",
51354 => "0111111010100000",
51355 => "0111111010100000",
51356 => "0111111010100000",
51357 => "0111111010100000",
51358 => "0111111010100000",
51359 => "0111111010100000",
51360 => "0111111010100000",
51361 => "0111111010100000",
51362 => "0111111010100000",
51363 => "0111111010100000",
51364 => "0111111010100000",
51365 => "0111111010100000",
51366 => "0111111010100000",
51367 => "0111111010100000",
51368 => "0111111010100000",
51369 => "0111111010100000",
51370 => "0111111010100000",
51371 => "0111111010100000",
51372 => "0111111010100000",
51373 => "0111111010100000",
51374 => "0111111010100000",
51375 => "0111111010100000",
51376 => "0111111010100000",
51377 => "0111111010100000",
51378 => "0111111010100000",
51379 => "0111111010100000",
51380 => "0111111010100000",
51381 => "0111111010100000",
51382 => "0111111010100000",
51383 => "0111111010100000",
51384 => "0111111010100000",
51385 => "0111111010100000",
51386 => "0111111010100000",
51387 => "0111111010100000",
51388 => "0111111010110000",
51389 => "0111111010110000",
51390 => "0111111010110000",
51391 => "0111111010110000",
51392 => "0111111010110000",
51393 => "0111111010110000",
51394 => "0111111010110000",
51395 => "0111111010110000",
51396 => "0111111010110000",
51397 => "0111111010110000",
51398 => "0111111010110000",
51399 => "0111111010110000",
51400 => "0111111010110000",
51401 => "0111111010110000",
51402 => "0111111010110000",
51403 => "0111111010110000",
51404 => "0111111010110000",
51405 => "0111111010110000",
51406 => "0111111010110000",
51407 => "0111111010110000",
51408 => "0111111010110000",
51409 => "0111111010110000",
51410 => "0111111010110000",
51411 => "0111111010110000",
51412 => "0111111010110000",
51413 => "0111111010110000",
51414 => "0111111010110000",
51415 => "0111111010110000",
51416 => "0111111010110000",
51417 => "0111111010110000",
51418 => "0111111010110000",
51419 => "0111111010110000",
51420 => "0111111010110000",
51421 => "0111111010110000",
51422 => "0111111010110000",
51423 => "0111111010110000",
51424 => "0111111010110000",
51425 => "0111111010110000",
51426 => "0111111010110000",
51427 => "0111111010110000",
51428 => "0111111010110000",
51429 => "0111111010110000",
51430 => "0111111010110000",
51431 => "0111111010110000",
51432 => "0111111010110000",
51433 => "0111111010110000",
51434 => "0111111010110000",
51435 => "0111111010110000",
51436 => "0111111010110000",
51437 => "0111111010110000",
51438 => "0111111010110000",
51439 => "0111111010110000",
51440 => "0111111010110000",
51441 => "0111111010110000",
51442 => "0111111010110000",
51443 => "0111111010110000",
51444 => "0111111010110000",
51445 => "0111111010110000",
51446 => "0111111010110000",
51447 => "0111111010110000",
51448 => "0111111010110000",
51449 => "0111111010110000",
51450 => "0111111010110000",
51451 => "0111111010110000",
51452 => "0111111010110000",
51453 => "0111111010110000",
51454 => "0111111010110000",
51455 => "0111111010110000",
51456 => "0111111010110000",
51457 => "0111111010110000",
51458 => "0111111010110000",
51459 => "0111111010110000",
51460 => "0111111010110000",
51461 => "0111111010110000",
51462 => "0111111010110000",
51463 => "0111111010110000",
51464 => "0111111010110000",
51465 => "0111111010110000",
51466 => "0111111010110000",
51467 => "0111111010110000",
51468 => "0111111010110000",
51469 => "0111111010110000",
51470 => "0111111010110000",
51471 => "0111111010110000",
51472 => "0111111010110000",
51473 => "0111111010110000",
51474 => "0111111010110000",
51475 => "0111111010110000",
51476 => "0111111010110000",
51477 => "0111111010110000",
51478 => "0111111010110000",
51479 => "0111111010110000",
51480 => "0111111010110000",
51481 => "0111111010110000",
51482 => "0111111010110000",
51483 => "0111111010110000",
51484 => "0111111010110000",
51485 => "0111111010110000",
51486 => "0111111010110000",
51487 => "0111111010110000",
51488 => "0111111010110000",
51489 => "0111111010110000",
51490 => "0111111010110000",
51491 => "0111111010110000",
51492 => "0111111010110000",
51493 => "0111111010110000",
51494 => "0111111010110000",
51495 => "0111111010110000",
51496 => "0111111010110000",
51497 => "0111111010110000",
51498 => "0111111010110000",
51499 => "0111111010110000",
51500 => "0111111010110000",
51501 => "0111111010110000",
51502 => "0111111010110000",
51503 => "0111111010110000",
51504 => "0111111010110000",
51505 => "0111111010110000",
51506 => "0111111010110000",
51507 => "0111111010110000",
51508 => "0111111010110000",
51509 => "0111111010110000",
51510 => "0111111010110000",
51511 => "0111111010110000",
51512 => "0111111010110000",
51513 => "0111111010110000",
51514 => "0111111010110000",
51515 => "0111111010110000",
51516 => "0111111010110000",
51517 => "0111111010110000",
51518 => "0111111010110000",
51519 => "0111111010110000",
51520 => "0111111010110000",
51521 => "0111111010110000",
51522 => "0111111010110000",
51523 => "0111111010110000",
51524 => "0111111010110000",
51525 => "0111111010110000",
51526 => "0111111010110000",
51527 => "0111111010110000",
51528 => "0111111010110000",
51529 => "0111111010110000",
51530 => "0111111010110000",
51531 => "0111111010110000",
51532 => "0111111010110000",
51533 => "0111111010110000",
51534 => "0111111010110000",
51535 => "0111111010110000",
51536 => "0111111010110000",
51537 => "0111111010110000",
51538 => "0111111010110000",
51539 => "0111111010110000",
51540 => "0111111010110000",
51541 => "0111111010110000",
51542 => "0111111010110000",
51543 => "0111111010110000",
51544 => "0111111010110000",
51545 => "0111111010110000",
51546 => "0111111010110000",
51547 => "0111111010110000",
51548 => "0111111010110000",
51549 => "0111111010110000",
51550 => "0111111010110000",
51551 => "0111111010110000",
51552 => "0111111010110000",
51553 => "0111111010110000",
51554 => "0111111010110000",
51555 => "0111111010110000",
51556 => "0111111010110000",
51557 => "0111111010110000",
51558 => "0111111010110000",
51559 => "0111111010110000",
51560 => "0111111010110000",
51561 => "0111111010110000",
51562 => "0111111010110000",
51563 => "0111111010110000",
51564 => "0111111010110000",
51565 => "0111111010110000",
51566 => "0111111010110000",
51567 => "0111111010110000",
51568 => "0111111010110000",
51569 => "0111111010110000",
51570 => "0111111010110000",
51571 => "0111111010110000",
51572 => "0111111010110000",
51573 => "0111111010110000",
51574 => "0111111010110000",
51575 => "0111111010110000",
51576 => "0111111010110000",
51577 => "0111111010110000",
51578 => "0111111010110000",
51579 => "0111111010110000",
51580 => "0111111010110000",
51581 => "0111111010110000",
51582 => "0111111010110000",
51583 => "0111111010110000",
51584 => "0111111010110000",
51585 => "0111111011000000",
51586 => "0111111011000000",
51587 => "0111111011000000",
51588 => "0111111011000000",
51589 => "0111111011000000",
51590 => "0111111011000000",
51591 => "0111111011000000",
51592 => "0111111011000000",
51593 => "0111111011000000",
51594 => "0111111011000000",
51595 => "0111111011000000",
51596 => "0111111011000000",
51597 => "0111111011000000",
51598 => "0111111011000000",
51599 => "0111111011000000",
51600 => "0111111011000000",
51601 => "0111111011000000",
51602 => "0111111011000000",
51603 => "0111111011000000",
51604 => "0111111011000000",
51605 => "0111111011000000",
51606 => "0111111011000000",
51607 => "0111111011000000",
51608 => "0111111011000000",
51609 => "0111111011000000",
51610 => "0111111011000000",
51611 => "0111111011000000",
51612 => "0111111011000000",
51613 => "0111111011000000",
51614 => "0111111011000000",
51615 => "0111111011000000",
51616 => "0111111011000000",
51617 => "0111111011000000",
51618 => "0111111011000000",
51619 => "0111111011000000",
51620 => "0111111011000000",
51621 => "0111111011000000",
51622 => "0111111011000000",
51623 => "0111111011000000",
51624 => "0111111011000000",
51625 => "0111111011000000",
51626 => "0111111011000000",
51627 => "0111111011000000",
51628 => "0111111011000000",
51629 => "0111111011000000",
51630 => "0111111011000000",
51631 => "0111111011000000",
51632 => "0111111011000000",
51633 => "0111111011000000",
51634 => "0111111011000000",
51635 => "0111111011000000",
51636 => "0111111011000000",
51637 => "0111111011000000",
51638 => "0111111011000000",
51639 => "0111111011000000",
51640 => "0111111011000000",
51641 => "0111111011000000",
51642 => "0111111011000000",
51643 => "0111111011000000",
51644 => "0111111011000000",
51645 => "0111111011000000",
51646 => "0111111011000000",
51647 => "0111111011000000",
51648 => "0111111011000000",
51649 => "0111111011000000",
51650 => "0111111011000000",
51651 => "0111111011000000",
51652 => "0111111011000000",
51653 => "0111111011000000",
51654 => "0111111011000000",
51655 => "0111111011000000",
51656 => "0111111011000000",
51657 => "0111111011000000",
51658 => "0111111011000000",
51659 => "0111111011000000",
51660 => "0111111011000000",
51661 => "0111111011000000",
51662 => "0111111011000000",
51663 => "0111111011000000",
51664 => "0111111011000000",
51665 => "0111111011000000",
51666 => "0111111011000000",
51667 => "0111111011000000",
51668 => "0111111011000000",
51669 => "0111111011000000",
51670 => "0111111011000000",
51671 => "0111111011000000",
51672 => "0111111011000000",
51673 => "0111111011000000",
51674 => "0111111011000000",
51675 => "0111111011000000",
51676 => "0111111011000000",
51677 => "0111111011000000",
51678 => "0111111011000000",
51679 => "0111111011000000",
51680 => "0111111011000000",
51681 => "0111111011000000",
51682 => "0111111011000000",
51683 => "0111111011000000",
51684 => "0111111011000000",
51685 => "0111111011000000",
51686 => "0111111011000000",
51687 => "0111111011000000",
51688 => "0111111011000000",
51689 => "0111111011000000",
51690 => "0111111011000000",
51691 => "0111111011000000",
51692 => "0111111011000000",
51693 => "0111111011000000",
51694 => "0111111011000000",
51695 => "0111111011000000",
51696 => "0111111011000000",
51697 => "0111111011000000",
51698 => "0111111011000000",
51699 => "0111111011000000",
51700 => "0111111011000000",
51701 => "0111111011000000",
51702 => "0111111011000000",
51703 => "0111111011000000",
51704 => "0111111011000000",
51705 => "0111111011000000",
51706 => "0111111011000000",
51707 => "0111111011000000",
51708 => "0111111011000000",
51709 => "0111111011000000",
51710 => "0111111011000000",
51711 => "0111111011000000",
51712 => "0111111011000000",
51713 => "0111111011000000",
51714 => "0111111011000000",
51715 => "0111111011000000",
51716 => "0111111011000000",
51717 => "0111111011000000",
51718 => "0111111011000000",
51719 => "0111111011000000",
51720 => "0111111011000000",
51721 => "0111111011000000",
51722 => "0111111011000000",
51723 => "0111111011000000",
51724 => "0111111011000000",
51725 => "0111111011000000",
51726 => "0111111011000000",
51727 => "0111111011000000",
51728 => "0111111011000000",
51729 => "0111111011000000",
51730 => "0111111011000000",
51731 => "0111111011000000",
51732 => "0111111011000000",
51733 => "0111111011000000",
51734 => "0111111011000000",
51735 => "0111111011000000",
51736 => "0111111011000000",
51737 => "0111111011000000",
51738 => "0111111011000000",
51739 => "0111111011000000",
51740 => "0111111011000000",
51741 => "0111111011000000",
51742 => "0111111011000000",
51743 => "0111111011000000",
51744 => "0111111011000000",
51745 => "0111111011000000",
51746 => "0111111011000000",
51747 => "0111111011000000",
51748 => "0111111011000000",
51749 => "0111111011000000",
51750 => "0111111011000000",
51751 => "0111111011000000",
51752 => "0111111011000000",
51753 => "0111111011000000",
51754 => "0111111011000000",
51755 => "0111111011000000",
51756 => "0111111011000000",
51757 => "0111111011000000",
51758 => "0111111011000000",
51759 => "0111111011000000",
51760 => "0111111011000000",
51761 => "0111111011000000",
51762 => "0111111011000000",
51763 => "0111111011000000",
51764 => "0111111011000000",
51765 => "0111111011000000",
51766 => "0111111011000000",
51767 => "0111111011000000",
51768 => "0111111011000000",
51769 => "0111111011000000",
51770 => "0111111011000000",
51771 => "0111111011000000",
51772 => "0111111011000000",
51773 => "0111111011000000",
51774 => "0111111011000000",
51775 => "0111111011000000",
51776 => "0111111011000000",
51777 => "0111111011000000",
51778 => "0111111011000000",
51779 => "0111111011000000",
51780 => "0111111011000000",
51781 => "0111111011000000",
51782 => "0111111011000000",
51783 => "0111111011000000",
51784 => "0111111011000000",
51785 => "0111111011000000",
51786 => "0111111011000000",
51787 => "0111111011000000",
51788 => "0111111011000000",
51789 => "0111111011000000",
51790 => "0111111011000000",
51791 => "0111111011000000",
51792 => "0111111011010000",
51793 => "0111111011010000",
51794 => "0111111011010000",
51795 => "0111111011010000",
51796 => "0111111011010000",
51797 => "0111111011010000",
51798 => "0111111011010000",
51799 => "0111111011010000",
51800 => "0111111011010000",
51801 => "0111111011010000",
51802 => "0111111011010000",
51803 => "0111111011010000",
51804 => "0111111011010000",
51805 => "0111111011010000",
51806 => "0111111011010000",
51807 => "0111111011010000",
51808 => "0111111011010000",
51809 => "0111111011010000",
51810 => "0111111011010000",
51811 => "0111111011010000",
51812 => "0111111011010000",
51813 => "0111111011010000",
51814 => "0111111011010000",
51815 => "0111111011010000",
51816 => "0111111011010000",
51817 => "0111111011010000",
51818 => "0111111011010000",
51819 => "0111111011010000",
51820 => "0111111011010000",
51821 => "0111111011010000",
51822 => "0111111011010000",
51823 => "0111111011010000",
51824 => "0111111011010000",
51825 => "0111111011010000",
51826 => "0111111011010000",
51827 => "0111111011010000",
51828 => "0111111011010000",
51829 => "0111111011010000",
51830 => "0111111011010000",
51831 => "0111111011010000",
51832 => "0111111011010000",
51833 => "0111111011010000",
51834 => "0111111011010000",
51835 => "0111111011010000",
51836 => "0111111011010000",
51837 => "0111111011010000",
51838 => "0111111011010000",
51839 => "0111111011010000",
51840 => "0111111011010000",
51841 => "0111111011010000",
51842 => "0111111011010000",
51843 => "0111111011010000",
51844 => "0111111011010000",
51845 => "0111111011010000",
51846 => "0111111011010000",
51847 => "0111111011010000",
51848 => "0111111011010000",
51849 => "0111111011010000",
51850 => "0111111011010000",
51851 => "0111111011010000",
51852 => "0111111011010000",
51853 => "0111111011010000",
51854 => "0111111011010000",
51855 => "0111111011010000",
51856 => "0111111011010000",
51857 => "0111111011010000",
51858 => "0111111011010000",
51859 => "0111111011010000",
51860 => "0111111011010000",
51861 => "0111111011010000",
51862 => "0111111011010000",
51863 => "0111111011010000",
51864 => "0111111011010000",
51865 => "0111111011010000",
51866 => "0111111011010000",
51867 => "0111111011010000",
51868 => "0111111011010000",
51869 => "0111111011010000",
51870 => "0111111011010000",
51871 => "0111111011010000",
51872 => "0111111011010000",
51873 => "0111111011010000",
51874 => "0111111011010000",
51875 => "0111111011010000",
51876 => "0111111011010000",
51877 => "0111111011010000",
51878 => "0111111011010000",
51879 => "0111111011010000",
51880 => "0111111011010000",
51881 => "0111111011010000",
51882 => "0111111011010000",
51883 => "0111111011010000",
51884 => "0111111011010000",
51885 => "0111111011010000",
51886 => "0111111011010000",
51887 => "0111111011010000",
51888 => "0111111011010000",
51889 => "0111111011010000",
51890 => "0111111011010000",
51891 => "0111111011010000",
51892 => "0111111011010000",
51893 => "0111111011010000",
51894 => "0111111011010000",
51895 => "0111111011010000",
51896 => "0111111011010000",
51897 => "0111111011010000",
51898 => "0111111011010000",
51899 => "0111111011010000",
51900 => "0111111011010000",
51901 => "0111111011010000",
51902 => "0111111011010000",
51903 => "0111111011010000",
51904 => "0111111011010000",
51905 => "0111111011010000",
51906 => "0111111011010000",
51907 => "0111111011010000",
51908 => "0111111011010000",
51909 => "0111111011010000",
51910 => "0111111011010000",
51911 => "0111111011010000",
51912 => "0111111011010000",
51913 => "0111111011010000",
51914 => "0111111011010000",
51915 => "0111111011010000",
51916 => "0111111011010000",
51917 => "0111111011010000",
51918 => "0111111011010000",
51919 => "0111111011010000",
51920 => "0111111011010000",
51921 => "0111111011010000",
51922 => "0111111011010000",
51923 => "0111111011010000",
51924 => "0111111011010000",
51925 => "0111111011010000",
51926 => "0111111011010000",
51927 => "0111111011010000",
51928 => "0111111011010000",
51929 => "0111111011010000",
51930 => "0111111011010000",
51931 => "0111111011010000",
51932 => "0111111011010000",
51933 => "0111111011010000",
51934 => "0111111011010000",
51935 => "0111111011010000",
51936 => "0111111011010000",
51937 => "0111111011010000",
51938 => "0111111011010000",
51939 => "0111111011010000",
51940 => "0111111011010000",
51941 => "0111111011010000",
51942 => "0111111011010000",
51943 => "0111111011010000",
51944 => "0111111011010000",
51945 => "0111111011010000",
51946 => "0111111011010000",
51947 => "0111111011010000",
51948 => "0111111011010000",
51949 => "0111111011010000",
51950 => "0111111011010000",
51951 => "0111111011010000",
51952 => "0111111011010000",
51953 => "0111111011010000",
51954 => "0111111011010000",
51955 => "0111111011010000",
51956 => "0111111011010000",
51957 => "0111111011010000",
51958 => "0111111011010000",
51959 => "0111111011010000",
51960 => "0111111011010000",
51961 => "0111111011010000",
51962 => "0111111011010000",
51963 => "0111111011010000",
51964 => "0111111011010000",
51965 => "0111111011010000",
51966 => "0111111011010000",
51967 => "0111111011010000",
51968 => "0111111011010000",
51969 => "0111111011010000",
51970 => "0111111011010000",
51971 => "0111111011010000",
51972 => "0111111011010000",
51973 => "0111111011010000",
51974 => "0111111011010000",
51975 => "0111111011010000",
51976 => "0111111011010000",
51977 => "0111111011010000",
51978 => "0111111011010000",
51979 => "0111111011010000",
51980 => "0111111011010000",
51981 => "0111111011010000",
51982 => "0111111011010000",
51983 => "0111111011010000",
51984 => "0111111011010000",
51985 => "0111111011010000",
51986 => "0111111011010000",
51987 => "0111111011010000",
51988 => "0111111011010000",
51989 => "0111111011010000",
51990 => "0111111011010000",
51991 => "0111111011010000",
51992 => "0111111011010000",
51993 => "0111111011010000",
51994 => "0111111011010000",
51995 => "0111111011010000",
51996 => "0111111011010000",
51997 => "0111111011010000",
51998 => "0111111011010000",
51999 => "0111111011010000",
52000 => "0111111011010000",
52001 => "0111111011010000",
52002 => "0111111011010000",
52003 => "0111111011010000",
52004 => "0111111011010000",
52005 => "0111111011010000",
52006 => "0111111011010000",
52007 => "0111111011010000",
52008 => "0111111011010000",
52009 => "0111111011010000",
52010 => "0111111011100000",
52011 => "0111111011100000",
52012 => "0111111011100000",
52013 => "0111111011100000",
52014 => "0111111011100000",
52015 => "0111111011100000",
52016 => "0111111011100000",
52017 => "0111111011100000",
52018 => "0111111011100000",
52019 => "0111111011100000",
52020 => "0111111011100000",
52021 => "0111111011100000",
52022 => "0111111011100000",
52023 => "0111111011100000",
52024 => "0111111011100000",
52025 => "0111111011100000",
52026 => "0111111011100000",
52027 => "0111111011100000",
52028 => "0111111011100000",
52029 => "0111111011100000",
52030 => "0111111011100000",
52031 => "0111111011100000",
52032 => "0111111011100000",
52033 => "0111111011100000",
52034 => "0111111011100000",
52035 => "0111111011100000",
52036 => "0111111011100000",
52037 => "0111111011100000",
52038 => "0111111011100000",
52039 => "0111111011100000",
52040 => "0111111011100000",
52041 => "0111111011100000",
52042 => "0111111011100000",
52043 => "0111111011100000",
52044 => "0111111011100000",
52045 => "0111111011100000",
52046 => "0111111011100000",
52047 => "0111111011100000",
52048 => "0111111011100000",
52049 => "0111111011100000",
52050 => "0111111011100000",
52051 => "0111111011100000",
52052 => "0111111011100000",
52053 => "0111111011100000",
52054 => "0111111011100000",
52055 => "0111111011100000",
52056 => "0111111011100000",
52057 => "0111111011100000",
52058 => "0111111011100000",
52059 => "0111111011100000",
52060 => "0111111011100000",
52061 => "0111111011100000",
52062 => "0111111011100000",
52063 => "0111111011100000",
52064 => "0111111011100000",
52065 => "0111111011100000",
52066 => "0111111011100000",
52067 => "0111111011100000",
52068 => "0111111011100000",
52069 => "0111111011100000",
52070 => "0111111011100000",
52071 => "0111111011100000",
52072 => "0111111011100000",
52073 => "0111111011100000",
52074 => "0111111011100000",
52075 => "0111111011100000",
52076 => "0111111011100000",
52077 => "0111111011100000",
52078 => "0111111011100000",
52079 => "0111111011100000",
52080 => "0111111011100000",
52081 => "0111111011100000",
52082 => "0111111011100000",
52083 => "0111111011100000",
52084 => "0111111011100000",
52085 => "0111111011100000",
52086 => "0111111011100000",
52087 => "0111111011100000",
52088 => "0111111011100000",
52089 => "0111111011100000",
52090 => "0111111011100000",
52091 => "0111111011100000",
52092 => "0111111011100000",
52093 => "0111111011100000",
52094 => "0111111011100000",
52095 => "0111111011100000",
52096 => "0111111011100000",
52097 => "0111111011100000",
52098 => "0111111011100000",
52099 => "0111111011100000",
52100 => "0111111011100000",
52101 => "0111111011100000",
52102 => "0111111011100000",
52103 => "0111111011100000",
52104 => "0111111011100000",
52105 => "0111111011100000",
52106 => "0111111011100000",
52107 => "0111111011100000",
52108 => "0111111011100000",
52109 => "0111111011100000",
52110 => "0111111011100000",
52111 => "0111111011100000",
52112 => "0111111011100000",
52113 => "0111111011100000",
52114 => "0111111011100000",
52115 => "0111111011100000",
52116 => "0111111011100000",
52117 => "0111111011100000",
52118 => "0111111011100000",
52119 => "0111111011100000",
52120 => "0111111011100000",
52121 => "0111111011100000",
52122 => "0111111011100000",
52123 => "0111111011100000",
52124 => "0111111011100000",
52125 => "0111111011100000",
52126 => "0111111011100000",
52127 => "0111111011100000",
52128 => "0111111011100000",
52129 => "0111111011100000",
52130 => "0111111011100000",
52131 => "0111111011100000",
52132 => "0111111011100000",
52133 => "0111111011100000",
52134 => "0111111011100000",
52135 => "0111111011100000",
52136 => "0111111011100000",
52137 => "0111111011100000",
52138 => "0111111011100000",
52139 => "0111111011100000",
52140 => "0111111011100000",
52141 => "0111111011100000",
52142 => "0111111011100000",
52143 => "0111111011100000",
52144 => "0111111011100000",
52145 => "0111111011100000",
52146 => "0111111011100000",
52147 => "0111111011100000",
52148 => "0111111011100000",
52149 => "0111111011100000",
52150 => "0111111011100000",
52151 => "0111111011100000",
52152 => "0111111011100000",
52153 => "0111111011100000",
52154 => "0111111011100000",
52155 => "0111111011100000",
52156 => "0111111011100000",
52157 => "0111111011100000",
52158 => "0111111011100000",
52159 => "0111111011100000",
52160 => "0111111011100000",
52161 => "0111111011100000",
52162 => "0111111011100000",
52163 => "0111111011100000",
52164 => "0111111011100000",
52165 => "0111111011100000",
52166 => "0111111011100000",
52167 => "0111111011100000",
52168 => "0111111011100000",
52169 => "0111111011100000",
52170 => "0111111011100000",
52171 => "0111111011100000",
52172 => "0111111011100000",
52173 => "0111111011100000",
52174 => "0111111011100000",
52175 => "0111111011100000",
52176 => "0111111011100000",
52177 => "0111111011100000",
52178 => "0111111011100000",
52179 => "0111111011100000",
52180 => "0111111011100000",
52181 => "0111111011100000",
52182 => "0111111011100000",
52183 => "0111111011100000",
52184 => "0111111011100000",
52185 => "0111111011100000",
52186 => "0111111011100000",
52187 => "0111111011100000",
52188 => "0111111011100000",
52189 => "0111111011100000",
52190 => "0111111011100000",
52191 => "0111111011100000",
52192 => "0111111011100000",
52193 => "0111111011100000",
52194 => "0111111011100000",
52195 => "0111111011100000",
52196 => "0111111011100000",
52197 => "0111111011100000",
52198 => "0111111011100000",
52199 => "0111111011100000",
52200 => "0111111011100000",
52201 => "0111111011100000",
52202 => "0111111011100000",
52203 => "0111111011100000",
52204 => "0111111011100000",
52205 => "0111111011100000",
52206 => "0111111011100000",
52207 => "0111111011100000",
52208 => "0111111011100000",
52209 => "0111111011100000",
52210 => "0111111011100000",
52211 => "0111111011100000",
52212 => "0111111011100000",
52213 => "0111111011100000",
52214 => "0111111011100000",
52215 => "0111111011100000",
52216 => "0111111011100000",
52217 => "0111111011100000",
52218 => "0111111011100000",
52219 => "0111111011100000",
52220 => "0111111011100000",
52221 => "0111111011100000",
52222 => "0111111011100000",
52223 => "0111111011100000",
52224 => "0111111011100000",
52225 => "0111111011100000",
52226 => "0111111011100000",
52227 => "0111111011100000",
52228 => "0111111011100000",
52229 => "0111111011100000",
52230 => "0111111011100000",
52231 => "0111111011100000",
52232 => "0111111011100000",
52233 => "0111111011100000",
52234 => "0111111011100000",
52235 => "0111111011100000",
52236 => "0111111011100000",
52237 => "0111111011100000",
52238 => "0111111011100000",
52239 => "0111111011110000",
52240 => "0111111011110000",
52241 => "0111111011110000",
52242 => "0111111011110000",
52243 => "0111111011110000",
52244 => "0111111011110000",
52245 => "0111111011110000",
52246 => "0111111011110000",
52247 => "0111111011110000",
52248 => "0111111011110000",
52249 => "0111111011110000",
52250 => "0111111011110000",
52251 => "0111111011110000",
52252 => "0111111011110000",
52253 => "0111111011110000",
52254 => "0111111011110000",
52255 => "0111111011110000",
52256 => "0111111011110000",
52257 => "0111111011110000",
52258 => "0111111011110000",
52259 => "0111111011110000",
52260 => "0111111011110000",
52261 => "0111111011110000",
52262 => "0111111011110000",
52263 => "0111111011110000",
52264 => "0111111011110000",
52265 => "0111111011110000",
52266 => "0111111011110000",
52267 => "0111111011110000",
52268 => "0111111011110000",
52269 => "0111111011110000",
52270 => "0111111011110000",
52271 => "0111111011110000",
52272 => "0111111011110000",
52273 => "0111111011110000",
52274 => "0111111011110000",
52275 => "0111111011110000",
52276 => "0111111011110000",
52277 => "0111111011110000",
52278 => "0111111011110000",
52279 => "0111111011110000",
52280 => "0111111011110000",
52281 => "0111111011110000",
52282 => "0111111011110000",
52283 => "0111111011110000",
52284 => "0111111011110000",
52285 => "0111111011110000",
52286 => "0111111011110000",
52287 => "0111111011110000",
52288 => "0111111011110000",
52289 => "0111111011110000",
52290 => "0111111011110000",
52291 => "0111111011110000",
52292 => "0111111011110000",
52293 => "0111111011110000",
52294 => "0111111011110000",
52295 => "0111111011110000",
52296 => "0111111011110000",
52297 => "0111111011110000",
52298 => "0111111011110000",
52299 => "0111111011110000",
52300 => "0111111011110000",
52301 => "0111111011110000",
52302 => "0111111011110000",
52303 => "0111111011110000",
52304 => "0111111011110000",
52305 => "0111111011110000",
52306 => "0111111011110000",
52307 => "0111111011110000",
52308 => "0111111011110000",
52309 => "0111111011110000",
52310 => "0111111011110000",
52311 => "0111111011110000",
52312 => "0111111011110000",
52313 => "0111111011110000",
52314 => "0111111011110000",
52315 => "0111111011110000",
52316 => "0111111011110000",
52317 => "0111111011110000",
52318 => "0111111011110000",
52319 => "0111111011110000",
52320 => "0111111011110000",
52321 => "0111111011110000",
52322 => "0111111011110000",
52323 => "0111111011110000",
52324 => "0111111011110000",
52325 => "0111111011110000",
52326 => "0111111011110000",
52327 => "0111111011110000",
52328 => "0111111011110000",
52329 => "0111111011110000",
52330 => "0111111011110000",
52331 => "0111111011110000",
52332 => "0111111011110000",
52333 => "0111111011110000",
52334 => "0111111011110000",
52335 => "0111111011110000",
52336 => "0111111011110000",
52337 => "0111111011110000",
52338 => "0111111011110000",
52339 => "0111111011110000",
52340 => "0111111011110000",
52341 => "0111111011110000",
52342 => "0111111011110000",
52343 => "0111111011110000",
52344 => "0111111011110000",
52345 => "0111111011110000",
52346 => "0111111011110000",
52347 => "0111111011110000",
52348 => "0111111011110000",
52349 => "0111111011110000",
52350 => "0111111011110000",
52351 => "0111111011110000",
52352 => "0111111011110000",
52353 => "0111111011110000",
52354 => "0111111011110000",
52355 => "0111111011110000",
52356 => "0111111011110000",
52357 => "0111111011110000",
52358 => "0111111011110000",
52359 => "0111111011110000",
52360 => "0111111011110000",
52361 => "0111111011110000",
52362 => "0111111011110000",
52363 => "0111111011110000",
52364 => "0111111011110000",
52365 => "0111111011110000",
52366 => "0111111011110000",
52367 => "0111111011110000",
52368 => "0111111011110000",
52369 => "0111111011110000",
52370 => "0111111011110000",
52371 => "0111111011110000",
52372 => "0111111011110000",
52373 => "0111111011110000",
52374 => "0111111011110000",
52375 => "0111111011110000",
52376 => "0111111011110000",
52377 => "0111111011110000",
52378 => "0111111011110000",
52379 => "0111111011110000",
52380 => "0111111011110000",
52381 => "0111111011110000",
52382 => "0111111011110000",
52383 => "0111111011110000",
52384 => "0111111011110000",
52385 => "0111111011110000",
52386 => "0111111011110000",
52387 => "0111111011110000",
52388 => "0111111011110000",
52389 => "0111111011110000",
52390 => "0111111011110000",
52391 => "0111111011110000",
52392 => "0111111011110000",
52393 => "0111111011110000",
52394 => "0111111011110000",
52395 => "0111111011110000",
52396 => "0111111011110000",
52397 => "0111111011110000",
52398 => "0111111011110000",
52399 => "0111111011110000",
52400 => "0111111011110000",
52401 => "0111111011110000",
52402 => "0111111011110000",
52403 => "0111111011110000",
52404 => "0111111011110000",
52405 => "0111111011110000",
52406 => "0111111011110000",
52407 => "0111111011110000",
52408 => "0111111011110000",
52409 => "0111111011110000",
52410 => "0111111011110000",
52411 => "0111111011110000",
52412 => "0111111011110000",
52413 => "0111111011110000",
52414 => "0111111011110000",
52415 => "0111111011110000",
52416 => "0111111011110000",
52417 => "0111111011110000",
52418 => "0111111011110000",
52419 => "0111111011110000",
52420 => "0111111011110000",
52421 => "0111111011110000",
52422 => "0111111011110000",
52423 => "0111111011110000",
52424 => "0111111011110000",
52425 => "0111111011110000",
52426 => "0111111011110000",
52427 => "0111111011110000",
52428 => "0111111011110000",
52429 => "0111111011110000",
52430 => "0111111011110000",
52431 => "0111111011110000",
52432 => "0111111011110000",
52433 => "0111111011110000",
52434 => "0111111011110000",
52435 => "0111111011110000",
52436 => "0111111011110000",
52437 => "0111111011110000",
52438 => "0111111011110000",
52439 => "0111111011110000",
52440 => "0111111011110000",
52441 => "0111111011110000",
52442 => "0111111011110000",
52443 => "0111111011110000",
52444 => "0111111011110000",
52445 => "0111111011110000",
52446 => "0111111011110000",
52447 => "0111111011110000",
52448 => "0111111011110000",
52449 => "0111111011110000",
52450 => "0111111011110000",
52451 => "0111111011110000",
52452 => "0111111011110000",
52453 => "0111111011110000",
52454 => "0111111011110000",
52455 => "0111111011110000",
52456 => "0111111011110000",
52457 => "0111111011110000",
52458 => "0111111011110000",
52459 => "0111111011110000",
52460 => "0111111011110000",
52461 => "0111111011110000",
52462 => "0111111011110000",
52463 => "0111111011110000",
52464 => "0111111011110000",
52465 => "0111111011110000",
52466 => "0111111011110000",
52467 => "0111111011110000",
52468 => "0111111011110000",
52469 => "0111111011110000",
52470 => "0111111011110000",
52471 => "0111111011110000",
52472 => "0111111011110000",
52473 => "0111111011110000",
52474 => "0111111011110000",
52475 => "0111111011110000",
52476 => "0111111011110000",
52477 => "0111111011110000",
52478 => "0111111011110000",
52479 => "0111111011110000",
52480 => "0111111011110000",
52481 => "0111111011110000",
52482 => "0111111100000000",
52483 => "0111111100000000",
52484 => "0111111100000000",
52485 => "0111111100000000",
52486 => "0111111100000000",
52487 => "0111111100000000",
52488 => "0111111100000000",
52489 => "0111111100000000",
52490 => "0111111100000000",
52491 => "0111111100000000",
52492 => "0111111100000000",
52493 => "0111111100000000",
52494 => "0111111100000000",
52495 => "0111111100000000",
52496 => "0111111100000000",
52497 => "0111111100000000",
52498 => "0111111100000000",
52499 => "0111111100000000",
52500 => "0111111100000000",
52501 => "0111111100000000",
52502 => "0111111100000000",
52503 => "0111111100000000",
52504 => "0111111100000000",
52505 => "0111111100000000",
52506 => "0111111100000000",
52507 => "0111111100000000",
52508 => "0111111100000000",
52509 => "0111111100000000",
52510 => "0111111100000000",
52511 => "0111111100000000",
52512 => "0111111100000000",
52513 => "0111111100000000",
52514 => "0111111100000000",
52515 => "0111111100000000",
52516 => "0111111100000000",
52517 => "0111111100000000",
52518 => "0111111100000000",
52519 => "0111111100000000",
52520 => "0111111100000000",
52521 => "0111111100000000",
52522 => "0111111100000000",
52523 => "0111111100000000",
52524 => "0111111100000000",
52525 => "0111111100000000",
52526 => "0111111100000000",
52527 => "0111111100000000",
52528 => "0111111100000000",
52529 => "0111111100000000",
52530 => "0111111100000000",
52531 => "0111111100000000",
52532 => "0111111100000000",
52533 => "0111111100000000",
52534 => "0111111100000000",
52535 => "0111111100000000",
52536 => "0111111100000000",
52537 => "0111111100000000",
52538 => "0111111100000000",
52539 => "0111111100000000",
52540 => "0111111100000000",
52541 => "0111111100000000",
52542 => "0111111100000000",
52543 => "0111111100000000",
52544 => "0111111100000000",
52545 => "0111111100000000",
52546 => "0111111100000000",
52547 => "0111111100000000",
52548 => "0111111100000000",
52549 => "0111111100000000",
52550 => "0111111100000000",
52551 => "0111111100000000",
52552 => "0111111100000000",
52553 => "0111111100000000",
52554 => "0111111100000000",
52555 => "0111111100000000",
52556 => "0111111100000000",
52557 => "0111111100000000",
52558 => "0111111100000000",
52559 => "0111111100000000",
52560 => "0111111100000000",
52561 => "0111111100000000",
52562 => "0111111100000000",
52563 => "0111111100000000",
52564 => "0111111100000000",
52565 => "0111111100000000",
52566 => "0111111100000000",
52567 => "0111111100000000",
52568 => "0111111100000000",
52569 => "0111111100000000",
52570 => "0111111100000000",
52571 => "0111111100000000",
52572 => "0111111100000000",
52573 => "0111111100000000",
52574 => "0111111100000000",
52575 => "0111111100000000",
52576 => "0111111100000000",
52577 => "0111111100000000",
52578 => "0111111100000000",
52579 => "0111111100000000",
52580 => "0111111100000000",
52581 => "0111111100000000",
52582 => "0111111100000000",
52583 => "0111111100000000",
52584 => "0111111100000000",
52585 => "0111111100000000",
52586 => "0111111100000000",
52587 => "0111111100000000",
52588 => "0111111100000000",
52589 => "0111111100000000",
52590 => "0111111100000000",
52591 => "0111111100000000",
52592 => "0111111100000000",
52593 => "0111111100000000",
52594 => "0111111100000000",
52595 => "0111111100000000",
52596 => "0111111100000000",
52597 => "0111111100000000",
52598 => "0111111100000000",
52599 => "0111111100000000",
52600 => "0111111100000000",
52601 => "0111111100000000",
52602 => "0111111100000000",
52603 => "0111111100000000",
52604 => "0111111100000000",
52605 => "0111111100000000",
52606 => "0111111100000000",
52607 => "0111111100000000",
52608 => "0111111100000000",
52609 => "0111111100000000",
52610 => "0111111100000000",
52611 => "0111111100000000",
52612 => "0111111100000000",
52613 => "0111111100000000",
52614 => "0111111100000000",
52615 => "0111111100000000",
52616 => "0111111100000000",
52617 => "0111111100000000",
52618 => "0111111100000000",
52619 => "0111111100000000",
52620 => "0111111100000000",
52621 => "0111111100000000",
52622 => "0111111100000000",
52623 => "0111111100000000",
52624 => "0111111100000000",
52625 => "0111111100000000",
52626 => "0111111100000000",
52627 => "0111111100000000",
52628 => "0111111100000000",
52629 => "0111111100000000",
52630 => "0111111100000000",
52631 => "0111111100000000",
52632 => "0111111100000000",
52633 => "0111111100000000",
52634 => "0111111100000000",
52635 => "0111111100000000",
52636 => "0111111100000000",
52637 => "0111111100000000",
52638 => "0111111100000000",
52639 => "0111111100000000",
52640 => "0111111100000000",
52641 => "0111111100000000",
52642 => "0111111100000000",
52643 => "0111111100000000",
52644 => "0111111100000000",
52645 => "0111111100000000",
52646 => "0111111100000000",
52647 => "0111111100000000",
52648 => "0111111100000000",
52649 => "0111111100000000",
52650 => "0111111100000000",
52651 => "0111111100000000",
52652 => "0111111100000000",
52653 => "0111111100000000",
52654 => "0111111100000000",
52655 => "0111111100000000",
52656 => "0111111100000000",
52657 => "0111111100000000",
52658 => "0111111100000000",
52659 => "0111111100000000",
52660 => "0111111100000000",
52661 => "0111111100000000",
52662 => "0111111100000000",
52663 => "0111111100000000",
52664 => "0111111100000000",
52665 => "0111111100000000",
52666 => "0111111100000000",
52667 => "0111111100000000",
52668 => "0111111100000000",
52669 => "0111111100000000",
52670 => "0111111100000000",
52671 => "0111111100000000",
52672 => "0111111100000000",
52673 => "0111111100000000",
52674 => "0111111100000000",
52675 => "0111111100000000",
52676 => "0111111100000000",
52677 => "0111111100000000",
52678 => "0111111100000000",
52679 => "0111111100000000",
52680 => "0111111100000000",
52681 => "0111111100000000",
52682 => "0111111100000000",
52683 => "0111111100000000",
52684 => "0111111100000000",
52685 => "0111111100000000",
52686 => "0111111100000000",
52687 => "0111111100000000",
52688 => "0111111100000000",
52689 => "0111111100000000",
52690 => "0111111100000000",
52691 => "0111111100000000",
52692 => "0111111100000000",
52693 => "0111111100000000",
52694 => "0111111100000000",
52695 => "0111111100000000",
52696 => "0111111100000000",
52697 => "0111111100000000",
52698 => "0111111100000000",
52699 => "0111111100000000",
52700 => "0111111100000000",
52701 => "0111111100000000",
52702 => "0111111100000000",
52703 => "0111111100000000",
52704 => "0111111100000000",
52705 => "0111111100000000",
52706 => "0111111100000000",
52707 => "0111111100000000",
52708 => "0111111100000000",
52709 => "0111111100000000",
52710 => "0111111100000000",
52711 => "0111111100000000",
52712 => "0111111100000000",
52713 => "0111111100000000",
52714 => "0111111100000000",
52715 => "0111111100000000",
52716 => "0111111100000000",
52717 => "0111111100000000",
52718 => "0111111100000000",
52719 => "0111111100000000",
52720 => "0111111100000000",
52721 => "0111111100000000",
52722 => "0111111100000000",
52723 => "0111111100000000",
52724 => "0111111100000000",
52725 => "0111111100000000",
52726 => "0111111100000000",
52727 => "0111111100000000",
52728 => "0111111100000000",
52729 => "0111111100000000",
52730 => "0111111100000000",
52731 => "0111111100000000",
52732 => "0111111100000000",
52733 => "0111111100000000",
52734 => "0111111100000000",
52735 => "0111111100000000",
52736 => "0111111100000000",
52737 => "0111111100000000",
52738 => "0111111100000000",
52739 => "0111111100000000",
52740 => "0111111100000000",
52741 => "0111111100010000",
52742 => "0111111100010000",
52743 => "0111111100010000",
52744 => "0111111100010000",
52745 => "0111111100010000",
52746 => "0111111100010000",
52747 => "0111111100010000",
52748 => "0111111100010000",
52749 => "0111111100010000",
52750 => "0111111100010000",
52751 => "0111111100010000",
52752 => "0111111100010000",
52753 => "0111111100010000",
52754 => "0111111100010000",
52755 => "0111111100010000",
52756 => "0111111100010000",
52757 => "0111111100010000",
52758 => "0111111100010000",
52759 => "0111111100010000",
52760 => "0111111100010000",
52761 => "0111111100010000",
52762 => "0111111100010000",
52763 => "0111111100010000",
52764 => "0111111100010000",
52765 => "0111111100010000",
52766 => "0111111100010000",
52767 => "0111111100010000",
52768 => "0111111100010000",
52769 => "0111111100010000",
52770 => "0111111100010000",
52771 => "0111111100010000",
52772 => "0111111100010000",
52773 => "0111111100010000",
52774 => "0111111100010000",
52775 => "0111111100010000",
52776 => "0111111100010000",
52777 => "0111111100010000",
52778 => "0111111100010000",
52779 => "0111111100010000",
52780 => "0111111100010000",
52781 => "0111111100010000",
52782 => "0111111100010000",
52783 => "0111111100010000",
52784 => "0111111100010000",
52785 => "0111111100010000",
52786 => "0111111100010000",
52787 => "0111111100010000",
52788 => "0111111100010000",
52789 => "0111111100010000",
52790 => "0111111100010000",
52791 => "0111111100010000",
52792 => "0111111100010000",
52793 => "0111111100010000",
52794 => "0111111100010000",
52795 => "0111111100010000",
52796 => "0111111100010000",
52797 => "0111111100010000",
52798 => "0111111100010000",
52799 => "0111111100010000",
52800 => "0111111100010000",
52801 => "0111111100010000",
52802 => "0111111100010000",
52803 => "0111111100010000",
52804 => "0111111100010000",
52805 => "0111111100010000",
52806 => "0111111100010000",
52807 => "0111111100010000",
52808 => "0111111100010000",
52809 => "0111111100010000",
52810 => "0111111100010000",
52811 => "0111111100010000",
52812 => "0111111100010000",
52813 => "0111111100010000",
52814 => "0111111100010000",
52815 => "0111111100010000",
52816 => "0111111100010000",
52817 => "0111111100010000",
52818 => "0111111100010000",
52819 => "0111111100010000",
52820 => "0111111100010000",
52821 => "0111111100010000",
52822 => "0111111100010000",
52823 => "0111111100010000",
52824 => "0111111100010000",
52825 => "0111111100010000",
52826 => "0111111100010000",
52827 => "0111111100010000",
52828 => "0111111100010000",
52829 => "0111111100010000",
52830 => "0111111100010000",
52831 => "0111111100010000",
52832 => "0111111100010000",
52833 => "0111111100010000",
52834 => "0111111100010000",
52835 => "0111111100010000",
52836 => "0111111100010000",
52837 => "0111111100010000",
52838 => "0111111100010000",
52839 => "0111111100010000",
52840 => "0111111100010000",
52841 => "0111111100010000",
52842 => "0111111100010000",
52843 => "0111111100010000",
52844 => "0111111100010000",
52845 => "0111111100010000",
52846 => "0111111100010000",
52847 => "0111111100010000",
52848 => "0111111100010000",
52849 => "0111111100010000",
52850 => "0111111100010000",
52851 => "0111111100010000",
52852 => "0111111100010000",
52853 => "0111111100010000",
52854 => "0111111100010000",
52855 => "0111111100010000",
52856 => "0111111100010000",
52857 => "0111111100010000",
52858 => "0111111100010000",
52859 => "0111111100010000",
52860 => "0111111100010000",
52861 => "0111111100010000",
52862 => "0111111100010000",
52863 => "0111111100010000",
52864 => "0111111100010000",
52865 => "0111111100010000",
52866 => "0111111100010000",
52867 => "0111111100010000",
52868 => "0111111100010000",
52869 => "0111111100010000",
52870 => "0111111100010000",
52871 => "0111111100010000",
52872 => "0111111100010000",
52873 => "0111111100010000",
52874 => "0111111100010000",
52875 => "0111111100010000",
52876 => "0111111100010000",
52877 => "0111111100010000",
52878 => "0111111100010000",
52879 => "0111111100010000",
52880 => "0111111100010000",
52881 => "0111111100010000",
52882 => "0111111100010000",
52883 => "0111111100010000",
52884 => "0111111100010000",
52885 => "0111111100010000",
52886 => "0111111100010000",
52887 => "0111111100010000",
52888 => "0111111100010000",
52889 => "0111111100010000",
52890 => "0111111100010000",
52891 => "0111111100010000",
52892 => "0111111100010000",
52893 => "0111111100010000",
52894 => "0111111100010000",
52895 => "0111111100010000",
52896 => "0111111100010000",
52897 => "0111111100010000",
52898 => "0111111100010000",
52899 => "0111111100010000",
52900 => "0111111100010000",
52901 => "0111111100010000",
52902 => "0111111100010000",
52903 => "0111111100010000",
52904 => "0111111100010000",
52905 => "0111111100010000",
52906 => "0111111100010000",
52907 => "0111111100010000",
52908 => "0111111100010000",
52909 => "0111111100010000",
52910 => "0111111100010000",
52911 => "0111111100010000",
52912 => "0111111100010000",
52913 => "0111111100010000",
52914 => "0111111100010000",
52915 => "0111111100010000",
52916 => "0111111100010000",
52917 => "0111111100010000",
52918 => "0111111100010000",
52919 => "0111111100010000",
52920 => "0111111100010000",
52921 => "0111111100010000",
52922 => "0111111100010000",
52923 => "0111111100010000",
52924 => "0111111100010000",
52925 => "0111111100010000",
52926 => "0111111100010000",
52927 => "0111111100010000",
52928 => "0111111100010000",
52929 => "0111111100010000",
52930 => "0111111100010000",
52931 => "0111111100010000",
52932 => "0111111100010000",
52933 => "0111111100010000",
52934 => "0111111100010000",
52935 => "0111111100010000",
52936 => "0111111100010000",
52937 => "0111111100010000",
52938 => "0111111100010000",
52939 => "0111111100010000",
52940 => "0111111100010000",
52941 => "0111111100010000",
52942 => "0111111100010000",
52943 => "0111111100010000",
52944 => "0111111100010000",
52945 => "0111111100010000",
52946 => "0111111100010000",
52947 => "0111111100010000",
52948 => "0111111100010000",
52949 => "0111111100010000",
52950 => "0111111100010000",
52951 => "0111111100010000",
52952 => "0111111100010000",
52953 => "0111111100010000",
52954 => "0111111100010000",
52955 => "0111111100010000",
52956 => "0111111100010000",
52957 => "0111111100010000",
52958 => "0111111100010000",
52959 => "0111111100010000",
52960 => "0111111100010000",
52961 => "0111111100010000",
52962 => "0111111100010000",
52963 => "0111111100010000",
52964 => "0111111100010000",
52965 => "0111111100010000",
52966 => "0111111100010000",
52967 => "0111111100010000",
52968 => "0111111100010000",
52969 => "0111111100010000",
52970 => "0111111100010000",
52971 => "0111111100010000",
52972 => "0111111100010000",
52973 => "0111111100010000",
52974 => "0111111100010000",
52975 => "0111111100010000",
52976 => "0111111100010000",
52977 => "0111111100010000",
52978 => "0111111100010000",
52979 => "0111111100010000",
52980 => "0111111100010000",
52981 => "0111111100010000",
52982 => "0111111100010000",
52983 => "0111111100010000",
52984 => "0111111100010000",
52985 => "0111111100010000",
52986 => "0111111100010000",
52987 => "0111111100010000",
52988 => "0111111100010000",
52989 => "0111111100010000",
52990 => "0111111100010000",
52991 => "0111111100010000",
52992 => "0111111100010000",
52993 => "0111111100010000",
52994 => "0111111100010000",
52995 => "0111111100010000",
52996 => "0111111100010000",
52997 => "0111111100010000",
52998 => "0111111100010000",
52999 => "0111111100010000",
53000 => "0111111100010000",
53001 => "0111111100010000",
53002 => "0111111100010000",
53003 => "0111111100010000",
53004 => "0111111100010000",
53005 => "0111111100010000",
53006 => "0111111100010000",
53007 => "0111111100010000",
53008 => "0111111100010000",
53009 => "0111111100010000",
53010 => "0111111100010000",
53011 => "0111111100010000",
53012 => "0111111100010000",
53013 => "0111111100010000",
53014 => "0111111100010000",
53015 => "0111111100010000",
53016 => "0111111100100000",
53017 => "0111111100100000",
53018 => "0111111100100000",
53019 => "0111111100100000",
53020 => "0111111100100000",
53021 => "0111111100100000",
53022 => "0111111100100000",
53023 => "0111111100100000",
53024 => "0111111100100000",
53025 => "0111111100100000",
53026 => "0111111100100000",
53027 => "0111111100100000",
53028 => "0111111100100000",
53029 => "0111111100100000",
53030 => "0111111100100000",
53031 => "0111111100100000",
53032 => "0111111100100000",
53033 => "0111111100100000",
53034 => "0111111100100000",
53035 => "0111111100100000",
53036 => "0111111100100000",
53037 => "0111111100100000",
53038 => "0111111100100000",
53039 => "0111111100100000",
53040 => "0111111100100000",
53041 => "0111111100100000",
53042 => "0111111100100000",
53043 => "0111111100100000",
53044 => "0111111100100000",
53045 => "0111111100100000",
53046 => "0111111100100000",
53047 => "0111111100100000",
53048 => "0111111100100000",
53049 => "0111111100100000",
53050 => "0111111100100000",
53051 => "0111111100100000",
53052 => "0111111100100000",
53053 => "0111111100100000",
53054 => "0111111100100000",
53055 => "0111111100100000",
53056 => "0111111100100000",
53057 => "0111111100100000",
53058 => "0111111100100000",
53059 => "0111111100100000",
53060 => "0111111100100000",
53061 => "0111111100100000",
53062 => "0111111100100000",
53063 => "0111111100100000",
53064 => "0111111100100000",
53065 => "0111111100100000",
53066 => "0111111100100000",
53067 => "0111111100100000",
53068 => "0111111100100000",
53069 => "0111111100100000",
53070 => "0111111100100000",
53071 => "0111111100100000",
53072 => "0111111100100000",
53073 => "0111111100100000",
53074 => "0111111100100000",
53075 => "0111111100100000",
53076 => "0111111100100000",
53077 => "0111111100100000",
53078 => "0111111100100000",
53079 => "0111111100100000",
53080 => "0111111100100000",
53081 => "0111111100100000",
53082 => "0111111100100000",
53083 => "0111111100100000",
53084 => "0111111100100000",
53085 => "0111111100100000",
53086 => "0111111100100000",
53087 => "0111111100100000",
53088 => "0111111100100000",
53089 => "0111111100100000",
53090 => "0111111100100000",
53091 => "0111111100100000",
53092 => "0111111100100000",
53093 => "0111111100100000",
53094 => "0111111100100000",
53095 => "0111111100100000",
53096 => "0111111100100000",
53097 => "0111111100100000",
53098 => "0111111100100000",
53099 => "0111111100100000",
53100 => "0111111100100000",
53101 => "0111111100100000",
53102 => "0111111100100000",
53103 => "0111111100100000",
53104 => "0111111100100000",
53105 => "0111111100100000",
53106 => "0111111100100000",
53107 => "0111111100100000",
53108 => "0111111100100000",
53109 => "0111111100100000",
53110 => "0111111100100000",
53111 => "0111111100100000",
53112 => "0111111100100000",
53113 => "0111111100100000",
53114 => "0111111100100000",
53115 => "0111111100100000",
53116 => "0111111100100000",
53117 => "0111111100100000",
53118 => "0111111100100000",
53119 => "0111111100100000",
53120 => "0111111100100000",
53121 => "0111111100100000",
53122 => "0111111100100000",
53123 => "0111111100100000",
53124 => "0111111100100000",
53125 => "0111111100100000",
53126 => "0111111100100000",
53127 => "0111111100100000",
53128 => "0111111100100000",
53129 => "0111111100100000",
53130 => "0111111100100000",
53131 => "0111111100100000",
53132 => "0111111100100000",
53133 => "0111111100100000",
53134 => "0111111100100000",
53135 => "0111111100100000",
53136 => "0111111100100000",
53137 => "0111111100100000",
53138 => "0111111100100000",
53139 => "0111111100100000",
53140 => "0111111100100000",
53141 => "0111111100100000",
53142 => "0111111100100000",
53143 => "0111111100100000",
53144 => "0111111100100000",
53145 => "0111111100100000",
53146 => "0111111100100000",
53147 => "0111111100100000",
53148 => "0111111100100000",
53149 => "0111111100100000",
53150 => "0111111100100000",
53151 => "0111111100100000",
53152 => "0111111100100000",
53153 => "0111111100100000",
53154 => "0111111100100000",
53155 => "0111111100100000",
53156 => "0111111100100000",
53157 => "0111111100100000",
53158 => "0111111100100000",
53159 => "0111111100100000",
53160 => "0111111100100000",
53161 => "0111111100100000",
53162 => "0111111100100000",
53163 => "0111111100100000",
53164 => "0111111100100000",
53165 => "0111111100100000",
53166 => "0111111100100000",
53167 => "0111111100100000",
53168 => "0111111100100000",
53169 => "0111111100100000",
53170 => "0111111100100000",
53171 => "0111111100100000",
53172 => "0111111100100000",
53173 => "0111111100100000",
53174 => "0111111100100000",
53175 => "0111111100100000",
53176 => "0111111100100000",
53177 => "0111111100100000",
53178 => "0111111100100000",
53179 => "0111111100100000",
53180 => "0111111100100000",
53181 => "0111111100100000",
53182 => "0111111100100000",
53183 => "0111111100100000",
53184 => "0111111100100000",
53185 => "0111111100100000",
53186 => "0111111100100000",
53187 => "0111111100100000",
53188 => "0111111100100000",
53189 => "0111111100100000",
53190 => "0111111100100000",
53191 => "0111111100100000",
53192 => "0111111100100000",
53193 => "0111111100100000",
53194 => "0111111100100000",
53195 => "0111111100100000",
53196 => "0111111100100000",
53197 => "0111111100100000",
53198 => "0111111100100000",
53199 => "0111111100100000",
53200 => "0111111100100000",
53201 => "0111111100100000",
53202 => "0111111100100000",
53203 => "0111111100100000",
53204 => "0111111100100000",
53205 => "0111111100100000",
53206 => "0111111100100000",
53207 => "0111111100100000",
53208 => "0111111100100000",
53209 => "0111111100100000",
53210 => "0111111100100000",
53211 => "0111111100100000",
53212 => "0111111100100000",
53213 => "0111111100100000",
53214 => "0111111100100000",
53215 => "0111111100100000",
53216 => "0111111100100000",
53217 => "0111111100100000",
53218 => "0111111100100000",
53219 => "0111111100100000",
53220 => "0111111100100000",
53221 => "0111111100100000",
53222 => "0111111100100000",
53223 => "0111111100100000",
53224 => "0111111100100000",
53225 => "0111111100100000",
53226 => "0111111100100000",
53227 => "0111111100100000",
53228 => "0111111100100000",
53229 => "0111111100100000",
53230 => "0111111100100000",
53231 => "0111111100100000",
53232 => "0111111100100000",
53233 => "0111111100100000",
53234 => "0111111100100000",
53235 => "0111111100100000",
53236 => "0111111100100000",
53237 => "0111111100100000",
53238 => "0111111100100000",
53239 => "0111111100100000",
53240 => "0111111100100000",
53241 => "0111111100100000",
53242 => "0111111100100000",
53243 => "0111111100100000",
53244 => "0111111100100000",
53245 => "0111111100100000",
53246 => "0111111100100000",
53247 => "0111111100100000",
53248 => "0111111100100000",
53249 => "0111111100100000",
53250 => "0111111100100000",
53251 => "0111111100100000",
53252 => "0111111100100000",
53253 => "0111111100100000",
53254 => "0111111100100000",
53255 => "0111111100100000",
53256 => "0111111100100000",
53257 => "0111111100100000",
53258 => "0111111100100000",
53259 => "0111111100100000",
53260 => "0111111100100000",
53261 => "0111111100100000",
53262 => "0111111100100000",
53263 => "0111111100100000",
53264 => "0111111100100000",
53265 => "0111111100100000",
53266 => "0111111100100000",
53267 => "0111111100100000",
53268 => "0111111100100000",
53269 => "0111111100100000",
53270 => "0111111100100000",
53271 => "0111111100100000",
53272 => "0111111100100000",
53273 => "0111111100100000",
53274 => "0111111100100000",
53275 => "0111111100100000",
53276 => "0111111100100000",
53277 => "0111111100100000",
53278 => "0111111100100000",
53279 => "0111111100100000",
53280 => "0111111100100000",
53281 => "0111111100100000",
53282 => "0111111100100000",
53283 => "0111111100100000",
53284 => "0111111100100000",
53285 => "0111111100100000",
53286 => "0111111100100000",
53287 => "0111111100100000",
53288 => "0111111100100000",
53289 => "0111111100100000",
53290 => "0111111100100000",
53291 => "0111111100100000",
53292 => "0111111100100000",
53293 => "0111111100100000",
53294 => "0111111100100000",
53295 => "0111111100100000",
53296 => "0111111100100000",
53297 => "0111111100100000",
53298 => "0111111100100000",
53299 => "0111111100100000",
53300 => "0111111100100000",
53301 => "0111111100100000",
53302 => "0111111100100000",
53303 => "0111111100100000",
53304 => "0111111100100000",
53305 => "0111111100100000",
53306 => "0111111100100000",
53307 => "0111111100100000",
53308 => "0111111100100000",
53309 => "0111111100100000",
53310 => "0111111100110000",
53311 => "0111111100110000",
53312 => "0111111100110000",
53313 => "0111111100110000",
53314 => "0111111100110000",
53315 => "0111111100110000",
53316 => "0111111100110000",
53317 => "0111111100110000",
53318 => "0111111100110000",
53319 => "0111111100110000",
53320 => "0111111100110000",
53321 => "0111111100110000",
53322 => "0111111100110000",
53323 => "0111111100110000",
53324 => "0111111100110000",
53325 => "0111111100110000",
53326 => "0111111100110000",
53327 => "0111111100110000",
53328 => "0111111100110000",
53329 => "0111111100110000",
53330 => "0111111100110000",
53331 => "0111111100110000",
53332 => "0111111100110000",
53333 => "0111111100110000",
53334 => "0111111100110000",
53335 => "0111111100110000",
53336 => "0111111100110000",
53337 => "0111111100110000",
53338 => "0111111100110000",
53339 => "0111111100110000",
53340 => "0111111100110000",
53341 => "0111111100110000",
53342 => "0111111100110000",
53343 => "0111111100110000",
53344 => "0111111100110000",
53345 => "0111111100110000",
53346 => "0111111100110000",
53347 => "0111111100110000",
53348 => "0111111100110000",
53349 => "0111111100110000",
53350 => "0111111100110000",
53351 => "0111111100110000",
53352 => "0111111100110000",
53353 => "0111111100110000",
53354 => "0111111100110000",
53355 => "0111111100110000",
53356 => "0111111100110000",
53357 => "0111111100110000",
53358 => "0111111100110000",
53359 => "0111111100110000",
53360 => "0111111100110000",
53361 => "0111111100110000",
53362 => "0111111100110000",
53363 => "0111111100110000",
53364 => "0111111100110000",
53365 => "0111111100110000",
53366 => "0111111100110000",
53367 => "0111111100110000",
53368 => "0111111100110000",
53369 => "0111111100110000",
53370 => "0111111100110000",
53371 => "0111111100110000",
53372 => "0111111100110000",
53373 => "0111111100110000",
53374 => "0111111100110000",
53375 => "0111111100110000",
53376 => "0111111100110000",
53377 => "0111111100110000",
53378 => "0111111100110000",
53379 => "0111111100110000",
53380 => "0111111100110000",
53381 => "0111111100110000",
53382 => "0111111100110000",
53383 => "0111111100110000",
53384 => "0111111100110000",
53385 => "0111111100110000",
53386 => "0111111100110000",
53387 => "0111111100110000",
53388 => "0111111100110000",
53389 => "0111111100110000",
53390 => "0111111100110000",
53391 => "0111111100110000",
53392 => "0111111100110000",
53393 => "0111111100110000",
53394 => "0111111100110000",
53395 => "0111111100110000",
53396 => "0111111100110000",
53397 => "0111111100110000",
53398 => "0111111100110000",
53399 => "0111111100110000",
53400 => "0111111100110000",
53401 => "0111111100110000",
53402 => "0111111100110000",
53403 => "0111111100110000",
53404 => "0111111100110000",
53405 => "0111111100110000",
53406 => "0111111100110000",
53407 => "0111111100110000",
53408 => "0111111100110000",
53409 => "0111111100110000",
53410 => "0111111100110000",
53411 => "0111111100110000",
53412 => "0111111100110000",
53413 => "0111111100110000",
53414 => "0111111100110000",
53415 => "0111111100110000",
53416 => "0111111100110000",
53417 => "0111111100110000",
53418 => "0111111100110000",
53419 => "0111111100110000",
53420 => "0111111100110000",
53421 => "0111111100110000",
53422 => "0111111100110000",
53423 => "0111111100110000",
53424 => "0111111100110000",
53425 => "0111111100110000",
53426 => "0111111100110000",
53427 => "0111111100110000",
53428 => "0111111100110000",
53429 => "0111111100110000",
53430 => "0111111100110000",
53431 => "0111111100110000",
53432 => "0111111100110000",
53433 => "0111111100110000",
53434 => "0111111100110000",
53435 => "0111111100110000",
53436 => "0111111100110000",
53437 => "0111111100110000",
53438 => "0111111100110000",
53439 => "0111111100110000",
53440 => "0111111100110000",
53441 => "0111111100110000",
53442 => "0111111100110000",
53443 => "0111111100110000",
53444 => "0111111100110000",
53445 => "0111111100110000",
53446 => "0111111100110000",
53447 => "0111111100110000",
53448 => "0111111100110000",
53449 => "0111111100110000",
53450 => "0111111100110000",
53451 => "0111111100110000",
53452 => "0111111100110000",
53453 => "0111111100110000",
53454 => "0111111100110000",
53455 => "0111111100110000",
53456 => "0111111100110000",
53457 => "0111111100110000",
53458 => "0111111100110000",
53459 => "0111111100110000",
53460 => "0111111100110000",
53461 => "0111111100110000",
53462 => "0111111100110000",
53463 => "0111111100110000",
53464 => "0111111100110000",
53465 => "0111111100110000",
53466 => "0111111100110000",
53467 => "0111111100110000",
53468 => "0111111100110000",
53469 => "0111111100110000",
53470 => "0111111100110000",
53471 => "0111111100110000",
53472 => "0111111100110000",
53473 => "0111111100110000",
53474 => "0111111100110000",
53475 => "0111111100110000",
53476 => "0111111100110000",
53477 => "0111111100110000",
53478 => "0111111100110000",
53479 => "0111111100110000",
53480 => "0111111100110000",
53481 => "0111111100110000",
53482 => "0111111100110000",
53483 => "0111111100110000",
53484 => "0111111100110000",
53485 => "0111111100110000",
53486 => "0111111100110000",
53487 => "0111111100110000",
53488 => "0111111100110000",
53489 => "0111111100110000",
53490 => "0111111100110000",
53491 => "0111111100110000",
53492 => "0111111100110000",
53493 => "0111111100110000",
53494 => "0111111100110000",
53495 => "0111111100110000",
53496 => "0111111100110000",
53497 => "0111111100110000",
53498 => "0111111100110000",
53499 => "0111111100110000",
53500 => "0111111100110000",
53501 => "0111111100110000",
53502 => "0111111100110000",
53503 => "0111111100110000",
53504 => "0111111100110000",
53505 => "0111111100110000",
53506 => "0111111100110000",
53507 => "0111111100110000",
53508 => "0111111100110000",
53509 => "0111111100110000",
53510 => "0111111100110000",
53511 => "0111111100110000",
53512 => "0111111100110000",
53513 => "0111111100110000",
53514 => "0111111100110000",
53515 => "0111111100110000",
53516 => "0111111100110000",
53517 => "0111111100110000",
53518 => "0111111100110000",
53519 => "0111111100110000",
53520 => "0111111100110000",
53521 => "0111111100110000",
53522 => "0111111100110000",
53523 => "0111111100110000",
53524 => "0111111100110000",
53525 => "0111111100110000",
53526 => "0111111100110000",
53527 => "0111111100110000",
53528 => "0111111100110000",
53529 => "0111111100110000",
53530 => "0111111100110000",
53531 => "0111111100110000",
53532 => "0111111100110000",
53533 => "0111111100110000",
53534 => "0111111100110000",
53535 => "0111111100110000",
53536 => "0111111100110000",
53537 => "0111111100110000",
53538 => "0111111100110000",
53539 => "0111111100110000",
53540 => "0111111100110000",
53541 => "0111111100110000",
53542 => "0111111100110000",
53543 => "0111111100110000",
53544 => "0111111100110000",
53545 => "0111111100110000",
53546 => "0111111100110000",
53547 => "0111111100110000",
53548 => "0111111100110000",
53549 => "0111111100110000",
53550 => "0111111100110000",
53551 => "0111111100110000",
53552 => "0111111100110000",
53553 => "0111111100110000",
53554 => "0111111100110000",
53555 => "0111111100110000",
53556 => "0111111100110000",
53557 => "0111111100110000",
53558 => "0111111100110000",
53559 => "0111111100110000",
53560 => "0111111100110000",
53561 => "0111111100110000",
53562 => "0111111100110000",
53563 => "0111111100110000",
53564 => "0111111100110000",
53565 => "0111111100110000",
53566 => "0111111100110000",
53567 => "0111111100110000",
53568 => "0111111100110000",
53569 => "0111111100110000",
53570 => "0111111100110000",
53571 => "0111111100110000",
53572 => "0111111100110000",
53573 => "0111111100110000",
53574 => "0111111100110000",
53575 => "0111111100110000",
53576 => "0111111100110000",
53577 => "0111111100110000",
53578 => "0111111100110000",
53579 => "0111111100110000",
53580 => "0111111100110000",
53581 => "0111111100110000",
53582 => "0111111100110000",
53583 => "0111111100110000",
53584 => "0111111100110000",
53585 => "0111111100110000",
53586 => "0111111100110000",
53587 => "0111111100110000",
53588 => "0111111100110000",
53589 => "0111111100110000",
53590 => "0111111100110000",
53591 => "0111111100110000",
53592 => "0111111100110000",
53593 => "0111111100110000",
53594 => "0111111100110000",
53595 => "0111111100110000",
53596 => "0111111100110000",
53597 => "0111111100110000",
53598 => "0111111100110000",
53599 => "0111111100110000",
53600 => "0111111100110000",
53601 => "0111111100110000",
53602 => "0111111100110000",
53603 => "0111111100110000",
53604 => "0111111100110000",
53605 => "0111111100110000",
53606 => "0111111100110000",
53607 => "0111111100110000",
53608 => "0111111100110000",
53609 => "0111111100110000",
53610 => "0111111100110000",
53611 => "0111111100110000",
53612 => "0111111100110000",
53613 => "0111111100110000",
53614 => "0111111100110000",
53615 => "0111111100110000",
53616 => "0111111100110000",
53617 => "0111111100110000",
53618 => "0111111100110000",
53619 => "0111111100110000",
53620 => "0111111100110000",
53621 => "0111111100110000",
53622 => "0111111100110000",
53623 => "0111111100110000",
53624 => "0111111100110000",
53625 => "0111111100110000",
53626 => "0111111100110000",
53627 => "0111111100110000",
53628 => "0111111101000000",
53629 => "0111111101000000",
53630 => "0111111101000000",
53631 => "0111111101000000",
53632 => "0111111101000000",
53633 => "0111111101000000",
53634 => "0111111101000000",
53635 => "0111111101000000",
53636 => "0111111101000000",
53637 => "0111111101000000",
53638 => "0111111101000000",
53639 => "0111111101000000",
53640 => "0111111101000000",
53641 => "0111111101000000",
53642 => "0111111101000000",
53643 => "0111111101000000",
53644 => "0111111101000000",
53645 => "0111111101000000",
53646 => "0111111101000000",
53647 => "0111111101000000",
53648 => "0111111101000000",
53649 => "0111111101000000",
53650 => "0111111101000000",
53651 => "0111111101000000",
53652 => "0111111101000000",
53653 => "0111111101000000",
53654 => "0111111101000000",
53655 => "0111111101000000",
53656 => "0111111101000000",
53657 => "0111111101000000",
53658 => "0111111101000000",
53659 => "0111111101000000",
53660 => "0111111101000000",
53661 => "0111111101000000",
53662 => "0111111101000000",
53663 => "0111111101000000",
53664 => "0111111101000000",
53665 => "0111111101000000",
53666 => "0111111101000000",
53667 => "0111111101000000",
53668 => "0111111101000000",
53669 => "0111111101000000",
53670 => "0111111101000000",
53671 => "0111111101000000",
53672 => "0111111101000000",
53673 => "0111111101000000",
53674 => "0111111101000000",
53675 => "0111111101000000",
53676 => "0111111101000000",
53677 => "0111111101000000",
53678 => "0111111101000000",
53679 => "0111111101000000",
53680 => "0111111101000000",
53681 => "0111111101000000",
53682 => "0111111101000000",
53683 => "0111111101000000",
53684 => "0111111101000000",
53685 => "0111111101000000",
53686 => "0111111101000000",
53687 => "0111111101000000",
53688 => "0111111101000000",
53689 => "0111111101000000",
53690 => "0111111101000000",
53691 => "0111111101000000",
53692 => "0111111101000000",
53693 => "0111111101000000",
53694 => "0111111101000000",
53695 => "0111111101000000",
53696 => "0111111101000000",
53697 => "0111111101000000",
53698 => "0111111101000000",
53699 => "0111111101000000",
53700 => "0111111101000000",
53701 => "0111111101000000",
53702 => "0111111101000000",
53703 => "0111111101000000",
53704 => "0111111101000000",
53705 => "0111111101000000",
53706 => "0111111101000000",
53707 => "0111111101000000",
53708 => "0111111101000000",
53709 => "0111111101000000",
53710 => "0111111101000000",
53711 => "0111111101000000",
53712 => "0111111101000000",
53713 => "0111111101000000",
53714 => "0111111101000000",
53715 => "0111111101000000",
53716 => "0111111101000000",
53717 => "0111111101000000",
53718 => "0111111101000000",
53719 => "0111111101000000",
53720 => "0111111101000000",
53721 => "0111111101000000",
53722 => "0111111101000000",
53723 => "0111111101000000",
53724 => "0111111101000000",
53725 => "0111111101000000",
53726 => "0111111101000000",
53727 => "0111111101000000",
53728 => "0111111101000000",
53729 => "0111111101000000",
53730 => "0111111101000000",
53731 => "0111111101000000",
53732 => "0111111101000000",
53733 => "0111111101000000",
53734 => "0111111101000000",
53735 => "0111111101000000",
53736 => "0111111101000000",
53737 => "0111111101000000",
53738 => "0111111101000000",
53739 => "0111111101000000",
53740 => "0111111101000000",
53741 => "0111111101000000",
53742 => "0111111101000000",
53743 => "0111111101000000",
53744 => "0111111101000000",
53745 => "0111111101000000",
53746 => "0111111101000000",
53747 => "0111111101000000",
53748 => "0111111101000000",
53749 => "0111111101000000",
53750 => "0111111101000000",
53751 => "0111111101000000",
53752 => "0111111101000000",
53753 => "0111111101000000",
53754 => "0111111101000000",
53755 => "0111111101000000",
53756 => "0111111101000000",
53757 => "0111111101000000",
53758 => "0111111101000000",
53759 => "0111111101000000",
53760 => "0111111101000000",
53761 => "0111111101000000",
53762 => "0111111101000000",
53763 => "0111111101000000",
53764 => "0111111101000000",
53765 => "0111111101000000",
53766 => "0111111101000000",
53767 => "0111111101000000",
53768 => "0111111101000000",
53769 => "0111111101000000",
53770 => "0111111101000000",
53771 => "0111111101000000",
53772 => "0111111101000000",
53773 => "0111111101000000",
53774 => "0111111101000000",
53775 => "0111111101000000",
53776 => "0111111101000000",
53777 => "0111111101000000",
53778 => "0111111101000000",
53779 => "0111111101000000",
53780 => "0111111101000000",
53781 => "0111111101000000",
53782 => "0111111101000000",
53783 => "0111111101000000",
53784 => "0111111101000000",
53785 => "0111111101000000",
53786 => "0111111101000000",
53787 => "0111111101000000",
53788 => "0111111101000000",
53789 => "0111111101000000",
53790 => "0111111101000000",
53791 => "0111111101000000",
53792 => "0111111101000000",
53793 => "0111111101000000",
53794 => "0111111101000000",
53795 => "0111111101000000",
53796 => "0111111101000000",
53797 => "0111111101000000",
53798 => "0111111101000000",
53799 => "0111111101000000",
53800 => "0111111101000000",
53801 => "0111111101000000",
53802 => "0111111101000000",
53803 => "0111111101000000",
53804 => "0111111101000000",
53805 => "0111111101000000",
53806 => "0111111101000000",
53807 => "0111111101000000",
53808 => "0111111101000000",
53809 => "0111111101000000",
53810 => "0111111101000000",
53811 => "0111111101000000",
53812 => "0111111101000000",
53813 => "0111111101000000",
53814 => "0111111101000000",
53815 => "0111111101000000",
53816 => "0111111101000000",
53817 => "0111111101000000",
53818 => "0111111101000000",
53819 => "0111111101000000",
53820 => "0111111101000000",
53821 => "0111111101000000",
53822 => "0111111101000000",
53823 => "0111111101000000",
53824 => "0111111101000000",
53825 => "0111111101000000",
53826 => "0111111101000000",
53827 => "0111111101000000",
53828 => "0111111101000000",
53829 => "0111111101000000",
53830 => "0111111101000000",
53831 => "0111111101000000",
53832 => "0111111101000000",
53833 => "0111111101000000",
53834 => "0111111101000000",
53835 => "0111111101000000",
53836 => "0111111101000000",
53837 => "0111111101000000",
53838 => "0111111101000000",
53839 => "0111111101000000",
53840 => "0111111101000000",
53841 => "0111111101000000",
53842 => "0111111101000000",
53843 => "0111111101000000",
53844 => "0111111101000000",
53845 => "0111111101000000",
53846 => "0111111101000000",
53847 => "0111111101000000",
53848 => "0111111101000000",
53849 => "0111111101000000",
53850 => "0111111101000000",
53851 => "0111111101000000",
53852 => "0111111101000000",
53853 => "0111111101000000",
53854 => "0111111101000000",
53855 => "0111111101000000",
53856 => "0111111101000000",
53857 => "0111111101000000",
53858 => "0111111101000000",
53859 => "0111111101000000",
53860 => "0111111101000000",
53861 => "0111111101000000",
53862 => "0111111101000000",
53863 => "0111111101000000",
53864 => "0111111101000000",
53865 => "0111111101000000",
53866 => "0111111101000000",
53867 => "0111111101000000",
53868 => "0111111101000000",
53869 => "0111111101000000",
53870 => "0111111101000000",
53871 => "0111111101000000",
53872 => "0111111101000000",
53873 => "0111111101000000",
53874 => "0111111101000000",
53875 => "0111111101000000",
53876 => "0111111101000000",
53877 => "0111111101000000",
53878 => "0111111101000000",
53879 => "0111111101000000",
53880 => "0111111101000000",
53881 => "0111111101000000",
53882 => "0111111101000000",
53883 => "0111111101000000",
53884 => "0111111101000000",
53885 => "0111111101000000",
53886 => "0111111101000000",
53887 => "0111111101000000",
53888 => "0111111101000000",
53889 => "0111111101000000",
53890 => "0111111101000000",
53891 => "0111111101000000",
53892 => "0111111101000000",
53893 => "0111111101000000",
53894 => "0111111101000000",
53895 => "0111111101000000",
53896 => "0111111101000000",
53897 => "0111111101000000",
53898 => "0111111101000000",
53899 => "0111111101000000",
53900 => "0111111101000000",
53901 => "0111111101000000",
53902 => "0111111101000000",
53903 => "0111111101000000",
53904 => "0111111101000000",
53905 => "0111111101000000",
53906 => "0111111101000000",
53907 => "0111111101000000",
53908 => "0111111101000000",
53909 => "0111111101000000",
53910 => "0111111101000000",
53911 => "0111111101000000",
53912 => "0111111101000000",
53913 => "0111111101000000",
53914 => "0111111101000000",
53915 => "0111111101000000",
53916 => "0111111101000000",
53917 => "0111111101000000",
53918 => "0111111101000000",
53919 => "0111111101000000",
53920 => "0111111101000000",
53921 => "0111111101000000",
53922 => "0111111101000000",
53923 => "0111111101000000",
53924 => "0111111101000000",
53925 => "0111111101000000",
53926 => "0111111101000000",
53927 => "0111111101000000",
53928 => "0111111101000000",
53929 => "0111111101000000",
53930 => "0111111101000000",
53931 => "0111111101000000",
53932 => "0111111101000000",
53933 => "0111111101000000",
53934 => "0111111101000000",
53935 => "0111111101000000",
53936 => "0111111101000000",
53937 => "0111111101000000",
53938 => "0111111101000000",
53939 => "0111111101000000",
53940 => "0111111101000000",
53941 => "0111111101000000",
53942 => "0111111101000000",
53943 => "0111111101000000",
53944 => "0111111101000000",
53945 => "0111111101000000",
53946 => "0111111101000000",
53947 => "0111111101000000",
53948 => "0111111101000000",
53949 => "0111111101000000",
53950 => "0111111101000000",
53951 => "0111111101000000",
53952 => "0111111101000000",
53953 => "0111111101000000",
53954 => "0111111101000000",
53955 => "0111111101000000",
53956 => "0111111101000000",
53957 => "0111111101000000",
53958 => "0111111101000000",
53959 => "0111111101000000",
53960 => "0111111101000000",
53961 => "0111111101000000",
53962 => "0111111101000000",
53963 => "0111111101000000",
53964 => "0111111101000000",
53965 => "0111111101000000",
53966 => "0111111101000000",
53967 => "0111111101000000",
53968 => "0111111101000000",
53969 => "0111111101000000",
53970 => "0111111101000000",
53971 => "0111111101010000",
53972 => "0111111101010000",
53973 => "0111111101010000",
53974 => "0111111101010000",
53975 => "0111111101010000",
53976 => "0111111101010000",
53977 => "0111111101010000",
53978 => "0111111101010000",
53979 => "0111111101010000",
53980 => "0111111101010000",
53981 => "0111111101010000",
53982 => "0111111101010000",
53983 => "0111111101010000",
53984 => "0111111101010000",
53985 => "0111111101010000",
53986 => "0111111101010000",
53987 => "0111111101010000",
53988 => "0111111101010000",
53989 => "0111111101010000",
53990 => "0111111101010000",
53991 => "0111111101010000",
53992 => "0111111101010000",
53993 => "0111111101010000",
53994 => "0111111101010000",
53995 => "0111111101010000",
53996 => "0111111101010000",
53997 => "0111111101010000",
53998 => "0111111101010000",
53999 => "0111111101010000",
54000 => "0111111101010000",
54001 => "0111111101010000",
54002 => "0111111101010000",
54003 => "0111111101010000",
54004 => "0111111101010000",
54005 => "0111111101010000",
54006 => "0111111101010000",
54007 => "0111111101010000",
54008 => "0111111101010000",
54009 => "0111111101010000",
54010 => "0111111101010000",
54011 => "0111111101010000",
54012 => "0111111101010000",
54013 => "0111111101010000",
54014 => "0111111101010000",
54015 => "0111111101010000",
54016 => "0111111101010000",
54017 => "0111111101010000",
54018 => "0111111101010000",
54019 => "0111111101010000",
54020 => "0111111101010000",
54021 => "0111111101010000",
54022 => "0111111101010000",
54023 => "0111111101010000",
54024 => "0111111101010000",
54025 => "0111111101010000",
54026 => "0111111101010000",
54027 => "0111111101010000",
54028 => "0111111101010000",
54029 => "0111111101010000",
54030 => "0111111101010000",
54031 => "0111111101010000",
54032 => "0111111101010000",
54033 => "0111111101010000",
54034 => "0111111101010000",
54035 => "0111111101010000",
54036 => "0111111101010000",
54037 => "0111111101010000",
54038 => "0111111101010000",
54039 => "0111111101010000",
54040 => "0111111101010000",
54041 => "0111111101010000",
54042 => "0111111101010000",
54043 => "0111111101010000",
54044 => "0111111101010000",
54045 => "0111111101010000",
54046 => "0111111101010000",
54047 => "0111111101010000",
54048 => "0111111101010000",
54049 => "0111111101010000",
54050 => "0111111101010000",
54051 => "0111111101010000",
54052 => "0111111101010000",
54053 => "0111111101010000",
54054 => "0111111101010000",
54055 => "0111111101010000",
54056 => "0111111101010000",
54057 => "0111111101010000",
54058 => "0111111101010000",
54059 => "0111111101010000",
54060 => "0111111101010000",
54061 => "0111111101010000",
54062 => "0111111101010000",
54063 => "0111111101010000",
54064 => "0111111101010000",
54065 => "0111111101010000",
54066 => "0111111101010000",
54067 => "0111111101010000",
54068 => "0111111101010000",
54069 => "0111111101010000",
54070 => "0111111101010000",
54071 => "0111111101010000",
54072 => "0111111101010000",
54073 => "0111111101010000",
54074 => "0111111101010000",
54075 => "0111111101010000",
54076 => "0111111101010000",
54077 => "0111111101010000",
54078 => "0111111101010000",
54079 => "0111111101010000",
54080 => "0111111101010000",
54081 => "0111111101010000",
54082 => "0111111101010000",
54083 => "0111111101010000",
54084 => "0111111101010000",
54085 => "0111111101010000",
54086 => "0111111101010000",
54087 => "0111111101010000",
54088 => "0111111101010000",
54089 => "0111111101010000",
54090 => "0111111101010000",
54091 => "0111111101010000",
54092 => "0111111101010000",
54093 => "0111111101010000",
54094 => "0111111101010000",
54095 => "0111111101010000",
54096 => "0111111101010000",
54097 => "0111111101010000",
54098 => "0111111101010000",
54099 => "0111111101010000",
54100 => "0111111101010000",
54101 => "0111111101010000",
54102 => "0111111101010000",
54103 => "0111111101010000",
54104 => "0111111101010000",
54105 => "0111111101010000",
54106 => "0111111101010000",
54107 => "0111111101010000",
54108 => "0111111101010000",
54109 => "0111111101010000",
54110 => "0111111101010000",
54111 => "0111111101010000",
54112 => "0111111101010000",
54113 => "0111111101010000",
54114 => "0111111101010000",
54115 => "0111111101010000",
54116 => "0111111101010000",
54117 => "0111111101010000",
54118 => "0111111101010000",
54119 => "0111111101010000",
54120 => "0111111101010000",
54121 => "0111111101010000",
54122 => "0111111101010000",
54123 => "0111111101010000",
54124 => "0111111101010000",
54125 => "0111111101010000",
54126 => "0111111101010000",
54127 => "0111111101010000",
54128 => "0111111101010000",
54129 => "0111111101010000",
54130 => "0111111101010000",
54131 => "0111111101010000",
54132 => "0111111101010000",
54133 => "0111111101010000",
54134 => "0111111101010000",
54135 => "0111111101010000",
54136 => "0111111101010000",
54137 => "0111111101010000",
54138 => "0111111101010000",
54139 => "0111111101010000",
54140 => "0111111101010000",
54141 => "0111111101010000",
54142 => "0111111101010000",
54143 => "0111111101010000",
54144 => "0111111101010000",
54145 => "0111111101010000",
54146 => "0111111101010000",
54147 => "0111111101010000",
54148 => "0111111101010000",
54149 => "0111111101010000",
54150 => "0111111101010000",
54151 => "0111111101010000",
54152 => "0111111101010000",
54153 => "0111111101010000",
54154 => "0111111101010000",
54155 => "0111111101010000",
54156 => "0111111101010000",
54157 => "0111111101010000",
54158 => "0111111101010000",
54159 => "0111111101010000",
54160 => "0111111101010000",
54161 => "0111111101010000",
54162 => "0111111101010000",
54163 => "0111111101010000",
54164 => "0111111101010000",
54165 => "0111111101010000",
54166 => "0111111101010000",
54167 => "0111111101010000",
54168 => "0111111101010000",
54169 => "0111111101010000",
54170 => "0111111101010000",
54171 => "0111111101010000",
54172 => "0111111101010000",
54173 => "0111111101010000",
54174 => "0111111101010000",
54175 => "0111111101010000",
54176 => "0111111101010000",
54177 => "0111111101010000",
54178 => "0111111101010000",
54179 => "0111111101010000",
54180 => "0111111101010000",
54181 => "0111111101010000",
54182 => "0111111101010000",
54183 => "0111111101010000",
54184 => "0111111101010000",
54185 => "0111111101010000",
54186 => "0111111101010000",
54187 => "0111111101010000",
54188 => "0111111101010000",
54189 => "0111111101010000",
54190 => "0111111101010000",
54191 => "0111111101010000",
54192 => "0111111101010000",
54193 => "0111111101010000",
54194 => "0111111101010000",
54195 => "0111111101010000",
54196 => "0111111101010000",
54197 => "0111111101010000",
54198 => "0111111101010000",
54199 => "0111111101010000",
54200 => "0111111101010000",
54201 => "0111111101010000",
54202 => "0111111101010000",
54203 => "0111111101010000",
54204 => "0111111101010000",
54205 => "0111111101010000",
54206 => "0111111101010000",
54207 => "0111111101010000",
54208 => "0111111101010000",
54209 => "0111111101010000",
54210 => "0111111101010000",
54211 => "0111111101010000",
54212 => "0111111101010000",
54213 => "0111111101010000",
54214 => "0111111101010000",
54215 => "0111111101010000",
54216 => "0111111101010000",
54217 => "0111111101010000",
54218 => "0111111101010000",
54219 => "0111111101010000",
54220 => "0111111101010000",
54221 => "0111111101010000",
54222 => "0111111101010000",
54223 => "0111111101010000",
54224 => "0111111101010000",
54225 => "0111111101010000",
54226 => "0111111101010000",
54227 => "0111111101010000",
54228 => "0111111101010000",
54229 => "0111111101010000",
54230 => "0111111101010000",
54231 => "0111111101010000",
54232 => "0111111101010000",
54233 => "0111111101010000",
54234 => "0111111101010000",
54235 => "0111111101010000",
54236 => "0111111101010000",
54237 => "0111111101010000",
54238 => "0111111101010000",
54239 => "0111111101010000",
54240 => "0111111101010000",
54241 => "0111111101010000",
54242 => "0111111101010000",
54243 => "0111111101010000",
54244 => "0111111101010000",
54245 => "0111111101010000",
54246 => "0111111101010000",
54247 => "0111111101010000",
54248 => "0111111101010000",
54249 => "0111111101010000",
54250 => "0111111101010000",
54251 => "0111111101010000",
54252 => "0111111101010000",
54253 => "0111111101010000",
54254 => "0111111101010000",
54255 => "0111111101010000",
54256 => "0111111101010000",
54257 => "0111111101010000",
54258 => "0111111101010000",
54259 => "0111111101010000",
54260 => "0111111101010000",
54261 => "0111111101010000",
54262 => "0111111101010000",
54263 => "0111111101010000",
54264 => "0111111101010000",
54265 => "0111111101010000",
54266 => "0111111101010000",
54267 => "0111111101010000",
54268 => "0111111101010000",
54269 => "0111111101010000",
54270 => "0111111101010000",
54271 => "0111111101010000",
54272 => "0111111101010000",
54273 => "0111111101010000",
54274 => "0111111101010000",
54275 => "0111111101010000",
54276 => "0111111101010000",
54277 => "0111111101010000",
54278 => "0111111101010000",
54279 => "0111111101010000",
54280 => "0111111101010000",
54281 => "0111111101010000",
54282 => "0111111101010000",
54283 => "0111111101010000",
54284 => "0111111101010000",
54285 => "0111111101010000",
54286 => "0111111101010000",
54287 => "0111111101010000",
54288 => "0111111101010000",
54289 => "0111111101010000",
54290 => "0111111101010000",
54291 => "0111111101010000",
54292 => "0111111101010000",
54293 => "0111111101010000",
54294 => "0111111101010000",
54295 => "0111111101010000",
54296 => "0111111101010000",
54297 => "0111111101010000",
54298 => "0111111101010000",
54299 => "0111111101010000",
54300 => "0111111101010000",
54301 => "0111111101010000",
54302 => "0111111101010000",
54303 => "0111111101010000",
54304 => "0111111101010000",
54305 => "0111111101010000",
54306 => "0111111101010000",
54307 => "0111111101010000",
54308 => "0111111101010000",
54309 => "0111111101010000",
54310 => "0111111101010000",
54311 => "0111111101010000",
54312 => "0111111101010000",
54313 => "0111111101010000",
54314 => "0111111101010000",
54315 => "0111111101010000",
54316 => "0111111101010000",
54317 => "0111111101010000",
54318 => "0111111101010000",
54319 => "0111111101010000",
54320 => "0111111101010000",
54321 => "0111111101010000",
54322 => "0111111101010000",
54323 => "0111111101010000",
54324 => "0111111101010000",
54325 => "0111111101010000",
54326 => "0111111101010000",
54327 => "0111111101010000",
54328 => "0111111101010000",
54329 => "0111111101010000",
54330 => "0111111101010000",
54331 => "0111111101010000",
54332 => "0111111101010000",
54333 => "0111111101010000",
54334 => "0111111101010000",
54335 => "0111111101010000",
54336 => "0111111101010000",
54337 => "0111111101010000",
54338 => "0111111101010000",
54339 => "0111111101010000",
54340 => "0111111101010000",
54341 => "0111111101010000",
54342 => "0111111101010000",
54343 => "0111111101010000",
54344 => "0111111101010000",
54345 => "0111111101010000",
54346 => "0111111101100000",
54347 => "0111111101100000",
54348 => "0111111101100000",
54349 => "0111111101100000",
54350 => "0111111101100000",
54351 => "0111111101100000",
54352 => "0111111101100000",
54353 => "0111111101100000",
54354 => "0111111101100000",
54355 => "0111111101100000",
54356 => "0111111101100000",
54357 => "0111111101100000",
54358 => "0111111101100000",
54359 => "0111111101100000",
54360 => "0111111101100000",
54361 => "0111111101100000",
54362 => "0111111101100000",
54363 => "0111111101100000",
54364 => "0111111101100000",
54365 => "0111111101100000",
54366 => "0111111101100000",
54367 => "0111111101100000",
54368 => "0111111101100000",
54369 => "0111111101100000",
54370 => "0111111101100000",
54371 => "0111111101100000",
54372 => "0111111101100000",
54373 => "0111111101100000",
54374 => "0111111101100000",
54375 => "0111111101100000",
54376 => "0111111101100000",
54377 => "0111111101100000",
54378 => "0111111101100000",
54379 => "0111111101100000",
54380 => "0111111101100000",
54381 => "0111111101100000",
54382 => "0111111101100000",
54383 => "0111111101100000",
54384 => "0111111101100000",
54385 => "0111111101100000",
54386 => "0111111101100000",
54387 => "0111111101100000",
54388 => "0111111101100000",
54389 => "0111111101100000",
54390 => "0111111101100000",
54391 => "0111111101100000",
54392 => "0111111101100000",
54393 => "0111111101100000",
54394 => "0111111101100000",
54395 => "0111111101100000",
54396 => "0111111101100000",
54397 => "0111111101100000",
54398 => "0111111101100000",
54399 => "0111111101100000",
54400 => "0111111101100000",
54401 => "0111111101100000",
54402 => "0111111101100000",
54403 => "0111111101100000",
54404 => "0111111101100000",
54405 => "0111111101100000",
54406 => "0111111101100000",
54407 => "0111111101100000",
54408 => "0111111101100000",
54409 => "0111111101100000",
54410 => "0111111101100000",
54411 => "0111111101100000",
54412 => "0111111101100000",
54413 => "0111111101100000",
54414 => "0111111101100000",
54415 => "0111111101100000",
54416 => "0111111101100000",
54417 => "0111111101100000",
54418 => "0111111101100000",
54419 => "0111111101100000",
54420 => "0111111101100000",
54421 => "0111111101100000",
54422 => "0111111101100000",
54423 => "0111111101100000",
54424 => "0111111101100000",
54425 => "0111111101100000",
54426 => "0111111101100000",
54427 => "0111111101100000",
54428 => "0111111101100000",
54429 => "0111111101100000",
54430 => "0111111101100000",
54431 => "0111111101100000",
54432 => "0111111101100000",
54433 => "0111111101100000",
54434 => "0111111101100000",
54435 => "0111111101100000",
54436 => "0111111101100000",
54437 => "0111111101100000",
54438 => "0111111101100000",
54439 => "0111111101100000",
54440 => "0111111101100000",
54441 => "0111111101100000",
54442 => "0111111101100000",
54443 => "0111111101100000",
54444 => "0111111101100000",
54445 => "0111111101100000",
54446 => "0111111101100000",
54447 => "0111111101100000",
54448 => "0111111101100000",
54449 => "0111111101100000",
54450 => "0111111101100000",
54451 => "0111111101100000",
54452 => "0111111101100000",
54453 => "0111111101100000",
54454 => "0111111101100000",
54455 => "0111111101100000",
54456 => "0111111101100000",
54457 => "0111111101100000",
54458 => "0111111101100000",
54459 => "0111111101100000",
54460 => "0111111101100000",
54461 => "0111111101100000",
54462 => "0111111101100000",
54463 => "0111111101100000",
54464 => "0111111101100000",
54465 => "0111111101100000",
54466 => "0111111101100000",
54467 => "0111111101100000",
54468 => "0111111101100000",
54469 => "0111111101100000",
54470 => "0111111101100000",
54471 => "0111111101100000",
54472 => "0111111101100000",
54473 => "0111111101100000",
54474 => "0111111101100000",
54475 => "0111111101100000",
54476 => "0111111101100000",
54477 => "0111111101100000",
54478 => "0111111101100000",
54479 => "0111111101100000",
54480 => "0111111101100000",
54481 => "0111111101100000",
54482 => "0111111101100000",
54483 => "0111111101100000",
54484 => "0111111101100000",
54485 => "0111111101100000",
54486 => "0111111101100000",
54487 => "0111111101100000",
54488 => "0111111101100000",
54489 => "0111111101100000",
54490 => "0111111101100000",
54491 => "0111111101100000",
54492 => "0111111101100000",
54493 => "0111111101100000",
54494 => "0111111101100000",
54495 => "0111111101100000",
54496 => "0111111101100000",
54497 => "0111111101100000",
54498 => "0111111101100000",
54499 => "0111111101100000",
54500 => "0111111101100000",
54501 => "0111111101100000",
54502 => "0111111101100000",
54503 => "0111111101100000",
54504 => "0111111101100000",
54505 => "0111111101100000",
54506 => "0111111101100000",
54507 => "0111111101100000",
54508 => "0111111101100000",
54509 => "0111111101100000",
54510 => "0111111101100000",
54511 => "0111111101100000",
54512 => "0111111101100000",
54513 => "0111111101100000",
54514 => "0111111101100000",
54515 => "0111111101100000",
54516 => "0111111101100000",
54517 => "0111111101100000",
54518 => "0111111101100000",
54519 => "0111111101100000",
54520 => "0111111101100000",
54521 => "0111111101100000",
54522 => "0111111101100000",
54523 => "0111111101100000",
54524 => "0111111101100000",
54525 => "0111111101100000",
54526 => "0111111101100000",
54527 => "0111111101100000",
54528 => "0111111101100000",
54529 => "0111111101100000",
54530 => "0111111101100000",
54531 => "0111111101100000",
54532 => "0111111101100000",
54533 => "0111111101100000",
54534 => "0111111101100000",
54535 => "0111111101100000",
54536 => "0111111101100000",
54537 => "0111111101100000",
54538 => "0111111101100000",
54539 => "0111111101100000",
54540 => "0111111101100000",
54541 => "0111111101100000",
54542 => "0111111101100000",
54543 => "0111111101100000",
54544 => "0111111101100000",
54545 => "0111111101100000",
54546 => "0111111101100000",
54547 => "0111111101100000",
54548 => "0111111101100000",
54549 => "0111111101100000",
54550 => "0111111101100000",
54551 => "0111111101100000",
54552 => "0111111101100000",
54553 => "0111111101100000",
54554 => "0111111101100000",
54555 => "0111111101100000",
54556 => "0111111101100000",
54557 => "0111111101100000",
54558 => "0111111101100000",
54559 => "0111111101100000",
54560 => "0111111101100000",
54561 => "0111111101100000",
54562 => "0111111101100000",
54563 => "0111111101100000",
54564 => "0111111101100000",
54565 => "0111111101100000",
54566 => "0111111101100000",
54567 => "0111111101100000",
54568 => "0111111101100000",
54569 => "0111111101100000",
54570 => "0111111101100000",
54571 => "0111111101100000",
54572 => "0111111101100000",
54573 => "0111111101100000",
54574 => "0111111101100000",
54575 => "0111111101100000",
54576 => "0111111101100000",
54577 => "0111111101100000",
54578 => "0111111101100000",
54579 => "0111111101100000",
54580 => "0111111101100000",
54581 => "0111111101100000",
54582 => "0111111101100000",
54583 => "0111111101100000",
54584 => "0111111101100000",
54585 => "0111111101100000",
54586 => "0111111101100000",
54587 => "0111111101100000",
54588 => "0111111101100000",
54589 => "0111111101100000",
54590 => "0111111101100000",
54591 => "0111111101100000",
54592 => "0111111101100000",
54593 => "0111111101100000",
54594 => "0111111101100000",
54595 => "0111111101100000",
54596 => "0111111101100000",
54597 => "0111111101100000",
54598 => "0111111101100000",
54599 => "0111111101100000",
54600 => "0111111101100000",
54601 => "0111111101100000",
54602 => "0111111101100000",
54603 => "0111111101100000",
54604 => "0111111101100000",
54605 => "0111111101100000",
54606 => "0111111101100000",
54607 => "0111111101100000",
54608 => "0111111101100000",
54609 => "0111111101100000",
54610 => "0111111101100000",
54611 => "0111111101100000",
54612 => "0111111101100000",
54613 => "0111111101100000",
54614 => "0111111101100000",
54615 => "0111111101100000",
54616 => "0111111101100000",
54617 => "0111111101100000",
54618 => "0111111101100000",
54619 => "0111111101100000",
54620 => "0111111101100000",
54621 => "0111111101100000",
54622 => "0111111101100000",
54623 => "0111111101100000",
54624 => "0111111101100000",
54625 => "0111111101100000",
54626 => "0111111101100000",
54627 => "0111111101100000",
54628 => "0111111101100000",
54629 => "0111111101100000",
54630 => "0111111101100000",
54631 => "0111111101100000",
54632 => "0111111101100000",
54633 => "0111111101100000",
54634 => "0111111101100000",
54635 => "0111111101100000",
54636 => "0111111101100000",
54637 => "0111111101100000",
54638 => "0111111101100000",
54639 => "0111111101100000",
54640 => "0111111101100000",
54641 => "0111111101100000",
54642 => "0111111101100000",
54643 => "0111111101100000",
54644 => "0111111101100000",
54645 => "0111111101100000",
54646 => "0111111101100000",
54647 => "0111111101100000",
54648 => "0111111101100000",
54649 => "0111111101100000",
54650 => "0111111101100000",
54651 => "0111111101100000",
54652 => "0111111101100000",
54653 => "0111111101100000",
54654 => "0111111101100000",
54655 => "0111111101100000",
54656 => "0111111101100000",
54657 => "0111111101100000",
54658 => "0111111101100000",
54659 => "0111111101100000",
54660 => "0111111101100000",
54661 => "0111111101100000",
54662 => "0111111101100000",
54663 => "0111111101100000",
54664 => "0111111101100000",
54665 => "0111111101100000",
54666 => "0111111101100000",
54667 => "0111111101100000",
54668 => "0111111101100000",
54669 => "0111111101100000",
54670 => "0111111101100000",
54671 => "0111111101100000",
54672 => "0111111101100000",
54673 => "0111111101100000",
54674 => "0111111101100000",
54675 => "0111111101100000",
54676 => "0111111101100000",
54677 => "0111111101100000",
54678 => "0111111101100000",
54679 => "0111111101100000",
54680 => "0111111101100000",
54681 => "0111111101100000",
54682 => "0111111101100000",
54683 => "0111111101100000",
54684 => "0111111101100000",
54685 => "0111111101100000",
54686 => "0111111101100000",
54687 => "0111111101100000",
54688 => "0111111101100000",
54689 => "0111111101100000",
54690 => "0111111101100000",
54691 => "0111111101100000",
54692 => "0111111101100000",
54693 => "0111111101100000",
54694 => "0111111101100000",
54695 => "0111111101100000",
54696 => "0111111101100000",
54697 => "0111111101100000",
54698 => "0111111101100000",
54699 => "0111111101100000",
54700 => "0111111101100000",
54701 => "0111111101100000",
54702 => "0111111101100000",
54703 => "0111111101100000",
54704 => "0111111101100000",
54705 => "0111111101100000",
54706 => "0111111101100000",
54707 => "0111111101100000",
54708 => "0111111101100000",
54709 => "0111111101100000",
54710 => "0111111101100000",
54711 => "0111111101100000",
54712 => "0111111101100000",
54713 => "0111111101100000",
54714 => "0111111101100000",
54715 => "0111111101100000",
54716 => "0111111101100000",
54717 => "0111111101100000",
54718 => "0111111101100000",
54719 => "0111111101100000",
54720 => "0111111101100000",
54721 => "0111111101100000",
54722 => "0111111101100000",
54723 => "0111111101100000",
54724 => "0111111101100000",
54725 => "0111111101100000",
54726 => "0111111101100000",
54727 => "0111111101100000",
54728 => "0111111101100000",
54729 => "0111111101100000",
54730 => "0111111101100000",
54731 => "0111111101100000",
54732 => "0111111101100000",
54733 => "0111111101100000",
54734 => "0111111101100000",
54735 => "0111111101100000",
54736 => "0111111101100000",
54737 => "0111111101100000",
54738 => "0111111101100000",
54739 => "0111111101100000",
54740 => "0111111101100000",
54741 => "0111111101100000",
54742 => "0111111101100000",
54743 => "0111111101100000",
54744 => "0111111101100000",
54745 => "0111111101100000",
54746 => "0111111101100000",
54747 => "0111111101100000",
54748 => "0111111101100000",
54749 => "0111111101100000",
54750 => "0111111101100000",
54751 => "0111111101100000",
54752 => "0111111101100000",
54753 => "0111111101100000",
54754 => "0111111101100000",
54755 => "0111111101100000",
54756 => "0111111101100000",
54757 => "0111111101100000",
54758 => "0111111101110000",
54759 => "0111111101110000",
54760 => "0111111101110000",
54761 => "0111111101110000",
54762 => "0111111101110000",
54763 => "0111111101110000",
54764 => "0111111101110000",
54765 => "0111111101110000",
54766 => "0111111101110000",
54767 => "0111111101110000",
54768 => "0111111101110000",
54769 => "0111111101110000",
54770 => "0111111101110000",
54771 => "0111111101110000",
54772 => "0111111101110000",
54773 => "0111111101110000",
54774 => "0111111101110000",
54775 => "0111111101110000",
54776 => "0111111101110000",
54777 => "0111111101110000",
54778 => "0111111101110000",
54779 => "0111111101110000",
54780 => "0111111101110000",
54781 => "0111111101110000",
54782 => "0111111101110000",
54783 => "0111111101110000",
54784 => "0111111101110000",
54785 => "0111111101110000",
54786 => "0111111101110000",
54787 => "0111111101110000",
54788 => "0111111101110000",
54789 => "0111111101110000",
54790 => "0111111101110000",
54791 => "0111111101110000",
54792 => "0111111101110000",
54793 => "0111111101110000",
54794 => "0111111101110000",
54795 => "0111111101110000",
54796 => "0111111101110000",
54797 => "0111111101110000",
54798 => "0111111101110000",
54799 => "0111111101110000",
54800 => "0111111101110000",
54801 => "0111111101110000",
54802 => "0111111101110000",
54803 => "0111111101110000",
54804 => "0111111101110000",
54805 => "0111111101110000",
54806 => "0111111101110000",
54807 => "0111111101110000",
54808 => "0111111101110000",
54809 => "0111111101110000",
54810 => "0111111101110000",
54811 => "0111111101110000",
54812 => "0111111101110000",
54813 => "0111111101110000",
54814 => "0111111101110000",
54815 => "0111111101110000",
54816 => "0111111101110000",
54817 => "0111111101110000",
54818 => "0111111101110000",
54819 => "0111111101110000",
54820 => "0111111101110000",
54821 => "0111111101110000",
54822 => "0111111101110000",
54823 => "0111111101110000",
54824 => "0111111101110000",
54825 => "0111111101110000",
54826 => "0111111101110000",
54827 => "0111111101110000",
54828 => "0111111101110000",
54829 => "0111111101110000",
54830 => "0111111101110000",
54831 => "0111111101110000",
54832 => "0111111101110000",
54833 => "0111111101110000",
54834 => "0111111101110000",
54835 => "0111111101110000",
54836 => "0111111101110000",
54837 => "0111111101110000",
54838 => "0111111101110000",
54839 => "0111111101110000",
54840 => "0111111101110000",
54841 => "0111111101110000",
54842 => "0111111101110000",
54843 => "0111111101110000",
54844 => "0111111101110000",
54845 => "0111111101110000",
54846 => "0111111101110000",
54847 => "0111111101110000",
54848 => "0111111101110000",
54849 => "0111111101110000",
54850 => "0111111101110000",
54851 => "0111111101110000",
54852 => "0111111101110000",
54853 => "0111111101110000",
54854 => "0111111101110000",
54855 => "0111111101110000",
54856 => "0111111101110000",
54857 => "0111111101110000",
54858 => "0111111101110000",
54859 => "0111111101110000",
54860 => "0111111101110000",
54861 => "0111111101110000",
54862 => "0111111101110000",
54863 => "0111111101110000",
54864 => "0111111101110000",
54865 => "0111111101110000",
54866 => "0111111101110000",
54867 => "0111111101110000",
54868 => "0111111101110000",
54869 => "0111111101110000",
54870 => "0111111101110000",
54871 => "0111111101110000",
54872 => "0111111101110000",
54873 => "0111111101110000",
54874 => "0111111101110000",
54875 => "0111111101110000",
54876 => "0111111101110000",
54877 => "0111111101110000",
54878 => "0111111101110000",
54879 => "0111111101110000",
54880 => "0111111101110000",
54881 => "0111111101110000",
54882 => "0111111101110000",
54883 => "0111111101110000",
54884 => "0111111101110000",
54885 => "0111111101110000",
54886 => "0111111101110000",
54887 => "0111111101110000",
54888 => "0111111101110000",
54889 => "0111111101110000",
54890 => "0111111101110000",
54891 => "0111111101110000",
54892 => "0111111101110000",
54893 => "0111111101110000",
54894 => "0111111101110000",
54895 => "0111111101110000",
54896 => "0111111101110000",
54897 => "0111111101110000",
54898 => "0111111101110000",
54899 => "0111111101110000",
54900 => "0111111101110000",
54901 => "0111111101110000",
54902 => "0111111101110000",
54903 => "0111111101110000",
54904 => "0111111101110000",
54905 => "0111111101110000",
54906 => "0111111101110000",
54907 => "0111111101110000",
54908 => "0111111101110000",
54909 => "0111111101110000",
54910 => "0111111101110000",
54911 => "0111111101110000",
54912 => "0111111101110000",
54913 => "0111111101110000",
54914 => "0111111101110000",
54915 => "0111111101110000",
54916 => "0111111101110000",
54917 => "0111111101110000",
54918 => "0111111101110000",
54919 => "0111111101110000",
54920 => "0111111101110000",
54921 => "0111111101110000",
54922 => "0111111101110000",
54923 => "0111111101110000",
54924 => "0111111101110000",
54925 => "0111111101110000",
54926 => "0111111101110000",
54927 => "0111111101110000",
54928 => "0111111101110000",
54929 => "0111111101110000",
54930 => "0111111101110000",
54931 => "0111111101110000",
54932 => "0111111101110000",
54933 => "0111111101110000",
54934 => "0111111101110000",
54935 => "0111111101110000",
54936 => "0111111101110000",
54937 => "0111111101110000",
54938 => "0111111101110000",
54939 => "0111111101110000",
54940 => "0111111101110000",
54941 => "0111111101110000",
54942 => "0111111101110000",
54943 => "0111111101110000",
54944 => "0111111101110000",
54945 => "0111111101110000",
54946 => "0111111101110000",
54947 => "0111111101110000",
54948 => "0111111101110000",
54949 => "0111111101110000",
54950 => "0111111101110000",
54951 => "0111111101110000",
54952 => "0111111101110000",
54953 => "0111111101110000",
54954 => "0111111101110000",
54955 => "0111111101110000",
54956 => "0111111101110000",
54957 => "0111111101110000",
54958 => "0111111101110000",
54959 => "0111111101110000",
54960 => "0111111101110000",
54961 => "0111111101110000",
54962 => "0111111101110000",
54963 => "0111111101110000",
54964 => "0111111101110000",
54965 => "0111111101110000",
54966 => "0111111101110000",
54967 => "0111111101110000",
54968 => "0111111101110000",
54969 => "0111111101110000",
54970 => "0111111101110000",
54971 => "0111111101110000",
54972 => "0111111101110000",
54973 => "0111111101110000",
54974 => "0111111101110000",
54975 => "0111111101110000",
54976 => "0111111101110000",
54977 => "0111111101110000",
54978 => "0111111101110000",
54979 => "0111111101110000",
54980 => "0111111101110000",
54981 => "0111111101110000",
54982 => "0111111101110000",
54983 => "0111111101110000",
54984 => "0111111101110000",
54985 => "0111111101110000",
54986 => "0111111101110000",
54987 => "0111111101110000",
54988 => "0111111101110000",
54989 => "0111111101110000",
54990 => "0111111101110000",
54991 => "0111111101110000",
54992 => "0111111101110000",
54993 => "0111111101110000",
54994 => "0111111101110000",
54995 => "0111111101110000",
54996 => "0111111101110000",
54997 => "0111111101110000",
54998 => "0111111101110000",
54999 => "0111111101110000",
55000 => "0111111101110000",
55001 => "0111111101110000",
55002 => "0111111101110000",
55003 => "0111111101110000",
55004 => "0111111101110000",
55005 => "0111111101110000",
55006 => "0111111101110000",
55007 => "0111111101110000",
55008 => "0111111101110000",
55009 => "0111111101110000",
55010 => "0111111101110000",
55011 => "0111111101110000",
55012 => "0111111101110000",
55013 => "0111111101110000",
55014 => "0111111101110000",
55015 => "0111111101110000",
55016 => "0111111101110000",
55017 => "0111111101110000",
55018 => "0111111101110000",
55019 => "0111111101110000",
55020 => "0111111101110000",
55021 => "0111111101110000",
55022 => "0111111101110000",
55023 => "0111111101110000",
55024 => "0111111101110000",
55025 => "0111111101110000",
55026 => "0111111101110000",
55027 => "0111111101110000",
55028 => "0111111101110000",
55029 => "0111111101110000",
55030 => "0111111101110000",
55031 => "0111111101110000",
55032 => "0111111101110000",
55033 => "0111111101110000",
55034 => "0111111101110000",
55035 => "0111111101110000",
55036 => "0111111101110000",
55037 => "0111111101110000",
55038 => "0111111101110000",
55039 => "0111111101110000",
55040 => "0111111101110000",
55041 => "0111111101110000",
55042 => "0111111101110000",
55043 => "0111111101110000",
55044 => "0111111101110000",
55045 => "0111111101110000",
55046 => "0111111101110000",
55047 => "0111111101110000",
55048 => "0111111101110000",
55049 => "0111111101110000",
55050 => "0111111101110000",
55051 => "0111111101110000",
55052 => "0111111101110000",
55053 => "0111111101110000",
55054 => "0111111101110000",
55055 => "0111111101110000",
55056 => "0111111101110000",
55057 => "0111111101110000",
55058 => "0111111101110000",
55059 => "0111111101110000",
55060 => "0111111101110000",
55061 => "0111111101110000",
55062 => "0111111101110000",
55063 => "0111111101110000",
55064 => "0111111101110000",
55065 => "0111111101110000",
55066 => "0111111101110000",
55067 => "0111111101110000",
55068 => "0111111101110000",
55069 => "0111111101110000",
55070 => "0111111101110000",
55071 => "0111111101110000",
55072 => "0111111101110000",
55073 => "0111111101110000",
55074 => "0111111101110000",
55075 => "0111111101110000",
55076 => "0111111101110000",
55077 => "0111111101110000",
55078 => "0111111101110000",
55079 => "0111111101110000",
55080 => "0111111101110000",
55081 => "0111111101110000",
55082 => "0111111101110000",
55083 => "0111111101110000",
55084 => "0111111101110000",
55085 => "0111111101110000",
55086 => "0111111101110000",
55087 => "0111111101110000",
55088 => "0111111101110000",
55089 => "0111111101110000",
55090 => "0111111101110000",
55091 => "0111111101110000",
55092 => "0111111101110000",
55093 => "0111111101110000",
55094 => "0111111101110000",
55095 => "0111111101110000",
55096 => "0111111101110000",
55097 => "0111111101110000",
55098 => "0111111101110000",
55099 => "0111111101110000",
55100 => "0111111101110000",
55101 => "0111111101110000",
55102 => "0111111101110000",
55103 => "0111111101110000",
55104 => "0111111101110000",
55105 => "0111111101110000",
55106 => "0111111101110000",
55107 => "0111111101110000",
55108 => "0111111101110000",
55109 => "0111111101110000",
55110 => "0111111101110000",
55111 => "0111111101110000",
55112 => "0111111101110000",
55113 => "0111111101110000",
55114 => "0111111101110000",
55115 => "0111111101110000",
55116 => "0111111101110000",
55117 => "0111111101110000",
55118 => "0111111101110000",
55119 => "0111111101110000",
55120 => "0111111101110000",
55121 => "0111111101110000",
55122 => "0111111101110000",
55123 => "0111111101110000",
55124 => "0111111101110000",
55125 => "0111111101110000",
55126 => "0111111101110000",
55127 => "0111111101110000",
55128 => "0111111101110000",
55129 => "0111111101110000",
55130 => "0111111101110000",
55131 => "0111111101110000",
55132 => "0111111101110000",
55133 => "0111111101110000",
55134 => "0111111101110000",
55135 => "0111111101110000",
55136 => "0111111101110000",
55137 => "0111111101110000",
55138 => "0111111101110000",
55139 => "0111111101110000",
55140 => "0111111101110000",
55141 => "0111111101110000",
55142 => "0111111101110000",
55143 => "0111111101110000",
55144 => "0111111101110000",
55145 => "0111111101110000",
55146 => "0111111101110000",
55147 => "0111111101110000",
55148 => "0111111101110000",
55149 => "0111111101110000",
55150 => "0111111101110000",
55151 => "0111111101110000",
55152 => "0111111101110000",
55153 => "0111111101110000",
55154 => "0111111101110000",
55155 => "0111111101110000",
55156 => "0111111101110000",
55157 => "0111111101110000",
55158 => "0111111101110000",
55159 => "0111111101110000",
55160 => "0111111101110000",
55161 => "0111111101110000",
55162 => "0111111101110000",
55163 => "0111111101110000",
55164 => "0111111101110000",
55165 => "0111111101110000",
55166 => "0111111101110000",
55167 => "0111111101110000",
55168 => "0111111101110000",
55169 => "0111111101110000",
55170 => "0111111101110000",
55171 => "0111111101110000",
55172 => "0111111101110000",
55173 => "0111111101110000",
55174 => "0111111101110000",
55175 => "0111111101110000",
55176 => "0111111101110000",
55177 => "0111111101110000",
55178 => "0111111101110000",
55179 => "0111111101110000",
55180 => "0111111101110000",
55181 => "0111111101110000",
55182 => "0111111101110000",
55183 => "0111111101110000",
55184 => "0111111101110000",
55185 => "0111111101110000",
55186 => "0111111101110000",
55187 => "0111111101110000",
55188 => "0111111101110000",
55189 => "0111111101110000",
55190 => "0111111101110000",
55191 => "0111111101110000",
55192 => "0111111101110000",
55193 => "0111111101110000",
55194 => "0111111101110000",
55195 => "0111111101110000",
55196 => "0111111101110000",
55197 => "0111111101110000",
55198 => "0111111101110000",
55199 => "0111111101110000",
55200 => "0111111101110000",
55201 => "0111111101110000",
55202 => "0111111101110000",
55203 => "0111111101110000",
55204 => "0111111101110000",
55205 => "0111111101110000",
55206 => "0111111101110000",
55207 => "0111111101110000",
55208 => "0111111101110000",
55209 => "0111111101110000",
55210 => "0111111101110000",
55211 => "0111111101110000",
55212 => "0111111101110000",
55213 => "0111111101110000",
55214 => "0111111101110000",
55215 => "0111111110000000",
55216 => "0111111110000000",
55217 => "0111111110000000",
55218 => "0111111110000000",
55219 => "0111111110000000",
55220 => "0111111110000000",
55221 => "0111111110000000",
55222 => "0111111110000000",
55223 => "0111111110000000",
55224 => "0111111110000000",
55225 => "0111111110000000",
55226 => "0111111110000000",
55227 => "0111111110000000",
55228 => "0111111110000000",
55229 => "0111111110000000",
55230 => "0111111110000000",
55231 => "0111111110000000",
55232 => "0111111110000000",
55233 => "0111111110000000",
55234 => "0111111110000000",
55235 => "0111111110000000",
55236 => "0111111110000000",
55237 => "0111111110000000",
55238 => "0111111110000000",
55239 => "0111111110000000",
55240 => "0111111110000000",
55241 => "0111111110000000",
55242 => "0111111110000000",
55243 => "0111111110000000",
55244 => "0111111110000000",
55245 => "0111111110000000",
55246 => "0111111110000000",
55247 => "0111111110000000",
55248 => "0111111110000000",
55249 => "0111111110000000",
55250 => "0111111110000000",
55251 => "0111111110000000",
55252 => "0111111110000000",
55253 => "0111111110000000",
55254 => "0111111110000000",
55255 => "0111111110000000",
55256 => "0111111110000000",
55257 => "0111111110000000",
55258 => "0111111110000000",
55259 => "0111111110000000",
55260 => "0111111110000000",
55261 => "0111111110000000",
55262 => "0111111110000000",
55263 => "0111111110000000",
55264 => "0111111110000000",
55265 => "0111111110000000",
55266 => "0111111110000000",
55267 => "0111111110000000",
55268 => "0111111110000000",
55269 => "0111111110000000",
55270 => "0111111110000000",
55271 => "0111111110000000",
55272 => "0111111110000000",
55273 => "0111111110000000",
55274 => "0111111110000000",
55275 => "0111111110000000",
55276 => "0111111110000000",
55277 => "0111111110000000",
55278 => "0111111110000000",
55279 => "0111111110000000",
55280 => "0111111110000000",
55281 => "0111111110000000",
55282 => "0111111110000000",
55283 => "0111111110000000",
55284 => "0111111110000000",
55285 => "0111111110000000",
55286 => "0111111110000000",
55287 => "0111111110000000",
55288 => "0111111110000000",
55289 => "0111111110000000",
55290 => "0111111110000000",
55291 => "0111111110000000",
55292 => "0111111110000000",
55293 => "0111111110000000",
55294 => "0111111110000000",
55295 => "0111111110000000",
55296 => "0111111110000000",
55297 => "0111111110000000",
55298 => "0111111110000000",
55299 => "0111111110000000",
55300 => "0111111110000000",
55301 => "0111111110000000",
55302 => "0111111110000000",
55303 => "0111111110000000",
55304 => "0111111110000000",
55305 => "0111111110000000",
55306 => "0111111110000000",
55307 => "0111111110000000",
55308 => "0111111110000000",
55309 => "0111111110000000",
55310 => "0111111110000000",
55311 => "0111111110000000",
55312 => "0111111110000000",
55313 => "0111111110000000",
55314 => "0111111110000000",
55315 => "0111111110000000",
55316 => "0111111110000000",
55317 => "0111111110000000",
55318 => "0111111110000000",
55319 => "0111111110000000",
55320 => "0111111110000000",
55321 => "0111111110000000",
55322 => "0111111110000000",
55323 => "0111111110000000",
55324 => "0111111110000000",
55325 => "0111111110000000",
55326 => "0111111110000000",
55327 => "0111111110000000",
55328 => "0111111110000000",
55329 => "0111111110000000",
55330 => "0111111110000000",
55331 => "0111111110000000",
55332 => "0111111110000000",
55333 => "0111111110000000",
55334 => "0111111110000000",
55335 => "0111111110000000",
55336 => "0111111110000000",
55337 => "0111111110000000",
55338 => "0111111110000000",
55339 => "0111111110000000",
55340 => "0111111110000000",
55341 => "0111111110000000",
55342 => "0111111110000000",
55343 => "0111111110000000",
55344 => "0111111110000000",
55345 => "0111111110000000",
55346 => "0111111110000000",
55347 => "0111111110000000",
55348 => "0111111110000000",
55349 => "0111111110000000",
55350 => "0111111110000000",
55351 => "0111111110000000",
55352 => "0111111110000000",
55353 => "0111111110000000",
55354 => "0111111110000000",
55355 => "0111111110000000",
55356 => "0111111110000000",
55357 => "0111111110000000",
55358 => "0111111110000000",
55359 => "0111111110000000",
55360 => "0111111110000000",
55361 => "0111111110000000",
55362 => "0111111110000000",
55363 => "0111111110000000",
55364 => "0111111110000000",
55365 => "0111111110000000",
55366 => "0111111110000000",
55367 => "0111111110000000",
55368 => "0111111110000000",
55369 => "0111111110000000",
55370 => "0111111110000000",
55371 => "0111111110000000",
55372 => "0111111110000000",
55373 => "0111111110000000",
55374 => "0111111110000000",
55375 => "0111111110000000",
55376 => "0111111110000000",
55377 => "0111111110000000",
55378 => "0111111110000000",
55379 => "0111111110000000",
55380 => "0111111110000000",
55381 => "0111111110000000",
55382 => "0111111110000000",
55383 => "0111111110000000",
55384 => "0111111110000000",
55385 => "0111111110000000",
55386 => "0111111110000000",
55387 => "0111111110000000",
55388 => "0111111110000000",
55389 => "0111111110000000",
55390 => "0111111110000000",
55391 => "0111111110000000",
55392 => "0111111110000000",
55393 => "0111111110000000",
55394 => "0111111110000000",
55395 => "0111111110000000",
55396 => "0111111110000000",
55397 => "0111111110000000",
55398 => "0111111110000000",
55399 => "0111111110000000",
55400 => "0111111110000000",
55401 => "0111111110000000",
55402 => "0111111110000000",
55403 => "0111111110000000",
55404 => "0111111110000000",
55405 => "0111111110000000",
55406 => "0111111110000000",
55407 => "0111111110000000",
55408 => "0111111110000000",
55409 => "0111111110000000",
55410 => "0111111110000000",
55411 => "0111111110000000",
55412 => "0111111110000000",
55413 => "0111111110000000",
55414 => "0111111110000000",
55415 => "0111111110000000",
55416 => "0111111110000000",
55417 => "0111111110000000",
55418 => "0111111110000000",
55419 => "0111111110000000",
55420 => "0111111110000000",
55421 => "0111111110000000",
55422 => "0111111110000000",
55423 => "0111111110000000",
55424 => "0111111110000000",
55425 => "0111111110000000",
55426 => "0111111110000000",
55427 => "0111111110000000",
55428 => "0111111110000000",
55429 => "0111111110000000",
55430 => "0111111110000000",
55431 => "0111111110000000",
55432 => "0111111110000000",
55433 => "0111111110000000",
55434 => "0111111110000000",
55435 => "0111111110000000",
55436 => "0111111110000000",
55437 => "0111111110000000",
55438 => "0111111110000000",
55439 => "0111111110000000",
55440 => "0111111110000000",
55441 => "0111111110000000",
55442 => "0111111110000000",
55443 => "0111111110000000",
55444 => "0111111110000000",
55445 => "0111111110000000",
55446 => "0111111110000000",
55447 => "0111111110000000",
55448 => "0111111110000000",
55449 => "0111111110000000",
55450 => "0111111110000000",
55451 => "0111111110000000",
55452 => "0111111110000000",
55453 => "0111111110000000",
55454 => "0111111110000000",
55455 => "0111111110000000",
55456 => "0111111110000000",
55457 => "0111111110000000",
55458 => "0111111110000000",
55459 => "0111111110000000",
55460 => "0111111110000000",
55461 => "0111111110000000",
55462 => "0111111110000000",
55463 => "0111111110000000",
55464 => "0111111110000000",
55465 => "0111111110000000",
55466 => "0111111110000000",
55467 => "0111111110000000",
55468 => "0111111110000000",
55469 => "0111111110000000",
55470 => "0111111110000000",
55471 => "0111111110000000",
55472 => "0111111110000000",
55473 => "0111111110000000",
55474 => "0111111110000000",
55475 => "0111111110000000",
55476 => "0111111110000000",
55477 => "0111111110000000",
55478 => "0111111110000000",
55479 => "0111111110000000",
55480 => "0111111110000000",
55481 => "0111111110000000",
55482 => "0111111110000000",
55483 => "0111111110000000",
55484 => "0111111110000000",
55485 => "0111111110000000",
55486 => "0111111110000000",
55487 => "0111111110000000",
55488 => "0111111110000000",
55489 => "0111111110000000",
55490 => "0111111110000000",
55491 => "0111111110000000",
55492 => "0111111110000000",
55493 => "0111111110000000",
55494 => "0111111110000000",
55495 => "0111111110000000",
55496 => "0111111110000000",
55497 => "0111111110000000",
55498 => "0111111110000000",
55499 => "0111111110000000",
55500 => "0111111110000000",
55501 => "0111111110000000",
55502 => "0111111110000000",
55503 => "0111111110000000",
55504 => "0111111110000000",
55505 => "0111111110000000",
55506 => "0111111110000000",
55507 => "0111111110000000",
55508 => "0111111110000000",
55509 => "0111111110000000",
55510 => "0111111110000000",
55511 => "0111111110000000",
55512 => "0111111110000000",
55513 => "0111111110000000",
55514 => "0111111110000000",
55515 => "0111111110000000",
55516 => "0111111110000000",
55517 => "0111111110000000",
55518 => "0111111110000000",
55519 => "0111111110000000",
55520 => "0111111110000000",
55521 => "0111111110000000",
55522 => "0111111110000000",
55523 => "0111111110000000",
55524 => "0111111110000000",
55525 => "0111111110000000",
55526 => "0111111110000000",
55527 => "0111111110000000",
55528 => "0111111110000000",
55529 => "0111111110000000",
55530 => "0111111110000000",
55531 => "0111111110000000",
55532 => "0111111110000000",
55533 => "0111111110000000",
55534 => "0111111110000000",
55535 => "0111111110000000",
55536 => "0111111110000000",
55537 => "0111111110000000",
55538 => "0111111110000000",
55539 => "0111111110000000",
55540 => "0111111110000000",
55541 => "0111111110000000",
55542 => "0111111110000000",
55543 => "0111111110000000",
55544 => "0111111110000000",
55545 => "0111111110000000",
55546 => "0111111110000000",
55547 => "0111111110000000",
55548 => "0111111110000000",
55549 => "0111111110000000",
55550 => "0111111110000000",
55551 => "0111111110000000",
55552 => "0111111110000000",
55553 => "0111111110000000",
55554 => "0111111110000000",
55555 => "0111111110000000",
55556 => "0111111110000000",
55557 => "0111111110000000",
55558 => "0111111110000000",
55559 => "0111111110000000",
55560 => "0111111110000000",
55561 => "0111111110000000",
55562 => "0111111110000000",
55563 => "0111111110000000",
55564 => "0111111110000000",
55565 => "0111111110000000",
55566 => "0111111110000000",
55567 => "0111111110000000",
55568 => "0111111110000000",
55569 => "0111111110000000",
55570 => "0111111110000000",
55571 => "0111111110000000",
55572 => "0111111110000000",
55573 => "0111111110000000",
55574 => "0111111110000000",
55575 => "0111111110000000",
55576 => "0111111110000000",
55577 => "0111111110000000",
55578 => "0111111110000000",
55579 => "0111111110000000",
55580 => "0111111110000000",
55581 => "0111111110000000",
55582 => "0111111110000000",
55583 => "0111111110000000",
55584 => "0111111110000000",
55585 => "0111111110000000",
55586 => "0111111110000000",
55587 => "0111111110000000",
55588 => "0111111110000000",
55589 => "0111111110000000",
55590 => "0111111110000000",
55591 => "0111111110000000",
55592 => "0111111110000000",
55593 => "0111111110000000",
55594 => "0111111110000000",
55595 => "0111111110000000",
55596 => "0111111110000000",
55597 => "0111111110000000",
55598 => "0111111110000000",
55599 => "0111111110000000",
55600 => "0111111110000000",
55601 => "0111111110000000",
55602 => "0111111110000000",
55603 => "0111111110000000",
55604 => "0111111110000000",
55605 => "0111111110000000",
55606 => "0111111110000000",
55607 => "0111111110000000",
55608 => "0111111110000000",
55609 => "0111111110000000",
55610 => "0111111110000000",
55611 => "0111111110000000",
55612 => "0111111110000000",
55613 => "0111111110000000",
55614 => "0111111110000000",
55615 => "0111111110000000",
55616 => "0111111110000000",
55617 => "0111111110000000",
55618 => "0111111110000000",
55619 => "0111111110000000",
55620 => "0111111110000000",
55621 => "0111111110000000",
55622 => "0111111110000000",
55623 => "0111111110000000",
55624 => "0111111110000000",
55625 => "0111111110000000",
55626 => "0111111110000000",
55627 => "0111111110000000",
55628 => "0111111110000000",
55629 => "0111111110000000",
55630 => "0111111110000000",
55631 => "0111111110000000",
55632 => "0111111110000000",
55633 => "0111111110000000",
55634 => "0111111110000000",
55635 => "0111111110000000",
55636 => "0111111110000000",
55637 => "0111111110000000",
55638 => "0111111110000000",
55639 => "0111111110000000",
55640 => "0111111110000000",
55641 => "0111111110000000",
55642 => "0111111110000000",
55643 => "0111111110000000",
55644 => "0111111110000000",
55645 => "0111111110000000",
55646 => "0111111110000000",
55647 => "0111111110000000",
55648 => "0111111110000000",
55649 => "0111111110000000",
55650 => "0111111110000000",
55651 => "0111111110000000",
55652 => "0111111110000000",
55653 => "0111111110000000",
55654 => "0111111110000000",
55655 => "0111111110000000",
55656 => "0111111110000000",
55657 => "0111111110000000",
55658 => "0111111110000000",
55659 => "0111111110000000",
55660 => "0111111110000000",
55661 => "0111111110000000",
55662 => "0111111110000000",
55663 => "0111111110000000",
55664 => "0111111110000000",
55665 => "0111111110000000",
55666 => "0111111110000000",
55667 => "0111111110000000",
55668 => "0111111110000000",
55669 => "0111111110000000",
55670 => "0111111110000000",
55671 => "0111111110000000",
55672 => "0111111110000000",
55673 => "0111111110000000",
55674 => "0111111110000000",
55675 => "0111111110000000",
55676 => "0111111110000000",
55677 => "0111111110000000",
55678 => "0111111110000000",
55679 => "0111111110000000",
55680 => "0111111110000000",
55681 => "0111111110000000",
55682 => "0111111110000000",
55683 => "0111111110000000",
55684 => "0111111110000000",
55685 => "0111111110000000",
55686 => "0111111110000000",
55687 => "0111111110000000",
55688 => "0111111110000000",
55689 => "0111111110000000",
55690 => "0111111110000000",
55691 => "0111111110000000",
55692 => "0111111110000000",
55693 => "0111111110000000",
55694 => "0111111110000000",
55695 => "0111111110000000",
55696 => "0111111110000000",
55697 => "0111111110000000",
55698 => "0111111110000000",
55699 => "0111111110000000",
55700 => "0111111110000000",
55701 => "0111111110000000",
55702 => "0111111110000000",
55703 => "0111111110000000",
55704 => "0111111110000000",
55705 => "0111111110000000",
55706 => "0111111110000000",
55707 => "0111111110000000",
55708 => "0111111110000000",
55709 => "0111111110000000",
55710 => "0111111110000000",
55711 => "0111111110000000",
55712 => "0111111110000000",
55713 => "0111111110000000",
55714 => "0111111110000000",
55715 => "0111111110000000",
55716 => "0111111110000000",
55717 => "0111111110000000",
55718 => "0111111110000000",
55719 => "0111111110000000",
55720 => "0111111110000000",
55721 => "0111111110000000",
55722 => "0111111110000000",
55723 => "0111111110000000",
55724 => "0111111110000000",
55725 => "0111111110000000",
55726 => "0111111110000000",
55727 => "0111111110000000",
55728 => "0111111110000000",
55729 => "0111111110000000",
55730 => "0111111110010000",
55731 => "0111111110010000",
55732 => "0111111110010000",
55733 => "0111111110010000",
55734 => "0111111110010000",
55735 => "0111111110010000",
55736 => "0111111110010000",
55737 => "0111111110010000",
55738 => "0111111110010000",
55739 => "0111111110010000",
55740 => "0111111110010000",
55741 => "0111111110010000",
55742 => "0111111110010000",
55743 => "0111111110010000",
55744 => "0111111110010000",
55745 => "0111111110010000",
55746 => "0111111110010000",
55747 => "0111111110010000",
55748 => "0111111110010000",
55749 => "0111111110010000",
55750 => "0111111110010000",
55751 => "0111111110010000",
55752 => "0111111110010000",
55753 => "0111111110010000",
55754 => "0111111110010000",
55755 => "0111111110010000",
55756 => "0111111110010000",
55757 => "0111111110010000",
55758 => "0111111110010000",
55759 => "0111111110010000",
55760 => "0111111110010000",
55761 => "0111111110010000",
55762 => "0111111110010000",
55763 => "0111111110010000",
55764 => "0111111110010000",
55765 => "0111111110010000",
55766 => "0111111110010000",
55767 => "0111111110010000",
55768 => "0111111110010000",
55769 => "0111111110010000",
55770 => "0111111110010000",
55771 => "0111111110010000",
55772 => "0111111110010000",
55773 => "0111111110010000",
55774 => "0111111110010000",
55775 => "0111111110010000",
55776 => "0111111110010000",
55777 => "0111111110010000",
55778 => "0111111110010000",
55779 => "0111111110010000",
55780 => "0111111110010000",
55781 => "0111111110010000",
55782 => "0111111110010000",
55783 => "0111111110010000",
55784 => "0111111110010000",
55785 => "0111111110010000",
55786 => "0111111110010000",
55787 => "0111111110010000",
55788 => "0111111110010000",
55789 => "0111111110010000",
55790 => "0111111110010000",
55791 => "0111111110010000",
55792 => "0111111110010000",
55793 => "0111111110010000",
55794 => "0111111110010000",
55795 => "0111111110010000",
55796 => "0111111110010000",
55797 => "0111111110010000",
55798 => "0111111110010000",
55799 => "0111111110010000",
55800 => "0111111110010000",
55801 => "0111111110010000",
55802 => "0111111110010000",
55803 => "0111111110010000",
55804 => "0111111110010000",
55805 => "0111111110010000",
55806 => "0111111110010000",
55807 => "0111111110010000",
55808 => "0111111110010000",
55809 => "0111111110010000",
55810 => "0111111110010000",
55811 => "0111111110010000",
55812 => "0111111110010000",
55813 => "0111111110010000",
55814 => "0111111110010000",
55815 => "0111111110010000",
55816 => "0111111110010000",
55817 => "0111111110010000",
55818 => "0111111110010000",
55819 => "0111111110010000",
55820 => "0111111110010000",
55821 => "0111111110010000",
55822 => "0111111110010000",
55823 => "0111111110010000",
55824 => "0111111110010000",
55825 => "0111111110010000",
55826 => "0111111110010000",
55827 => "0111111110010000",
55828 => "0111111110010000",
55829 => "0111111110010000",
55830 => "0111111110010000",
55831 => "0111111110010000",
55832 => "0111111110010000",
55833 => "0111111110010000",
55834 => "0111111110010000",
55835 => "0111111110010000",
55836 => "0111111110010000",
55837 => "0111111110010000",
55838 => "0111111110010000",
55839 => "0111111110010000",
55840 => "0111111110010000",
55841 => "0111111110010000",
55842 => "0111111110010000",
55843 => "0111111110010000",
55844 => "0111111110010000",
55845 => "0111111110010000",
55846 => "0111111110010000",
55847 => "0111111110010000",
55848 => "0111111110010000",
55849 => "0111111110010000",
55850 => "0111111110010000",
55851 => "0111111110010000",
55852 => "0111111110010000",
55853 => "0111111110010000",
55854 => "0111111110010000",
55855 => "0111111110010000",
55856 => "0111111110010000",
55857 => "0111111110010000",
55858 => "0111111110010000",
55859 => "0111111110010000",
55860 => "0111111110010000",
55861 => "0111111110010000",
55862 => "0111111110010000",
55863 => "0111111110010000",
55864 => "0111111110010000",
55865 => "0111111110010000",
55866 => "0111111110010000",
55867 => "0111111110010000",
55868 => "0111111110010000",
55869 => "0111111110010000",
55870 => "0111111110010000",
55871 => "0111111110010000",
55872 => "0111111110010000",
55873 => "0111111110010000",
55874 => "0111111110010000",
55875 => "0111111110010000",
55876 => "0111111110010000",
55877 => "0111111110010000",
55878 => "0111111110010000",
55879 => "0111111110010000",
55880 => "0111111110010000",
55881 => "0111111110010000",
55882 => "0111111110010000",
55883 => "0111111110010000",
55884 => "0111111110010000",
55885 => "0111111110010000",
55886 => "0111111110010000",
55887 => "0111111110010000",
55888 => "0111111110010000",
55889 => "0111111110010000",
55890 => "0111111110010000",
55891 => "0111111110010000",
55892 => "0111111110010000",
55893 => "0111111110010000",
55894 => "0111111110010000",
55895 => "0111111110010000",
55896 => "0111111110010000",
55897 => "0111111110010000",
55898 => "0111111110010000",
55899 => "0111111110010000",
55900 => "0111111110010000",
55901 => "0111111110010000",
55902 => "0111111110010000",
55903 => "0111111110010000",
55904 => "0111111110010000",
55905 => "0111111110010000",
55906 => "0111111110010000",
55907 => "0111111110010000",
55908 => "0111111110010000",
55909 => "0111111110010000",
55910 => "0111111110010000",
55911 => "0111111110010000",
55912 => "0111111110010000",
55913 => "0111111110010000",
55914 => "0111111110010000",
55915 => "0111111110010000",
55916 => "0111111110010000",
55917 => "0111111110010000",
55918 => "0111111110010000",
55919 => "0111111110010000",
55920 => "0111111110010000",
55921 => "0111111110010000",
55922 => "0111111110010000",
55923 => "0111111110010000",
55924 => "0111111110010000",
55925 => "0111111110010000",
55926 => "0111111110010000",
55927 => "0111111110010000",
55928 => "0111111110010000",
55929 => "0111111110010000",
55930 => "0111111110010000",
55931 => "0111111110010000",
55932 => "0111111110010000",
55933 => "0111111110010000",
55934 => "0111111110010000",
55935 => "0111111110010000",
55936 => "0111111110010000",
55937 => "0111111110010000",
55938 => "0111111110010000",
55939 => "0111111110010000",
55940 => "0111111110010000",
55941 => "0111111110010000",
55942 => "0111111110010000",
55943 => "0111111110010000",
55944 => "0111111110010000",
55945 => "0111111110010000",
55946 => "0111111110010000",
55947 => "0111111110010000",
55948 => "0111111110010000",
55949 => "0111111110010000",
55950 => "0111111110010000",
55951 => "0111111110010000",
55952 => "0111111110010000",
55953 => "0111111110010000",
55954 => "0111111110010000",
55955 => "0111111110010000",
55956 => "0111111110010000",
55957 => "0111111110010000",
55958 => "0111111110010000",
55959 => "0111111110010000",
55960 => "0111111110010000",
55961 => "0111111110010000",
55962 => "0111111110010000",
55963 => "0111111110010000",
55964 => "0111111110010000",
55965 => "0111111110010000",
55966 => "0111111110010000",
55967 => "0111111110010000",
55968 => "0111111110010000",
55969 => "0111111110010000",
55970 => "0111111110010000",
55971 => "0111111110010000",
55972 => "0111111110010000",
55973 => "0111111110010000",
55974 => "0111111110010000",
55975 => "0111111110010000",
55976 => "0111111110010000",
55977 => "0111111110010000",
55978 => "0111111110010000",
55979 => "0111111110010000",
55980 => "0111111110010000",
55981 => "0111111110010000",
55982 => "0111111110010000",
55983 => "0111111110010000",
55984 => "0111111110010000",
55985 => "0111111110010000",
55986 => "0111111110010000",
55987 => "0111111110010000",
55988 => "0111111110010000",
55989 => "0111111110010000",
55990 => "0111111110010000",
55991 => "0111111110010000",
55992 => "0111111110010000",
55993 => "0111111110010000",
55994 => "0111111110010000",
55995 => "0111111110010000",
55996 => "0111111110010000",
55997 => "0111111110010000",
55998 => "0111111110010000",
55999 => "0111111110010000",
56000 => "0111111110010000",
56001 => "0111111110010000",
56002 => "0111111110010000",
56003 => "0111111110010000",
56004 => "0111111110010000",
56005 => "0111111110010000",
56006 => "0111111110010000",
56007 => "0111111110010000",
56008 => "0111111110010000",
56009 => "0111111110010000",
56010 => "0111111110010000",
56011 => "0111111110010000",
56012 => "0111111110010000",
56013 => "0111111110010000",
56014 => "0111111110010000",
56015 => "0111111110010000",
56016 => "0111111110010000",
56017 => "0111111110010000",
56018 => "0111111110010000",
56019 => "0111111110010000",
56020 => "0111111110010000",
56021 => "0111111110010000",
56022 => "0111111110010000",
56023 => "0111111110010000",
56024 => "0111111110010000",
56025 => "0111111110010000",
56026 => "0111111110010000",
56027 => "0111111110010000",
56028 => "0111111110010000",
56029 => "0111111110010000",
56030 => "0111111110010000",
56031 => "0111111110010000",
56032 => "0111111110010000",
56033 => "0111111110010000",
56034 => "0111111110010000",
56035 => "0111111110010000",
56036 => "0111111110010000",
56037 => "0111111110010000",
56038 => "0111111110010000",
56039 => "0111111110010000",
56040 => "0111111110010000",
56041 => "0111111110010000",
56042 => "0111111110010000",
56043 => "0111111110010000",
56044 => "0111111110010000",
56045 => "0111111110010000",
56046 => "0111111110010000",
56047 => "0111111110010000",
56048 => "0111111110010000",
56049 => "0111111110010000",
56050 => "0111111110010000",
56051 => "0111111110010000",
56052 => "0111111110010000",
56053 => "0111111110010000",
56054 => "0111111110010000",
56055 => "0111111110010000",
56056 => "0111111110010000",
56057 => "0111111110010000",
56058 => "0111111110010000",
56059 => "0111111110010000",
56060 => "0111111110010000",
56061 => "0111111110010000",
56062 => "0111111110010000",
56063 => "0111111110010000",
56064 => "0111111110010000",
56065 => "0111111110010000",
56066 => "0111111110010000",
56067 => "0111111110010000",
56068 => "0111111110010000",
56069 => "0111111110010000",
56070 => "0111111110010000",
56071 => "0111111110010000",
56072 => "0111111110010000",
56073 => "0111111110010000",
56074 => "0111111110010000",
56075 => "0111111110010000",
56076 => "0111111110010000",
56077 => "0111111110010000",
56078 => "0111111110010000",
56079 => "0111111110010000",
56080 => "0111111110010000",
56081 => "0111111110010000",
56082 => "0111111110010000",
56083 => "0111111110010000",
56084 => "0111111110010000",
56085 => "0111111110010000",
56086 => "0111111110010000",
56087 => "0111111110010000",
56088 => "0111111110010000",
56089 => "0111111110010000",
56090 => "0111111110010000",
56091 => "0111111110010000",
56092 => "0111111110010000",
56093 => "0111111110010000",
56094 => "0111111110010000",
56095 => "0111111110010000",
56096 => "0111111110010000",
56097 => "0111111110010000",
56098 => "0111111110010000",
56099 => "0111111110010000",
56100 => "0111111110010000",
56101 => "0111111110010000",
56102 => "0111111110010000",
56103 => "0111111110010000",
56104 => "0111111110010000",
56105 => "0111111110010000",
56106 => "0111111110010000",
56107 => "0111111110010000",
56108 => "0111111110010000",
56109 => "0111111110010000",
56110 => "0111111110010000",
56111 => "0111111110010000",
56112 => "0111111110010000",
56113 => "0111111110010000",
56114 => "0111111110010000",
56115 => "0111111110010000",
56116 => "0111111110010000",
56117 => "0111111110010000",
56118 => "0111111110010000",
56119 => "0111111110010000",
56120 => "0111111110010000",
56121 => "0111111110010000",
56122 => "0111111110010000",
56123 => "0111111110010000",
56124 => "0111111110010000",
56125 => "0111111110010000",
56126 => "0111111110010000",
56127 => "0111111110010000",
56128 => "0111111110010000",
56129 => "0111111110010000",
56130 => "0111111110010000",
56131 => "0111111110010000",
56132 => "0111111110010000",
56133 => "0111111110010000",
56134 => "0111111110010000",
56135 => "0111111110010000",
56136 => "0111111110010000",
56137 => "0111111110010000",
56138 => "0111111110010000",
56139 => "0111111110010000",
56140 => "0111111110010000",
56141 => "0111111110010000",
56142 => "0111111110010000",
56143 => "0111111110010000",
56144 => "0111111110010000",
56145 => "0111111110010000",
56146 => "0111111110010000",
56147 => "0111111110010000",
56148 => "0111111110010000",
56149 => "0111111110010000",
56150 => "0111111110010000",
56151 => "0111111110010000",
56152 => "0111111110010000",
56153 => "0111111110010000",
56154 => "0111111110010000",
56155 => "0111111110010000",
56156 => "0111111110010000",
56157 => "0111111110010000",
56158 => "0111111110010000",
56159 => "0111111110010000",
56160 => "0111111110010000",
56161 => "0111111110010000",
56162 => "0111111110010000",
56163 => "0111111110010000",
56164 => "0111111110010000",
56165 => "0111111110010000",
56166 => "0111111110010000",
56167 => "0111111110010000",
56168 => "0111111110010000",
56169 => "0111111110010000",
56170 => "0111111110010000",
56171 => "0111111110010000",
56172 => "0111111110010000",
56173 => "0111111110010000",
56174 => "0111111110010000",
56175 => "0111111110010000",
56176 => "0111111110010000",
56177 => "0111111110010000",
56178 => "0111111110010000",
56179 => "0111111110010000",
56180 => "0111111110010000",
56181 => "0111111110010000",
56182 => "0111111110010000",
56183 => "0111111110010000",
56184 => "0111111110010000",
56185 => "0111111110010000",
56186 => "0111111110010000",
56187 => "0111111110010000",
56188 => "0111111110010000",
56189 => "0111111110010000",
56190 => "0111111110010000",
56191 => "0111111110010000",
56192 => "0111111110010000",
56193 => "0111111110010000",
56194 => "0111111110010000",
56195 => "0111111110010000",
56196 => "0111111110010000",
56197 => "0111111110010000",
56198 => "0111111110010000",
56199 => "0111111110010000",
56200 => "0111111110010000",
56201 => "0111111110010000",
56202 => "0111111110010000",
56203 => "0111111110010000",
56204 => "0111111110010000",
56205 => "0111111110010000",
56206 => "0111111110010000",
56207 => "0111111110010000",
56208 => "0111111110010000",
56209 => "0111111110010000",
56210 => "0111111110010000",
56211 => "0111111110010000",
56212 => "0111111110010000",
56213 => "0111111110010000",
56214 => "0111111110010000",
56215 => "0111111110010000",
56216 => "0111111110010000",
56217 => "0111111110010000",
56218 => "0111111110010000",
56219 => "0111111110010000",
56220 => "0111111110010000",
56221 => "0111111110010000",
56222 => "0111111110010000",
56223 => "0111111110010000",
56224 => "0111111110010000",
56225 => "0111111110010000",
56226 => "0111111110010000",
56227 => "0111111110010000",
56228 => "0111111110010000",
56229 => "0111111110010000",
56230 => "0111111110010000",
56231 => "0111111110010000",
56232 => "0111111110010000",
56233 => "0111111110010000",
56234 => "0111111110010000",
56235 => "0111111110010000",
56236 => "0111111110010000",
56237 => "0111111110010000",
56238 => "0111111110010000",
56239 => "0111111110010000",
56240 => "0111111110010000",
56241 => "0111111110010000",
56242 => "0111111110010000",
56243 => "0111111110010000",
56244 => "0111111110010000",
56245 => "0111111110010000",
56246 => "0111111110010000",
56247 => "0111111110010000",
56248 => "0111111110010000",
56249 => "0111111110010000",
56250 => "0111111110010000",
56251 => "0111111110010000",
56252 => "0111111110010000",
56253 => "0111111110010000",
56254 => "0111111110010000",
56255 => "0111111110010000",
56256 => "0111111110010000",
56257 => "0111111110010000",
56258 => "0111111110010000",
56259 => "0111111110010000",
56260 => "0111111110010000",
56261 => "0111111110010000",
56262 => "0111111110010000",
56263 => "0111111110010000",
56264 => "0111111110010000",
56265 => "0111111110010000",
56266 => "0111111110010000",
56267 => "0111111110010000",
56268 => "0111111110010000",
56269 => "0111111110010000",
56270 => "0111111110010000",
56271 => "0111111110010000",
56272 => "0111111110010000",
56273 => "0111111110010000",
56274 => "0111111110010000",
56275 => "0111111110010000",
56276 => "0111111110010000",
56277 => "0111111110010000",
56278 => "0111111110010000",
56279 => "0111111110010000",
56280 => "0111111110010000",
56281 => "0111111110010000",
56282 => "0111111110010000",
56283 => "0111111110010000",
56284 => "0111111110010000",
56285 => "0111111110010000",
56286 => "0111111110010000",
56287 => "0111111110010000",
56288 => "0111111110010000",
56289 => "0111111110010000",
56290 => "0111111110010000",
56291 => "0111111110010000",
56292 => "0111111110010000",
56293 => "0111111110010000",
56294 => "0111111110010000",
56295 => "0111111110010000",
56296 => "0111111110010000",
56297 => "0111111110010000",
56298 => "0111111110010000",
56299 => "0111111110010000",
56300 => "0111111110010000",
56301 => "0111111110010000",
56302 => "0111111110010000",
56303 => "0111111110010000",
56304 => "0111111110010000",
56305 => "0111111110010000",
56306 => "0111111110010000",
56307 => "0111111110010000",
56308 => "0111111110010000",
56309 => "0111111110010000",
56310 => "0111111110010000",
56311 => "0111111110010000",
56312 => "0111111110010000",
56313 => "0111111110010000",
56314 => "0111111110010000",
56315 => "0111111110010000",
56316 => "0111111110010000",
56317 => "0111111110010000",
56318 => "0111111110100000",
56319 => "0111111110100000",
56320 => "0111111110100000",
56321 => "0111111110100000",
56322 => "0111111110100000",
56323 => "0111111110100000",
56324 => "0111111110100000",
56325 => "0111111110100000",
56326 => "0111111110100000",
56327 => "0111111110100000",
56328 => "0111111110100000",
56329 => "0111111110100000",
56330 => "0111111110100000",
56331 => "0111111110100000",
56332 => "0111111110100000",
56333 => "0111111110100000",
56334 => "0111111110100000",
56335 => "0111111110100000",
56336 => "0111111110100000",
56337 => "0111111110100000",
56338 => "0111111110100000",
56339 => "0111111110100000",
56340 => "0111111110100000",
56341 => "0111111110100000",
56342 => "0111111110100000",
56343 => "0111111110100000",
56344 => "0111111110100000",
56345 => "0111111110100000",
56346 => "0111111110100000",
56347 => "0111111110100000",
56348 => "0111111110100000",
56349 => "0111111110100000",
56350 => "0111111110100000",
56351 => "0111111110100000",
56352 => "0111111110100000",
56353 => "0111111110100000",
56354 => "0111111110100000",
56355 => "0111111110100000",
56356 => "0111111110100000",
56357 => "0111111110100000",
56358 => "0111111110100000",
56359 => "0111111110100000",
56360 => "0111111110100000",
56361 => "0111111110100000",
56362 => "0111111110100000",
56363 => "0111111110100000",
56364 => "0111111110100000",
56365 => "0111111110100000",
56366 => "0111111110100000",
56367 => "0111111110100000",
56368 => "0111111110100000",
56369 => "0111111110100000",
56370 => "0111111110100000",
56371 => "0111111110100000",
56372 => "0111111110100000",
56373 => "0111111110100000",
56374 => "0111111110100000",
56375 => "0111111110100000",
56376 => "0111111110100000",
56377 => "0111111110100000",
56378 => "0111111110100000",
56379 => "0111111110100000",
56380 => "0111111110100000",
56381 => "0111111110100000",
56382 => "0111111110100000",
56383 => "0111111110100000",
56384 => "0111111110100000",
56385 => "0111111110100000",
56386 => "0111111110100000",
56387 => "0111111110100000",
56388 => "0111111110100000",
56389 => "0111111110100000",
56390 => "0111111110100000",
56391 => "0111111110100000",
56392 => "0111111110100000",
56393 => "0111111110100000",
56394 => "0111111110100000",
56395 => "0111111110100000",
56396 => "0111111110100000",
56397 => "0111111110100000",
56398 => "0111111110100000",
56399 => "0111111110100000",
56400 => "0111111110100000",
56401 => "0111111110100000",
56402 => "0111111110100000",
56403 => "0111111110100000",
56404 => "0111111110100000",
56405 => "0111111110100000",
56406 => "0111111110100000",
56407 => "0111111110100000",
56408 => "0111111110100000",
56409 => "0111111110100000",
56410 => "0111111110100000",
56411 => "0111111110100000",
56412 => "0111111110100000",
56413 => "0111111110100000",
56414 => "0111111110100000",
56415 => "0111111110100000",
56416 => "0111111110100000",
56417 => "0111111110100000",
56418 => "0111111110100000",
56419 => "0111111110100000",
56420 => "0111111110100000",
56421 => "0111111110100000",
56422 => "0111111110100000",
56423 => "0111111110100000",
56424 => "0111111110100000",
56425 => "0111111110100000",
56426 => "0111111110100000",
56427 => "0111111110100000",
56428 => "0111111110100000",
56429 => "0111111110100000",
56430 => "0111111110100000",
56431 => "0111111110100000",
56432 => "0111111110100000",
56433 => "0111111110100000",
56434 => "0111111110100000",
56435 => "0111111110100000",
56436 => "0111111110100000",
56437 => "0111111110100000",
56438 => "0111111110100000",
56439 => "0111111110100000",
56440 => "0111111110100000",
56441 => "0111111110100000",
56442 => "0111111110100000",
56443 => "0111111110100000",
56444 => "0111111110100000",
56445 => "0111111110100000",
56446 => "0111111110100000",
56447 => "0111111110100000",
56448 => "0111111110100000",
56449 => "0111111110100000",
56450 => "0111111110100000",
56451 => "0111111110100000",
56452 => "0111111110100000",
56453 => "0111111110100000",
56454 => "0111111110100000",
56455 => "0111111110100000",
56456 => "0111111110100000",
56457 => "0111111110100000",
56458 => "0111111110100000",
56459 => "0111111110100000",
56460 => "0111111110100000",
56461 => "0111111110100000",
56462 => "0111111110100000",
56463 => "0111111110100000",
56464 => "0111111110100000",
56465 => "0111111110100000",
56466 => "0111111110100000",
56467 => "0111111110100000",
56468 => "0111111110100000",
56469 => "0111111110100000",
56470 => "0111111110100000",
56471 => "0111111110100000",
56472 => "0111111110100000",
56473 => "0111111110100000",
56474 => "0111111110100000",
56475 => "0111111110100000",
56476 => "0111111110100000",
56477 => "0111111110100000",
56478 => "0111111110100000",
56479 => "0111111110100000",
56480 => "0111111110100000",
56481 => "0111111110100000",
56482 => "0111111110100000",
56483 => "0111111110100000",
56484 => "0111111110100000",
56485 => "0111111110100000",
56486 => "0111111110100000",
56487 => "0111111110100000",
56488 => "0111111110100000",
56489 => "0111111110100000",
56490 => "0111111110100000",
56491 => "0111111110100000",
56492 => "0111111110100000",
56493 => "0111111110100000",
56494 => "0111111110100000",
56495 => "0111111110100000",
56496 => "0111111110100000",
56497 => "0111111110100000",
56498 => "0111111110100000",
56499 => "0111111110100000",
56500 => "0111111110100000",
56501 => "0111111110100000",
56502 => "0111111110100000",
56503 => "0111111110100000",
56504 => "0111111110100000",
56505 => "0111111110100000",
56506 => "0111111110100000",
56507 => "0111111110100000",
56508 => "0111111110100000",
56509 => "0111111110100000",
56510 => "0111111110100000",
56511 => "0111111110100000",
56512 => "0111111110100000",
56513 => "0111111110100000",
56514 => "0111111110100000",
56515 => "0111111110100000",
56516 => "0111111110100000",
56517 => "0111111110100000",
56518 => "0111111110100000",
56519 => "0111111110100000",
56520 => "0111111110100000",
56521 => "0111111110100000",
56522 => "0111111110100000",
56523 => "0111111110100000",
56524 => "0111111110100000",
56525 => "0111111110100000",
56526 => "0111111110100000",
56527 => "0111111110100000",
56528 => "0111111110100000",
56529 => "0111111110100000",
56530 => "0111111110100000",
56531 => "0111111110100000",
56532 => "0111111110100000",
56533 => "0111111110100000",
56534 => "0111111110100000",
56535 => "0111111110100000",
56536 => "0111111110100000",
56537 => "0111111110100000",
56538 => "0111111110100000",
56539 => "0111111110100000",
56540 => "0111111110100000",
56541 => "0111111110100000",
56542 => "0111111110100000",
56543 => "0111111110100000",
56544 => "0111111110100000",
56545 => "0111111110100000",
56546 => "0111111110100000",
56547 => "0111111110100000",
56548 => "0111111110100000",
56549 => "0111111110100000",
56550 => "0111111110100000",
56551 => "0111111110100000",
56552 => "0111111110100000",
56553 => "0111111110100000",
56554 => "0111111110100000",
56555 => "0111111110100000",
56556 => "0111111110100000",
56557 => "0111111110100000",
56558 => "0111111110100000",
56559 => "0111111110100000",
56560 => "0111111110100000",
56561 => "0111111110100000",
56562 => "0111111110100000",
56563 => "0111111110100000",
56564 => "0111111110100000",
56565 => "0111111110100000",
56566 => "0111111110100000",
56567 => "0111111110100000",
56568 => "0111111110100000",
56569 => "0111111110100000",
56570 => "0111111110100000",
56571 => "0111111110100000",
56572 => "0111111110100000",
56573 => "0111111110100000",
56574 => "0111111110100000",
56575 => "0111111110100000",
56576 => "0111111110100000",
56577 => "0111111110100000",
56578 => "0111111110100000",
56579 => "0111111110100000",
56580 => "0111111110100000",
56581 => "0111111110100000",
56582 => "0111111110100000",
56583 => "0111111110100000",
56584 => "0111111110100000",
56585 => "0111111110100000",
56586 => "0111111110100000",
56587 => "0111111110100000",
56588 => "0111111110100000",
56589 => "0111111110100000",
56590 => "0111111110100000",
56591 => "0111111110100000",
56592 => "0111111110100000",
56593 => "0111111110100000",
56594 => "0111111110100000",
56595 => "0111111110100000",
56596 => "0111111110100000",
56597 => "0111111110100000",
56598 => "0111111110100000",
56599 => "0111111110100000",
56600 => "0111111110100000",
56601 => "0111111110100000",
56602 => "0111111110100000",
56603 => "0111111110100000",
56604 => "0111111110100000",
56605 => "0111111110100000",
56606 => "0111111110100000",
56607 => "0111111110100000",
56608 => "0111111110100000",
56609 => "0111111110100000",
56610 => "0111111110100000",
56611 => "0111111110100000",
56612 => "0111111110100000",
56613 => "0111111110100000",
56614 => "0111111110100000",
56615 => "0111111110100000",
56616 => "0111111110100000",
56617 => "0111111110100000",
56618 => "0111111110100000",
56619 => "0111111110100000",
56620 => "0111111110100000",
56621 => "0111111110100000",
56622 => "0111111110100000",
56623 => "0111111110100000",
56624 => "0111111110100000",
56625 => "0111111110100000",
56626 => "0111111110100000",
56627 => "0111111110100000",
56628 => "0111111110100000",
56629 => "0111111110100000",
56630 => "0111111110100000",
56631 => "0111111110100000",
56632 => "0111111110100000",
56633 => "0111111110100000",
56634 => "0111111110100000",
56635 => "0111111110100000",
56636 => "0111111110100000",
56637 => "0111111110100000",
56638 => "0111111110100000",
56639 => "0111111110100000",
56640 => "0111111110100000",
56641 => "0111111110100000",
56642 => "0111111110100000",
56643 => "0111111110100000",
56644 => "0111111110100000",
56645 => "0111111110100000",
56646 => "0111111110100000",
56647 => "0111111110100000",
56648 => "0111111110100000",
56649 => "0111111110100000",
56650 => "0111111110100000",
56651 => "0111111110100000",
56652 => "0111111110100000",
56653 => "0111111110100000",
56654 => "0111111110100000",
56655 => "0111111110100000",
56656 => "0111111110100000",
56657 => "0111111110100000",
56658 => "0111111110100000",
56659 => "0111111110100000",
56660 => "0111111110100000",
56661 => "0111111110100000",
56662 => "0111111110100000",
56663 => "0111111110100000",
56664 => "0111111110100000",
56665 => "0111111110100000",
56666 => "0111111110100000",
56667 => "0111111110100000",
56668 => "0111111110100000",
56669 => "0111111110100000",
56670 => "0111111110100000",
56671 => "0111111110100000",
56672 => "0111111110100000",
56673 => "0111111110100000",
56674 => "0111111110100000",
56675 => "0111111110100000",
56676 => "0111111110100000",
56677 => "0111111110100000",
56678 => "0111111110100000",
56679 => "0111111110100000",
56680 => "0111111110100000",
56681 => "0111111110100000",
56682 => "0111111110100000",
56683 => "0111111110100000",
56684 => "0111111110100000",
56685 => "0111111110100000",
56686 => "0111111110100000",
56687 => "0111111110100000",
56688 => "0111111110100000",
56689 => "0111111110100000",
56690 => "0111111110100000",
56691 => "0111111110100000",
56692 => "0111111110100000",
56693 => "0111111110100000",
56694 => "0111111110100000",
56695 => "0111111110100000",
56696 => "0111111110100000",
56697 => "0111111110100000",
56698 => "0111111110100000",
56699 => "0111111110100000",
56700 => "0111111110100000",
56701 => "0111111110100000",
56702 => "0111111110100000",
56703 => "0111111110100000",
56704 => "0111111110100000",
56705 => "0111111110100000",
56706 => "0111111110100000",
56707 => "0111111110100000",
56708 => "0111111110100000",
56709 => "0111111110100000",
56710 => "0111111110100000",
56711 => "0111111110100000",
56712 => "0111111110100000",
56713 => "0111111110100000",
56714 => "0111111110100000",
56715 => "0111111110100000",
56716 => "0111111110100000",
56717 => "0111111110100000",
56718 => "0111111110100000",
56719 => "0111111110100000",
56720 => "0111111110100000",
56721 => "0111111110100000",
56722 => "0111111110100000",
56723 => "0111111110100000",
56724 => "0111111110100000",
56725 => "0111111110100000",
56726 => "0111111110100000",
56727 => "0111111110100000",
56728 => "0111111110100000",
56729 => "0111111110100000",
56730 => "0111111110100000",
56731 => "0111111110100000",
56732 => "0111111110100000",
56733 => "0111111110100000",
56734 => "0111111110100000",
56735 => "0111111110100000",
56736 => "0111111110100000",
56737 => "0111111110100000",
56738 => "0111111110100000",
56739 => "0111111110100000",
56740 => "0111111110100000",
56741 => "0111111110100000",
56742 => "0111111110100000",
56743 => "0111111110100000",
56744 => "0111111110100000",
56745 => "0111111110100000",
56746 => "0111111110100000",
56747 => "0111111110100000",
56748 => "0111111110100000",
56749 => "0111111110100000",
56750 => "0111111110100000",
56751 => "0111111110100000",
56752 => "0111111110100000",
56753 => "0111111110100000",
56754 => "0111111110100000",
56755 => "0111111110100000",
56756 => "0111111110100000",
56757 => "0111111110100000",
56758 => "0111111110100000",
56759 => "0111111110100000",
56760 => "0111111110100000",
56761 => "0111111110100000",
56762 => "0111111110100000",
56763 => "0111111110100000",
56764 => "0111111110100000",
56765 => "0111111110100000",
56766 => "0111111110100000",
56767 => "0111111110100000",
56768 => "0111111110100000",
56769 => "0111111110100000",
56770 => "0111111110100000",
56771 => "0111111110100000",
56772 => "0111111110100000",
56773 => "0111111110100000",
56774 => "0111111110100000",
56775 => "0111111110100000",
56776 => "0111111110100000",
56777 => "0111111110100000",
56778 => "0111111110100000",
56779 => "0111111110100000",
56780 => "0111111110100000",
56781 => "0111111110100000",
56782 => "0111111110100000",
56783 => "0111111110100000",
56784 => "0111111110100000",
56785 => "0111111110100000",
56786 => "0111111110100000",
56787 => "0111111110100000",
56788 => "0111111110100000",
56789 => "0111111110100000",
56790 => "0111111110100000",
56791 => "0111111110100000",
56792 => "0111111110100000",
56793 => "0111111110100000",
56794 => "0111111110100000",
56795 => "0111111110100000",
56796 => "0111111110100000",
56797 => "0111111110100000",
56798 => "0111111110100000",
56799 => "0111111110100000",
56800 => "0111111110100000",
56801 => "0111111110100000",
56802 => "0111111110100000",
56803 => "0111111110100000",
56804 => "0111111110100000",
56805 => "0111111110100000",
56806 => "0111111110100000",
56807 => "0111111110100000",
56808 => "0111111110100000",
56809 => "0111111110100000",
56810 => "0111111110100000",
56811 => "0111111110100000",
56812 => "0111111110100000",
56813 => "0111111110100000",
56814 => "0111111110100000",
56815 => "0111111110100000",
56816 => "0111111110100000",
56817 => "0111111110100000",
56818 => "0111111110100000",
56819 => "0111111110100000",
56820 => "0111111110100000",
56821 => "0111111110100000",
56822 => "0111111110100000",
56823 => "0111111110100000",
56824 => "0111111110100000",
56825 => "0111111110100000",
56826 => "0111111110100000",
56827 => "0111111110100000",
56828 => "0111111110100000",
56829 => "0111111110100000",
56830 => "0111111110100000",
56831 => "0111111110100000",
56832 => "0111111110100000",
56833 => "0111111110100000",
56834 => "0111111110100000",
56835 => "0111111110100000",
56836 => "0111111110100000",
56837 => "0111111110100000",
56838 => "0111111110100000",
56839 => "0111111110100000",
56840 => "0111111110100000",
56841 => "0111111110100000",
56842 => "0111111110100000",
56843 => "0111111110100000",
56844 => "0111111110100000",
56845 => "0111111110100000",
56846 => "0111111110100000",
56847 => "0111111110100000",
56848 => "0111111110100000",
56849 => "0111111110100000",
56850 => "0111111110100000",
56851 => "0111111110100000",
56852 => "0111111110100000",
56853 => "0111111110100000",
56854 => "0111111110100000",
56855 => "0111111110100000",
56856 => "0111111110100000",
56857 => "0111111110100000",
56858 => "0111111110100000",
56859 => "0111111110100000",
56860 => "0111111110100000",
56861 => "0111111110100000",
56862 => "0111111110100000",
56863 => "0111111110100000",
56864 => "0111111110100000",
56865 => "0111111110100000",
56866 => "0111111110100000",
56867 => "0111111110100000",
56868 => "0111111110100000",
56869 => "0111111110100000",
56870 => "0111111110100000",
56871 => "0111111110100000",
56872 => "0111111110100000",
56873 => "0111111110100000",
56874 => "0111111110100000",
56875 => "0111111110100000",
56876 => "0111111110100000",
56877 => "0111111110100000",
56878 => "0111111110100000",
56879 => "0111111110100000",
56880 => "0111111110100000",
56881 => "0111111110100000",
56882 => "0111111110100000",
56883 => "0111111110100000",
56884 => "0111111110100000",
56885 => "0111111110100000",
56886 => "0111111110100000",
56887 => "0111111110100000",
56888 => "0111111110100000",
56889 => "0111111110100000",
56890 => "0111111110100000",
56891 => "0111111110100000",
56892 => "0111111110100000",
56893 => "0111111110100000",
56894 => "0111111110100000",
56895 => "0111111110100000",
56896 => "0111111110100000",
56897 => "0111111110100000",
56898 => "0111111110100000",
56899 => "0111111110100000",
56900 => "0111111110100000",
56901 => "0111111110100000",
56902 => "0111111110100000",
56903 => "0111111110100000",
56904 => "0111111110100000",
56905 => "0111111110100000",
56906 => "0111111110100000",
56907 => "0111111110100000",
56908 => "0111111110100000",
56909 => "0111111110100000",
56910 => "0111111110100000",
56911 => "0111111110100000",
56912 => "0111111110100000",
56913 => "0111111110100000",
56914 => "0111111110100000",
56915 => "0111111110100000",
56916 => "0111111110100000",
56917 => "0111111110100000",
56918 => "0111111110100000",
56919 => "0111111110100000",
56920 => "0111111110100000",
56921 => "0111111110100000",
56922 => "0111111110100000",
56923 => "0111111110100000",
56924 => "0111111110100000",
56925 => "0111111110100000",
56926 => "0111111110100000",
56927 => "0111111110100000",
56928 => "0111111110100000",
56929 => "0111111110100000",
56930 => "0111111110100000",
56931 => "0111111110100000",
56932 => "0111111110100000",
56933 => "0111111110100000",
56934 => "0111111110100000",
56935 => "0111111110100000",
56936 => "0111111110100000",
56937 => "0111111110100000",
56938 => "0111111110100000",
56939 => "0111111110100000",
56940 => "0111111110100000",
56941 => "0111111110100000",
56942 => "0111111110100000",
56943 => "0111111110100000",
56944 => "0111111110100000",
56945 => "0111111110100000",
56946 => "0111111110100000",
56947 => "0111111110100000",
56948 => "0111111110100000",
56949 => "0111111110100000",
56950 => "0111111110100000",
56951 => "0111111110100000",
56952 => "0111111110100000",
56953 => "0111111110100000",
56954 => "0111111110100000",
56955 => "0111111110100000",
56956 => "0111111110100000",
56957 => "0111111110100000",
56958 => "0111111110100000",
56959 => "0111111110100000",
56960 => "0111111110100000",
56961 => "0111111110100000",
56962 => "0111111110100000",
56963 => "0111111110100000",
56964 => "0111111110100000",
56965 => "0111111110100000",
56966 => "0111111110100000",
56967 => "0111111110100000",
56968 => "0111111110100000",
56969 => "0111111110100000",
56970 => "0111111110100000",
56971 => "0111111110100000",
56972 => "0111111110100000",
56973 => "0111111110100000",
56974 => "0111111110100000",
56975 => "0111111110100000",
56976 => "0111111110100000",
56977 => "0111111110100000",
56978 => "0111111110100000",
56979 => "0111111110100000",
56980 => "0111111110100000",
56981 => "0111111110100000",
56982 => "0111111110100000",
56983 => "0111111110100000",
56984 => "0111111110100000",
56985 => "0111111110100000",
56986 => "0111111110100000",
56987 => "0111111110100000",
56988 => "0111111110100000",
56989 => "0111111110100000",
56990 => "0111111110100000",
56991 => "0111111110100000",
56992 => "0111111110100000",
56993 => "0111111110100000",
56994 => "0111111110100000",
56995 => "0111111110100000",
56996 => "0111111110100000",
56997 => "0111111110100000",
56998 => "0111111110100000",
56999 => "0111111110100000",
57000 => "0111111110100000",
57001 => "0111111110100000",
57002 => "0111111110100000",
57003 => "0111111110100000",
57004 => "0111111110110000",
57005 => "0111111110110000",
57006 => "0111111110110000",
57007 => "0111111110110000",
57008 => "0111111110110000",
57009 => "0111111110110000",
57010 => "0111111110110000",
57011 => "0111111110110000",
57012 => "0111111110110000",
57013 => "0111111110110000",
57014 => "0111111110110000",
57015 => "0111111110110000",
57016 => "0111111110110000",
57017 => "0111111110110000",
57018 => "0111111110110000",
57019 => "0111111110110000",
57020 => "0111111110110000",
57021 => "0111111110110000",
57022 => "0111111110110000",
57023 => "0111111110110000",
57024 => "0111111110110000",
57025 => "0111111110110000",
57026 => "0111111110110000",
57027 => "0111111110110000",
57028 => "0111111110110000",
57029 => "0111111110110000",
57030 => "0111111110110000",
57031 => "0111111110110000",
57032 => "0111111110110000",
57033 => "0111111110110000",
57034 => "0111111110110000",
57035 => "0111111110110000",
57036 => "0111111110110000",
57037 => "0111111110110000",
57038 => "0111111110110000",
57039 => "0111111110110000",
57040 => "0111111110110000",
57041 => "0111111110110000",
57042 => "0111111110110000",
57043 => "0111111110110000",
57044 => "0111111110110000",
57045 => "0111111110110000",
57046 => "0111111110110000",
57047 => "0111111110110000",
57048 => "0111111110110000",
57049 => "0111111110110000",
57050 => "0111111110110000",
57051 => "0111111110110000",
57052 => "0111111110110000",
57053 => "0111111110110000",
57054 => "0111111110110000",
57055 => "0111111110110000",
57056 => "0111111110110000",
57057 => "0111111110110000",
57058 => "0111111110110000",
57059 => "0111111110110000",
57060 => "0111111110110000",
57061 => "0111111110110000",
57062 => "0111111110110000",
57063 => "0111111110110000",
57064 => "0111111110110000",
57065 => "0111111110110000",
57066 => "0111111110110000",
57067 => "0111111110110000",
57068 => "0111111110110000",
57069 => "0111111110110000",
57070 => "0111111110110000",
57071 => "0111111110110000",
57072 => "0111111110110000",
57073 => "0111111110110000",
57074 => "0111111110110000",
57075 => "0111111110110000",
57076 => "0111111110110000",
57077 => "0111111110110000",
57078 => "0111111110110000",
57079 => "0111111110110000",
57080 => "0111111110110000",
57081 => "0111111110110000",
57082 => "0111111110110000",
57083 => "0111111110110000",
57084 => "0111111110110000",
57085 => "0111111110110000",
57086 => "0111111110110000",
57087 => "0111111110110000",
57088 => "0111111110110000",
57089 => "0111111110110000",
57090 => "0111111110110000",
57091 => "0111111110110000",
57092 => "0111111110110000",
57093 => "0111111110110000",
57094 => "0111111110110000",
57095 => "0111111110110000",
57096 => "0111111110110000",
57097 => "0111111110110000",
57098 => "0111111110110000",
57099 => "0111111110110000",
57100 => "0111111110110000",
57101 => "0111111110110000",
57102 => "0111111110110000",
57103 => "0111111110110000",
57104 => "0111111110110000",
57105 => "0111111110110000",
57106 => "0111111110110000",
57107 => "0111111110110000",
57108 => "0111111110110000",
57109 => "0111111110110000",
57110 => "0111111110110000",
57111 => "0111111110110000",
57112 => "0111111110110000",
57113 => "0111111110110000",
57114 => "0111111110110000",
57115 => "0111111110110000",
57116 => "0111111110110000",
57117 => "0111111110110000",
57118 => "0111111110110000",
57119 => "0111111110110000",
57120 => "0111111110110000",
57121 => "0111111110110000",
57122 => "0111111110110000",
57123 => "0111111110110000",
57124 => "0111111110110000",
57125 => "0111111110110000",
57126 => "0111111110110000",
57127 => "0111111110110000",
57128 => "0111111110110000",
57129 => "0111111110110000",
57130 => "0111111110110000",
57131 => "0111111110110000",
57132 => "0111111110110000",
57133 => "0111111110110000",
57134 => "0111111110110000",
57135 => "0111111110110000",
57136 => "0111111110110000",
57137 => "0111111110110000",
57138 => "0111111110110000",
57139 => "0111111110110000",
57140 => "0111111110110000",
57141 => "0111111110110000",
57142 => "0111111110110000",
57143 => "0111111110110000",
57144 => "0111111110110000",
57145 => "0111111110110000",
57146 => "0111111110110000",
57147 => "0111111110110000",
57148 => "0111111110110000",
57149 => "0111111110110000",
57150 => "0111111110110000",
57151 => "0111111110110000",
57152 => "0111111110110000",
57153 => "0111111110110000",
57154 => "0111111110110000",
57155 => "0111111110110000",
57156 => "0111111110110000",
57157 => "0111111110110000",
57158 => "0111111110110000",
57159 => "0111111110110000",
57160 => "0111111110110000",
57161 => "0111111110110000",
57162 => "0111111110110000",
57163 => "0111111110110000",
57164 => "0111111110110000",
57165 => "0111111110110000",
57166 => "0111111110110000",
57167 => "0111111110110000",
57168 => "0111111110110000",
57169 => "0111111110110000",
57170 => "0111111110110000",
57171 => "0111111110110000",
57172 => "0111111110110000",
57173 => "0111111110110000",
57174 => "0111111110110000",
57175 => "0111111110110000",
57176 => "0111111110110000",
57177 => "0111111110110000",
57178 => "0111111110110000",
57179 => "0111111110110000",
57180 => "0111111110110000",
57181 => "0111111110110000",
57182 => "0111111110110000",
57183 => "0111111110110000",
57184 => "0111111110110000",
57185 => "0111111110110000",
57186 => "0111111110110000",
57187 => "0111111110110000",
57188 => "0111111110110000",
57189 => "0111111110110000",
57190 => "0111111110110000",
57191 => "0111111110110000",
57192 => "0111111110110000",
57193 => "0111111110110000",
57194 => "0111111110110000",
57195 => "0111111110110000",
57196 => "0111111110110000",
57197 => "0111111110110000",
57198 => "0111111110110000",
57199 => "0111111110110000",
57200 => "0111111110110000",
57201 => "0111111110110000",
57202 => "0111111110110000",
57203 => "0111111110110000",
57204 => "0111111110110000",
57205 => "0111111110110000",
57206 => "0111111110110000",
57207 => "0111111110110000",
57208 => "0111111110110000",
57209 => "0111111110110000",
57210 => "0111111110110000",
57211 => "0111111110110000",
57212 => "0111111110110000",
57213 => "0111111110110000",
57214 => "0111111110110000",
57215 => "0111111110110000",
57216 => "0111111110110000",
57217 => "0111111110110000",
57218 => "0111111110110000",
57219 => "0111111110110000",
57220 => "0111111110110000",
57221 => "0111111110110000",
57222 => "0111111110110000",
57223 => "0111111110110000",
57224 => "0111111110110000",
57225 => "0111111110110000",
57226 => "0111111110110000",
57227 => "0111111110110000",
57228 => "0111111110110000",
57229 => "0111111110110000",
57230 => "0111111110110000",
57231 => "0111111110110000",
57232 => "0111111110110000",
57233 => "0111111110110000",
57234 => "0111111110110000",
57235 => "0111111110110000",
57236 => "0111111110110000",
57237 => "0111111110110000",
57238 => "0111111110110000",
57239 => "0111111110110000",
57240 => "0111111110110000",
57241 => "0111111110110000",
57242 => "0111111110110000",
57243 => "0111111110110000",
57244 => "0111111110110000",
57245 => "0111111110110000",
57246 => "0111111110110000",
57247 => "0111111110110000",
57248 => "0111111110110000",
57249 => "0111111110110000",
57250 => "0111111110110000",
57251 => "0111111110110000",
57252 => "0111111110110000",
57253 => "0111111110110000",
57254 => "0111111110110000",
57255 => "0111111110110000",
57256 => "0111111110110000",
57257 => "0111111110110000",
57258 => "0111111110110000",
57259 => "0111111110110000",
57260 => "0111111110110000",
57261 => "0111111110110000",
57262 => "0111111110110000",
57263 => "0111111110110000",
57264 => "0111111110110000",
57265 => "0111111110110000",
57266 => "0111111110110000",
57267 => "0111111110110000",
57268 => "0111111110110000",
57269 => "0111111110110000",
57270 => "0111111110110000",
57271 => "0111111110110000",
57272 => "0111111110110000",
57273 => "0111111110110000",
57274 => "0111111110110000",
57275 => "0111111110110000",
57276 => "0111111110110000",
57277 => "0111111110110000",
57278 => "0111111110110000",
57279 => "0111111110110000",
57280 => "0111111110110000",
57281 => "0111111110110000",
57282 => "0111111110110000",
57283 => "0111111110110000",
57284 => "0111111110110000",
57285 => "0111111110110000",
57286 => "0111111110110000",
57287 => "0111111110110000",
57288 => "0111111110110000",
57289 => "0111111110110000",
57290 => "0111111110110000",
57291 => "0111111110110000",
57292 => "0111111110110000",
57293 => "0111111110110000",
57294 => "0111111110110000",
57295 => "0111111110110000",
57296 => "0111111110110000",
57297 => "0111111110110000",
57298 => "0111111110110000",
57299 => "0111111110110000",
57300 => "0111111110110000",
57301 => "0111111110110000",
57302 => "0111111110110000",
57303 => "0111111110110000",
57304 => "0111111110110000",
57305 => "0111111110110000",
57306 => "0111111110110000",
57307 => "0111111110110000",
57308 => "0111111110110000",
57309 => "0111111110110000",
57310 => "0111111110110000",
57311 => "0111111110110000",
57312 => "0111111110110000",
57313 => "0111111110110000",
57314 => "0111111110110000",
57315 => "0111111110110000",
57316 => "0111111110110000",
57317 => "0111111110110000",
57318 => "0111111110110000",
57319 => "0111111110110000",
57320 => "0111111110110000",
57321 => "0111111110110000",
57322 => "0111111110110000",
57323 => "0111111110110000",
57324 => "0111111110110000",
57325 => "0111111110110000",
57326 => "0111111110110000",
57327 => "0111111110110000",
57328 => "0111111110110000",
57329 => "0111111110110000",
57330 => "0111111110110000",
57331 => "0111111110110000",
57332 => "0111111110110000",
57333 => "0111111110110000",
57334 => "0111111110110000",
57335 => "0111111110110000",
57336 => "0111111110110000",
57337 => "0111111110110000",
57338 => "0111111110110000",
57339 => "0111111110110000",
57340 => "0111111110110000",
57341 => "0111111110110000",
57342 => "0111111110110000",
57343 => "0111111110110000",
57344 => "0111111110110000",
57345 => "0111111110110000",
57346 => "0111111110110000",
57347 => "0111111110110000",
57348 => "0111111110110000",
57349 => "0111111110110000",
57350 => "0111111110110000",
57351 => "0111111110110000",
57352 => "0111111110110000",
57353 => "0111111110110000",
57354 => "0111111110110000",
57355 => "0111111110110000",
57356 => "0111111110110000",
57357 => "0111111110110000",
57358 => "0111111110110000",
57359 => "0111111110110000",
57360 => "0111111110110000",
57361 => "0111111110110000",
57362 => "0111111110110000",
57363 => "0111111110110000",
57364 => "0111111110110000",
57365 => "0111111110110000",
57366 => "0111111110110000",
57367 => "0111111110110000",
57368 => "0111111110110000",
57369 => "0111111110110000",
57370 => "0111111110110000",
57371 => "0111111110110000",
57372 => "0111111110110000",
57373 => "0111111110110000",
57374 => "0111111110110000",
57375 => "0111111110110000",
57376 => "0111111110110000",
57377 => "0111111110110000",
57378 => "0111111110110000",
57379 => "0111111110110000",
57380 => "0111111110110000",
57381 => "0111111110110000",
57382 => "0111111110110000",
57383 => "0111111110110000",
57384 => "0111111110110000",
57385 => "0111111110110000",
57386 => "0111111110110000",
57387 => "0111111110110000",
57388 => "0111111110110000",
57389 => "0111111110110000",
57390 => "0111111110110000",
57391 => "0111111110110000",
57392 => "0111111110110000",
57393 => "0111111110110000",
57394 => "0111111110110000",
57395 => "0111111110110000",
57396 => "0111111110110000",
57397 => "0111111110110000",
57398 => "0111111110110000",
57399 => "0111111110110000",
57400 => "0111111110110000",
57401 => "0111111110110000",
57402 => "0111111110110000",
57403 => "0111111110110000",
57404 => "0111111110110000",
57405 => "0111111110110000",
57406 => "0111111110110000",
57407 => "0111111110110000",
57408 => "0111111110110000",
57409 => "0111111110110000",
57410 => "0111111110110000",
57411 => "0111111110110000",
57412 => "0111111110110000",
57413 => "0111111110110000",
57414 => "0111111110110000",
57415 => "0111111110110000",
57416 => "0111111110110000",
57417 => "0111111110110000",
57418 => "0111111110110000",
57419 => "0111111110110000",
57420 => "0111111110110000",
57421 => "0111111110110000",
57422 => "0111111110110000",
57423 => "0111111110110000",
57424 => "0111111110110000",
57425 => "0111111110110000",
57426 => "0111111110110000",
57427 => "0111111110110000",
57428 => "0111111110110000",
57429 => "0111111110110000",
57430 => "0111111110110000",
57431 => "0111111110110000",
57432 => "0111111110110000",
57433 => "0111111110110000",
57434 => "0111111110110000",
57435 => "0111111110110000",
57436 => "0111111110110000",
57437 => "0111111110110000",
57438 => "0111111110110000",
57439 => "0111111110110000",
57440 => "0111111110110000",
57441 => "0111111110110000",
57442 => "0111111110110000",
57443 => "0111111110110000",
57444 => "0111111110110000",
57445 => "0111111110110000",
57446 => "0111111110110000",
57447 => "0111111110110000",
57448 => "0111111110110000",
57449 => "0111111110110000",
57450 => "0111111110110000",
57451 => "0111111110110000",
57452 => "0111111110110000",
57453 => "0111111110110000",
57454 => "0111111110110000",
57455 => "0111111110110000",
57456 => "0111111110110000",
57457 => "0111111110110000",
57458 => "0111111110110000",
57459 => "0111111110110000",
57460 => "0111111110110000",
57461 => "0111111110110000",
57462 => "0111111110110000",
57463 => "0111111110110000",
57464 => "0111111110110000",
57465 => "0111111110110000",
57466 => "0111111110110000",
57467 => "0111111110110000",
57468 => "0111111110110000",
57469 => "0111111110110000",
57470 => "0111111110110000",
57471 => "0111111110110000",
57472 => "0111111110110000",
57473 => "0111111110110000",
57474 => "0111111110110000",
57475 => "0111111110110000",
57476 => "0111111110110000",
57477 => "0111111110110000",
57478 => "0111111110110000",
57479 => "0111111110110000",
57480 => "0111111110110000",
57481 => "0111111110110000",
57482 => "0111111110110000",
57483 => "0111111110110000",
57484 => "0111111110110000",
57485 => "0111111110110000",
57486 => "0111111110110000",
57487 => "0111111110110000",
57488 => "0111111110110000",
57489 => "0111111110110000",
57490 => "0111111110110000",
57491 => "0111111110110000",
57492 => "0111111110110000",
57493 => "0111111110110000",
57494 => "0111111110110000",
57495 => "0111111110110000",
57496 => "0111111110110000",
57497 => "0111111110110000",
57498 => "0111111110110000",
57499 => "0111111110110000",
57500 => "0111111110110000",
57501 => "0111111110110000",
57502 => "0111111110110000",
57503 => "0111111110110000",
57504 => "0111111110110000",
57505 => "0111111110110000",
57506 => "0111111110110000",
57507 => "0111111110110000",
57508 => "0111111110110000",
57509 => "0111111110110000",
57510 => "0111111110110000",
57511 => "0111111110110000",
57512 => "0111111110110000",
57513 => "0111111110110000",
57514 => "0111111110110000",
57515 => "0111111110110000",
57516 => "0111111110110000",
57517 => "0111111110110000",
57518 => "0111111110110000",
57519 => "0111111110110000",
57520 => "0111111110110000",
57521 => "0111111110110000",
57522 => "0111111110110000",
57523 => "0111111110110000",
57524 => "0111111110110000",
57525 => "0111111110110000",
57526 => "0111111110110000",
57527 => "0111111110110000",
57528 => "0111111110110000",
57529 => "0111111110110000",
57530 => "0111111110110000",
57531 => "0111111110110000",
57532 => "0111111110110000",
57533 => "0111111110110000",
57534 => "0111111110110000",
57535 => "0111111110110000",
57536 => "0111111110110000",
57537 => "0111111110110000",
57538 => "0111111110110000",
57539 => "0111111110110000",
57540 => "0111111110110000",
57541 => "0111111110110000",
57542 => "0111111110110000",
57543 => "0111111110110000",
57544 => "0111111110110000",
57545 => "0111111110110000",
57546 => "0111111110110000",
57547 => "0111111110110000",
57548 => "0111111110110000",
57549 => "0111111110110000",
57550 => "0111111110110000",
57551 => "0111111110110000",
57552 => "0111111110110000",
57553 => "0111111110110000",
57554 => "0111111110110000",
57555 => "0111111110110000",
57556 => "0111111110110000",
57557 => "0111111110110000",
57558 => "0111111110110000",
57559 => "0111111110110000",
57560 => "0111111110110000",
57561 => "0111111110110000",
57562 => "0111111110110000",
57563 => "0111111110110000",
57564 => "0111111110110000",
57565 => "0111111110110000",
57566 => "0111111110110000",
57567 => "0111111110110000",
57568 => "0111111110110000",
57569 => "0111111110110000",
57570 => "0111111110110000",
57571 => "0111111110110000",
57572 => "0111111110110000",
57573 => "0111111110110000",
57574 => "0111111110110000",
57575 => "0111111110110000",
57576 => "0111111110110000",
57577 => "0111111110110000",
57578 => "0111111110110000",
57579 => "0111111110110000",
57580 => "0111111110110000",
57581 => "0111111110110000",
57582 => "0111111110110000",
57583 => "0111111110110000",
57584 => "0111111110110000",
57585 => "0111111110110000",
57586 => "0111111110110000",
57587 => "0111111110110000",
57588 => "0111111110110000",
57589 => "0111111110110000",
57590 => "0111111110110000",
57591 => "0111111110110000",
57592 => "0111111110110000",
57593 => "0111111110110000",
57594 => "0111111110110000",
57595 => "0111111110110000",
57596 => "0111111110110000",
57597 => "0111111110110000",
57598 => "0111111110110000",
57599 => "0111111110110000",
57600 => "0111111110110000",
57601 => "0111111110110000",
57602 => "0111111110110000",
57603 => "0111111110110000",
57604 => "0111111110110000",
57605 => "0111111110110000",
57606 => "0111111110110000",
57607 => "0111111110110000",
57608 => "0111111110110000",
57609 => "0111111110110000",
57610 => "0111111110110000",
57611 => "0111111110110000",
57612 => "0111111110110000",
57613 => "0111111110110000",
57614 => "0111111110110000",
57615 => "0111111110110000",
57616 => "0111111110110000",
57617 => "0111111110110000",
57618 => "0111111110110000",
57619 => "0111111110110000",
57620 => "0111111110110000",
57621 => "0111111110110000",
57622 => "0111111110110000",
57623 => "0111111110110000",
57624 => "0111111110110000",
57625 => "0111111110110000",
57626 => "0111111110110000",
57627 => "0111111110110000",
57628 => "0111111110110000",
57629 => "0111111110110000",
57630 => "0111111110110000",
57631 => "0111111110110000",
57632 => "0111111110110000",
57633 => "0111111110110000",
57634 => "0111111110110000",
57635 => "0111111110110000",
57636 => "0111111110110000",
57637 => "0111111110110000",
57638 => "0111111110110000",
57639 => "0111111110110000",
57640 => "0111111110110000",
57641 => "0111111110110000",
57642 => "0111111110110000",
57643 => "0111111110110000",
57644 => "0111111110110000",
57645 => "0111111110110000",
57646 => "0111111110110000",
57647 => "0111111110110000",
57648 => "0111111110110000",
57649 => "0111111110110000",
57650 => "0111111110110000",
57651 => "0111111110110000",
57652 => "0111111110110000",
57653 => "0111111110110000",
57654 => "0111111110110000",
57655 => "0111111110110000",
57656 => "0111111110110000",
57657 => "0111111110110000",
57658 => "0111111110110000",
57659 => "0111111110110000",
57660 => "0111111110110000",
57661 => "0111111110110000",
57662 => "0111111110110000",
57663 => "0111111110110000",
57664 => "0111111110110000",
57665 => "0111111110110000",
57666 => "0111111110110000",
57667 => "0111111110110000",
57668 => "0111111110110000",
57669 => "0111111110110000",
57670 => "0111111110110000",
57671 => "0111111110110000",
57672 => "0111111110110000",
57673 => "0111111110110000",
57674 => "0111111110110000",
57675 => "0111111110110000",
57676 => "0111111110110000",
57677 => "0111111110110000",
57678 => "0111111110110000",
57679 => "0111111110110000",
57680 => "0111111110110000",
57681 => "0111111110110000",
57682 => "0111111110110000",
57683 => "0111111110110000",
57684 => "0111111110110000",
57685 => "0111111110110000",
57686 => "0111111110110000",
57687 => "0111111110110000",
57688 => "0111111110110000",
57689 => "0111111110110000",
57690 => "0111111110110000",
57691 => "0111111110110000",
57692 => "0111111110110000",
57693 => "0111111110110000",
57694 => "0111111110110000",
57695 => "0111111110110000",
57696 => "0111111110110000",
57697 => "0111111110110000",
57698 => "0111111110110000",
57699 => "0111111110110000",
57700 => "0111111110110000",
57701 => "0111111110110000",
57702 => "0111111110110000",
57703 => "0111111110110000",
57704 => "0111111110110000",
57705 => "0111111110110000",
57706 => "0111111110110000",
57707 => "0111111110110000",
57708 => "0111111110110000",
57709 => "0111111110110000",
57710 => "0111111110110000",
57711 => "0111111110110000",
57712 => "0111111110110000",
57713 => "0111111110110000",
57714 => "0111111110110000",
57715 => "0111111110110000",
57716 => "0111111110110000",
57717 => "0111111110110000",
57718 => "0111111110110000",
57719 => "0111111110110000",
57720 => "0111111110110000",
57721 => "0111111110110000",
57722 => "0111111110110000",
57723 => "0111111110110000",
57724 => "0111111110110000",
57725 => "0111111110110000",
57726 => "0111111110110000",
57727 => "0111111110110000",
57728 => "0111111110110000",
57729 => "0111111110110000",
57730 => "0111111110110000",
57731 => "0111111110110000",
57732 => "0111111110110000",
57733 => "0111111110110000",
57734 => "0111111110110000",
57735 => "0111111110110000",
57736 => "0111111110110000",
57737 => "0111111110110000",
57738 => "0111111110110000",
57739 => "0111111110110000",
57740 => "0111111110110000",
57741 => "0111111110110000",
57742 => "0111111110110000",
57743 => "0111111110110000",
57744 => "0111111110110000",
57745 => "0111111110110000",
57746 => "0111111110110000",
57747 => "0111111110110000",
57748 => "0111111110110000",
57749 => "0111111110110000",
57750 => "0111111110110000",
57751 => "0111111110110000",
57752 => "0111111110110000",
57753 => "0111111110110000",
57754 => "0111111110110000",
57755 => "0111111110110000",
57756 => "0111111110110000",
57757 => "0111111110110000",
57758 => "0111111110110000",
57759 => "0111111110110000",
57760 => "0111111110110000",
57761 => "0111111110110000",
57762 => "0111111110110000",
57763 => "0111111110110000",
57764 => "0111111110110000",
57765 => "0111111110110000",
57766 => "0111111110110000",
57767 => "0111111110110000",
57768 => "0111111110110000",
57769 => "0111111110110000",
57770 => "0111111110110000",
57771 => "0111111110110000",
57772 => "0111111110110000",
57773 => "0111111110110000",
57774 => "0111111110110000",
57775 => "0111111110110000",
57776 => "0111111110110000",
57777 => "0111111110110000",
57778 => "0111111110110000",
57779 => "0111111110110000",
57780 => "0111111110110000",
57781 => "0111111110110000",
57782 => "0111111110110000",
57783 => "0111111110110000",
57784 => "0111111110110000",
57785 => "0111111110110000",
57786 => "0111111110110000",
57787 => "0111111110110000",
57788 => "0111111110110000",
57789 => "0111111110110000",
57790 => "0111111110110000",
57791 => "0111111110110000",
57792 => "0111111110110000",
57793 => "0111111110110000",
57794 => "0111111110110000",
57795 => "0111111110110000",
57796 => "0111111110110000",
57797 => "0111111110110000",
57798 => "0111111110110000",
57799 => "0111111110110000",
57800 => "0111111110110000",
57801 => "0111111110110000",
57802 => "0111111110110000",
57803 => "0111111110110000",
57804 => "0111111110110000",
57805 => "0111111110110000",
57806 => "0111111110110000",
57807 => "0111111110110000",
57808 => "0111111110110000",
57809 => "0111111110110000",
57810 => "0111111110110000",
57811 => "0111111110110000",
57812 => "0111111110110000",
57813 => "0111111110110000",
57814 => "0111111110110000",
57815 => "0111111110110000",
57816 => "0111111110110000",
57817 => "0111111110110000",
57818 => "0111111110110000",
57819 => "0111111110110000",
57820 => "0111111110110000",
57821 => "0111111110110000",
57822 => "0111111110110000",
57823 => "0111111110110000",
57824 => "0111111110110000",
57825 => "0111111110110000",
57826 => "0111111110110000",
57827 => "0111111110110000",
57828 => "0111111111000000",
57829 => "0111111111000000",
57830 => "0111111111000000",
57831 => "0111111111000000",
57832 => "0111111111000000",
57833 => "0111111111000000",
57834 => "0111111111000000",
57835 => "0111111111000000",
57836 => "0111111111000000",
57837 => "0111111111000000",
57838 => "0111111111000000",
57839 => "0111111111000000",
57840 => "0111111111000000",
57841 => "0111111111000000",
57842 => "0111111111000000",
57843 => "0111111111000000",
57844 => "0111111111000000",
57845 => "0111111111000000",
57846 => "0111111111000000",
57847 => "0111111111000000",
57848 => "0111111111000000",
57849 => "0111111111000000",
57850 => "0111111111000000",
57851 => "0111111111000000",
57852 => "0111111111000000",
57853 => "0111111111000000",
57854 => "0111111111000000",
57855 => "0111111111000000",
57856 => "0111111111000000",
57857 => "0111111111000000",
57858 => "0111111111000000",
57859 => "0111111111000000",
57860 => "0111111111000000",
57861 => "0111111111000000",
57862 => "0111111111000000",
57863 => "0111111111000000",
57864 => "0111111111000000",
57865 => "0111111111000000",
57866 => "0111111111000000",
57867 => "0111111111000000",
57868 => "0111111111000000",
57869 => "0111111111000000",
57870 => "0111111111000000",
57871 => "0111111111000000",
57872 => "0111111111000000",
57873 => "0111111111000000",
57874 => "0111111111000000",
57875 => "0111111111000000",
57876 => "0111111111000000",
57877 => "0111111111000000",
57878 => "0111111111000000",
57879 => "0111111111000000",
57880 => "0111111111000000",
57881 => "0111111111000000",
57882 => "0111111111000000",
57883 => "0111111111000000",
57884 => "0111111111000000",
57885 => "0111111111000000",
57886 => "0111111111000000",
57887 => "0111111111000000",
57888 => "0111111111000000",
57889 => "0111111111000000",
57890 => "0111111111000000",
57891 => "0111111111000000",
57892 => "0111111111000000",
57893 => "0111111111000000",
57894 => "0111111111000000",
57895 => "0111111111000000",
57896 => "0111111111000000",
57897 => "0111111111000000",
57898 => "0111111111000000",
57899 => "0111111111000000",
57900 => "0111111111000000",
57901 => "0111111111000000",
57902 => "0111111111000000",
57903 => "0111111111000000",
57904 => "0111111111000000",
57905 => "0111111111000000",
57906 => "0111111111000000",
57907 => "0111111111000000",
57908 => "0111111111000000",
57909 => "0111111111000000",
57910 => "0111111111000000",
57911 => "0111111111000000",
57912 => "0111111111000000",
57913 => "0111111111000000",
57914 => "0111111111000000",
57915 => "0111111111000000",
57916 => "0111111111000000",
57917 => "0111111111000000",
57918 => "0111111111000000",
57919 => "0111111111000000",
57920 => "0111111111000000",
57921 => "0111111111000000",
57922 => "0111111111000000",
57923 => "0111111111000000",
57924 => "0111111111000000",
57925 => "0111111111000000",
57926 => "0111111111000000",
57927 => "0111111111000000",
57928 => "0111111111000000",
57929 => "0111111111000000",
57930 => "0111111111000000",
57931 => "0111111111000000",
57932 => "0111111111000000",
57933 => "0111111111000000",
57934 => "0111111111000000",
57935 => "0111111111000000",
57936 => "0111111111000000",
57937 => "0111111111000000",
57938 => "0111111111000000",
57939 => "0111111111000000",
57940 => "0111111111000000",
57941 => "0111111111000000",
57942 => "0111111111000000",
57943 => "0111111111000000",
57944 => "0111111111000000",
57945 => "0111111111000000",
57946 => "0111111111000000",
57947 => "0111111111000000",
57948 => "0111111111000000",
57949 => "0111111111000000",
57950 => "0111111111000000",
57951 => "0111111111000000",
57952 => "0111111111000000",
57953 => "0111111111000000",
57954 => "0111111111000000",
57955 => "0111111111000000",
57956 => "0111111111000000",
57957 => "0111111111000000",
57958 => "0111111111000000",
57959 => "0111111111000000",
57960 => "0111111111000000",
57961 => "0111111111000000",
57962 => "0111111111000000",
57963 => "0111111111000000",
57964 => "0111111111000000",
57965 => "0111111111000000",
57966 => "0111111111000000",
57967 => "0111111111000000",
57968 => "0111111111000000",
57969 => "0111111111000000",
57970 => "0111111111000000",
57971 => "0111111111000000",
57972 => "0111111111000000",
57973 => "0111111111000000",
57974 => "0111111111000000",
57975 => "0111111111000000",
57976 => "0111111111000000",
57977 => "0111111111000000",
57978 => "0111111111000000",
57979 => "0111111111000000",
57980 => "0111111111000000",
57981 => "0111111111000000",
57982 => "0111111111000000",
57983 => "0111111111000000",
57984 => "0111111111000000",
57985 => "0111111111000000",
57986 => "0111111111000000",
57987 => "0111111111000000",
57988 => "0111111111000000",
57989 => "0111111111000000",
57990 => "0111111111000000",
57991 => "0111111111000000",
57992 => "0111111111000000",
57993 => "0111111111000000",
57994 => "0111111111000000",
57995 => "0111111111000000",
57996 => "0111111111000000",
57997 => "0111111111000000",
57998 => "0111111111000000",
57999 => "0111111111000000",
58000 => "0111111111000000",
58001 => "0111111111000000",
58002 => "0111111111000000",
58003 => "0111111111000000",
58004 => "0111111111000000",
58005 => "0111111111000000",
58006 => "0111111111000000",
58007 => "0111111111000000",
58008 => "0111111111000000",
58009 => "0111111111000000",
58010 => "0111111111000000",
58011 => "0111111111000000",
58012 => "0111111111000000",
58013 => "0111111111000000",
58014 => "0111111111000000",
58015 => "0111111111000000",
58016 => "0111111111000000",
58017 => "0111111111000000",
58018 => "0111111111000000",
58019 => "0111111111000000",
58020 => "0111111111000000",
58021 => "0111111111000000",
58022 => "0111111111000000",
58023 => "0111111111000000",
58024 => "0111111111000000",
58025 => "0111111111000000",
58026 => "0111111111000000",
58027 => "0111111111000000",
58028 => "0111111111000000",
58029 => "0111111111000000",
58030 => "0111111111000000",
58031 => "0111111111000000",
58032 => "0111111111000000",
58033 => "0111111111000000",
58034 => "0111111111000000",
58035 => "0111111111000000",
58036 => "0111111111000000",
58037 => "0111111111000000",
58038 => "0111111111000000",
58039 => "0111111111000000",
58040 => "0111111111000000",
58041 => "0111111111000000",
58042 => "0111111111000000",
58043 => "0111111111000000",
58044 => "0111111111000000",
58045 => "0111111111000000",
58046 => "0111111111000000",
58047 => "0111111111000000",
58048 => "0111111111000000",
58049 => "0111111111000000",
58050 => "0111111111000000",
58051 => "0111111111000000",
58052 => "0111111111000000",
58053 => "0111111111000000",
58054 => "0111111111000000",
58055 => "0111111111000000",
58056 => "0111111111000000",
58057 => "0111111111000000",
58058 => "0111111111000000",
58059 => "0111111111000000",
58060 => "0111111111000000",
58061 => "0111111111000000",
58062 => "0111111111000000",
58063 => "0111111111000000",
58064 => "0111111111000000",
58065 => "0111111111000000",
58066 => "0111111111000000",
58067 => "0111111111000000",
58068 => "0111111111000000",
58069 => "0111111111000000",
58070 => "0111111111000000",
58071 => "0111111111000000",
58072 => "0111111111000000",
58073 => "0111111111000000",
58074 => "0111111111000000",
58075 => "0111111111000000",
58076 => "0111111111000000",
58077 => "0111111111000000",
58078 => "0111111111000000",
58079 => "0111111111000000",
58080 => "0111111111000000",
58081 => "0111111111000000",
58082 => "0111111111000000",
58083 => "0111111111000000",
58084 => "0111111111000000",
58085 => "0111111111000000",
58086 => "0111111111000000",
58087 => "0111111111000000",
58088 => "0111111111000000",
58089 => "0111111111000000",
58090 => "0111111111000000",
58091 => "0111111111000000",
58092 => "0111111111000000",
58093 => "0111111111000000",
58094 => "0111111111000000",
58095 => "0111111111000000",
58096 => "0111111111000000",
58097 => "0111111111000000",
58098 => "0111111111000000",
58099 => "0111111111000000",
58100 => "0111111111000000",
58101 => "0111111111000000",
58102 => "0111111111000000",
58103 => "0111111111000000",
58104 => "0111111111000000",
58105 => "0111111111000000",
58106 => "0111111111000000",
58107 => "0111111111000000",
58108 => "0111111111000000",
58109 => "0111111111000000",
58110 => "0111111111000000",
58111 => "0111111111000000",
58112 => "0111111111000000",
58113 => "0111111111000000",
58114 => "0111111111000000",
58115 => "0111111111000000",
58116 => "0111111111000000",
58117 => "0111111111000000",
58118 => "0111111111000000",
58119 => "0111111111000000",
58120 => "0111111111000000",
58121 => "0111111111000000",
58122 => "0111111111000000",
58123 => "0111111111000000",
58124 => "0111111111000000",
58125 => "0111111111000000",
58126 => "0111111111000000",
58127 => "0111111111000000",
58128 => "0111111111000000",
58129 => "0111111111000000",
58130 => "0111111111000000",
58131 => "0111111111000000",
58132 => "0111111111000000",
58133 => "0111111111000000",
58134 => "0111111111000000",
58135 => "0111111111000000",
58136 => "0111111111000000",
58137 => "0111111111000000",
58138 => "0111111111000000",
58139 => "0111111111000000",
58140 => "0111111111000000",
58141 => "0111111111000000",
58142 => "0111111111000000",
58143 => "0111111111000000",
58144 => "0111111111000000",
58145 => "0111111111000000",
58146 => "0111111111000000",
58147 => "0111111111000000",
58148 => "0111111111000000",
58149 => "0111111111000000",
58150 => "0111111111000000",
58151 => "0111111111000000",
58152 => "0111111111000000",
58153 => "0111111111000000",
58154 => "0111111111000000",
58155 => "0111111111000000",
58156 => "0111111111000000",
58157 => "0111111111000000",
58158 => "0111111111000000",
58159 => "0111111111000000",
58160 => "0111111111000000",
58161 => "0111111111000000",
58162 => "0111111111000000",
58163 => "0111111111000000",
58164 => "0111111111000000",
58165 => "0111111111000000",
58166 => "0111111111000000",
58167 => "0111111111000000",
58168 => "0111111111000000",
58169 => "0111111111000000",
58170 => "0111111111000000",
58171 => "0111111111000000",
58172 => "0111111111000000",
58173 => "0111111111000000",
58174 => "0111111111000000",
58175 => "0111111111000000",
58176 => "0111111111000000",
58177 => "0111111111000000",
58178 => "0111111111000000",
58179 => "0111111111000000",
58180 => "0111111111000000",
58181 => "0111111111000000",
58182 => "0111111111000000",
58183 => "0111111111000000",
58184 => "0111111111000000",
58185 => "0111111111000000",
58186 => "0111111111000000",
58187 => "0111111111000000",
58188 => "0111111111000000",
58189 => "0111111111000000",
58190 => "0111111111000000",
58191 => "0111111111000000",
58192 => "0111111111000000",
58193 => "0111111111000000",
58194 => "0111111111000000",
58195 => "0111111111000000",
58196 => "0111111111000000",
58197 => "0111111111000000",
58198 => "0111111111000000",
58199 => "0111111111000000",
58200 => "0111111111000000",
58201 => "0111111111000000",
58202 => "0111111111000000",
58203 => "0111111111000000",
58204 => "0111111111000000",
58205 => "0111111111000000",
58206 => "0111111111000000",
58207 => "0111111111000000",
58208 => "0111111111000000",
58209 => "0111111111000000",
58210 => "0111111111000000",
58211 => "0111111111000000",
58212 => "0111111111000000",
58213 => "0111111111000000",
58214 => "0111111111000000",
58215 => "0111111111000000",
58216 => "0111111111000000",
58217 => "0111111111000000",
58218 => "0111111111000000",
58219 => "0111111111000000",
58220 => "0111111111000000",
58221 => "0111111111000000",
58222 => "0111111111000000",
58223 => "0111111111000000",
58224 => "0111111111000000",
58225 => "0111111111000000",
58226 => "0111111111000000",
58227 => "0111111111000000",
58228 => "0111111111000000",
58229 => "0111111111000000",
58230 => "0111111111000000",
58231 => "0111111111000000",
58232 => "0111111111000000",
58233 => "0111111111000000",
58234 => "0111111111000000",
58235 => "0111111111000000",
58236 => "0111111111000000",
58237 => "0111111111000000",
58238 => "0111111111000000",
58239 => "0111111111000000",
58240 => "0111111111000000",
58241 => "0111111111000000",
58242 => "0111111111000000",
58243 => "0111111111000000",
58244 => "0111111111000000",
58245 => "0111111111000000",
58246 => "0111111111000000",
58247 => "0111111111000000",
58248 => "0111111111000000",
58249 => "0111111111000000",
58250 => "0111111111000000",
58251 => "0111111111000000",
58252 => "0111111111000000",
58253 => "0111111111000000",
58254 => "0111111111000000",
58255 => "0111111111000000",
58256 => "0111111111000000",
58257 => "0111111111000000",
58258 => "0111111111000000",
58259 => "0111111111000000",
58260 => "0111111111000000",
58261 => "0111111111000000",
58262 => "0111111111000000",
58263 => "0111111111000000",
58264 => "0111111111000000",
58265 => "0111111111000000",
58266 => "0111111111000000",
58267 => "0111111111000000",
58268 => "0111111111000000",
58269 => "0111111111000000",
58270 => "0111111111000000",
58271 => "0111111111000000",
58272 => "0111111111000000",
58273 => "0111111111000000",
58274 => "0111111111000000",
58275 => "0111111111000000",
58276 => "0111111111000000",
58277 => "0111111111000000",
58278 => "0111111111000000",
58279 => "0111111111000000",
58280 => "0111111111000000",
58281 => "0111111111000000",
58282 => "0111111111000000",
58283 => "0111111111000000",
58284 => "0111111111000000",
58285 => "0111111111000000",
58286 => "0111111111000000",
58287 => "0111111111000000",
58288 => "0111111111000000",
58289 => "0111111111000000",
58290 => "0111111111000000",
58291 => "0111111111000000",
58292 => "0111111111000000",
58293 => "0111111111000000",
58294 => "0111111111000000",
58295 => "0111111111000000",
58296 => "0111111111000000",
58297 => "0111111111000000",
58298 => "0111111111000000",
58299 => "0111111111000000",
58300 => "0111111111000000",
58301 => "0111111111000000",
58302 => "0111111111000000",
58303 => "0111111111000000",
58304 => "0111111111000000",
58305 => "0111111111000000",
58306 => "0111111111000000",
58307 => "0111111111000000",
58308 => "0111111111000000",
58309 => "0111111111000000",
58310 => "0111111111000000",
58311 => "0111111111000000",
58312 => "0111111111000000",
58313 => "0111111111000000",
58314 => "0111111111000000",
58315 => "0111111111000000",
58316 => "0111111111000000",
58317 => "0111111111000000",
58318 => "0111111111000000",
58319 => "0111111111000000",
58320 => "0111111111000000",
58321 => "0111111111000000",
58322 => "0111111111000000",
58323 => "0111111111000000",
58324 => "0111111111000000",
58325 => "0111111111000000",
58326 => "0111111111000000",
58327 => "0111111111000000",
58328 => "0111111111000000",
58329 => "0111111111000000",
58330 => "0111111111000000",
58331 => "0111111111000000",
58332 => "0111111111000000",
58333 => "0111111111000000",
58334 => "0111111111000000",
58335 => "0111111111000000",
58336 => "0111111111000000",
58337 => "0111111111000000",
58338 => "0111111111000000",
58339 => "0111111111000000",
58340 => "0111111111000000",
58341 => "0111111111000000",
58342 => "0111111111000000",
58343 => "0111111111000000",
58344 => "0111111111000000",
58345 => "0111111111000000",
58346 => "0111111111000000",
58347 => "0111111111000000",
58348 => "0111111111000000",
58349 => "0111111111000000",
58350 => "0111111111000000",
58351 => "0111111111000000",
58352 => "0111111111000000",
58353 => "0111111111000000",
58354 => "0111111111000000",
58355 => "0111111111000000",
58356 => "0111111111000000",
58357 => "0111111111000000",
58358 => "0111111111000000",
58359 => "0111111111000000",
58360 => "0111111111000000",
58361 => "0111111111000000",
58362 => "0111111111000000",
58363 => "0111111111000000",
58364 => "0111111111000000",
58365 => "0111111111000000",
58366 => "0111111111000000",
58367 => "0111111111000000",
58368 => "0111111111000000",
58369 => "0111111111000000",
58370 => "0111111111000000",
58371 => "0111111111000000",
58372 => "0111111111000000",
58373 => "0111111111000000",
58374 => "0111111111000000",
58375 => "0111111111000000",
58376 => "0111111111000000",
58377 => "0111111111000000",
58378 => "0111111111000000",
58379 => "0111111111000000",
58380 => "0111111111000000",
58381 => "0111111111000000",
58382 => "0111111111000000",
58383 => "0111111111000000",
58384 => "0111111111000000",
58385 => "0111111111000000",
58386 => "0111111111000000",
58387 => "0111111111000000",
58388 => "0111111111000000",
58389 => "0111111111000000",
58390 => "0111111111000000",
58391 => "0111111111000000",
58392 => "0111111111000000",
58393 => "0111111111000000",
58394 => "0111111111000000",
58395 => "0111111111000000",
58396 => "0111111111000000",
58397 => "0111111111000000",
58398 => "0111111111000000",
58399 => "0111111111000000",
58400 => "0111111111000000",
58401 => "0111111111000000",
58402 => "0111111111000000",
58403 => "0111111111000000",
58404 => "0111111111000000",
58405 => "0111111111000000",
58406 => "0111111111000000",
58407 => "0111111111000000",
58408 => "0111111111000000",
58409 => "0111111111000000",
58410 => "0111111111000000",
58411 => "0111111111000000",
58412 => "0111111111000000",
58413 => "0111111111000000",
58414 => "0111111111000000",
58415 => "0111111111000000",
58416 => "0111111111000000",
58417 => "0111111111000000",
58418 => "0111111111000000",
58419 => "0111111111000000",
58420 => "0111111111000000",
58421 => "0111111111000000",
58422 => "0111111111000000",
58423 => "0111111111000000",
58424 => "0111111111000000",
58425 => "0111111111000000",
58426 => "0111111111000000",
58427 => "0111111111000000",
58428 => "0111111111000000",
58429 => "0111111111000000",
58430 => "0111111111000000",
58431 => "0111111111000000",
58432 => "0111111111000000",
58433 => "0111111111000000",
58434 => "0111111111000000",
58435 => "0111111111000000",
58436 => "0111111111000000",
58437 => "0111111111000000",
58438 => "0111111111000000",
58439 => "0111111111000000",
58440 => "0111111111000000",
58441 => "0111111111000000",
58442 => "0111111111000000",
58443 => "0111111111000000",
58444 => "0111111111000000",
58445 => "0111111111000000",
58446 => "0111111111000000",
58447 => "0111111111000000",
58448 => "0111111111000000",
58449 => "0111111111000000",
58450 => "0111111111000000",
58451 => "0111111111000000",
58452 => "0111111111000000",
58453 => "0111111111000000",
58454 => "0111111111000000",
58455 => "0111111111000000",
58456 => "0111111111000000",
58457 => "0111111111000000",
58458 => "0111111111000000",
58459 => "0111111111000000",
58460 => "0111111111000000",
58461 => "0111111111000000",
58462 => "0111111111000000",
58463 => "0111111111000000",
58464 => "0111111111000000",
58465 => "0111111111000000",
58466 => "0111111111000000",
58467 => "0111111111000000",
58468 => "0111111111000000",
58469 => "0111111111000000",
58470 => "0111111111000000",
58471 => "0111111111000000",
58472 => "0111111111000000",
58473 => "0111111111000000",
58474 => "0111111111000000",
58475 => "0111111111000000",
58476 => "0111111111000000",
58477 => "0111111111000000",
58478 => "0111111111000000",
58479 => "0111111111000000",
58480 => "0111111111000000",
58481 => "0111111111000000",
58482 => "0111111111000000",
58483 => "0111111111000000",
58484 => "0111111111000000",
58485 => "0111111111000000",
58486 => "0111111111000000",
58487 => "0111111111000000",
58488 => "0111111111000000",
58489 => "0111111111000000",
58490 => "0111111111000000",
58491 => "0111111111000000",
58492 => "0111111111000000",
58493 => "0111111111000000",
58494 => "0111111111000000",
58495 => "0111111111000000",
58496 => "0111111111000000",
58497 => "0111111111000000",
58498 => "0111111111000000",
58499 => "0111111111000000",
58500 => "0111111111000000",
58501 => "0111111111000000",
58502 => "0111111111000000",
58503 => "0111111111000000",
58504 => "0111111111000000",
58505 => "0111111111000000",
58506 => "0111111111000000",
58507 => "0111111111000000",
58508 => "0111111111000000",
58509 => "0111111111000000",
58510 => "0111111111000000",
58511 => "0111111111000000",
58512 => "0111111111000000",
58513 => "0111111111000000",
58514 => "0111111111000000",
58515 => "0111111111000000",
58516 => "0111111111000000",
58517 => "0111111111000000",
58518 => "0111111111000000",
58519 => "0111111111000000",
58520 => "0111111111000000",
58521 => "0111111111000000",
58522 => "0111111111000000",
58523 => "0111111111000000",
58524 => "0111111111000000",
58525 => "0111111111000000",
58526 => "0111111111000000",
58527 => "0111111111000000",
58528 => "0111111111000000",
58529 => "0111111111000000",
58530 => "0111111111000000",
58531 => "0111111111000000",
58532 => "0111111111000000",
58533 => "0111111111000000",
58534 => "0111111111000000",
58535 => "0111111111000000",
58536 => "0111111111000000",
58537 => "0111111111000000",
58538 => "0111111111000000",
58539 => "0111111111000000",
58540 => "0111111111000000",
58541 => "0111111111000000",
58542 => "0111111111000000",
58543 => "0111111111000000",
58544 => "0111111111000000",
58545 => "0111111111000000",
58546 => "0111111111000000",
58547 => "0111111111000000",
58548 => "0111111111000000",
58549 => "0111111111000000",
58550 => "0111111111000000",
58551 => "0111111111000000",
58552 => "0111111111000000",
58553 => "0111111111000000",
58554 => "0111111111000000",
58555 => "0111111111000000",
58556 => "0111111111000000",
58557 => "0111111111000000",
58558 => "0111111111000000",
58559 => "0111111111000000",
58560 => "0111111111000000",
58561 => "0111111111000000",
58562 => "0111111111000000",
58563 => "0111111111000000",
58564 => "0111111111000000",
58565 => "0111111111000000",
58566 => "0111111111000000",
58567 => "0111111111000000",
58568 => "0111111111000000",
58569 => "0111111111000000",
58570 => "0111111111000000",
58571 => "0111111111000000",
58572 => "0111111111000000",
58573 => "0111111111000000",
58574 => "0111111111000000",
58575 => "0111111111000000",
58576 => "0111111111000000",
58577 => "0111111111000000",
58578 => "0111111111000000",
58579 => "0111111111000000",
58580 => "0111111111000000",
58581 => "0111111111000000",
58582 => "0111111111000000",
58583 => "0111111111000000",
58584 => "0111111111000000",
58585 => "0111111111000000",
58586 => "0111111111000000",
58587 => "0111111111000000",
58588 => "0111111111000000",
58589 => "0111111111000000",
58590 => "0111111111000000",
58591 => "0111111111000000",
58592 => "0111111111000000",
58593 => "0111111111000000",
58594 => "0111111111000000",
58595 => "0111111111000000",
58596 => "0111111111000000",
58597 => "0111111111000000",
58598 => "0111111111000000",
58599 => "0111111111000000",
58600 => "0111111111000000",
58601 => "0111111111000000",
58602 => "0111111111000000",
58603 => "0111111111000000",
58604 => "0111111111000000",
58605 => "0111111111000000",
58606 => "0111111111000000",
58607 => "0111111111000000",
58608 => "0111111111000000",
58609 => "0111111111000000",
58610 => "0111111111000000",
58611 => "0111111111000000",
58612 => "0111111111000000",
58613 => "0111111111000000",
58614 => "0111111111000000",
58615 => "0111111111000000",
58616 => "0111111111000000",
58617 => "0111111111000000",
58618 => "0111111111000000",
58619 => "0111111111000000",
58620 => "0111111111000000",
58621 => "0111111111000000",
58622 => "0111111111000000",
58623 => "0111111111000000",
58624 => "0111111111000000",
58625 => "0111111111000000",
58626 => "0111111111000000",
58627 => "0111111111000000",
58628 => "0111111111000000",
58629 => "0111111111000000",
58630 => "0111111111000000",
58631 => "0111111111000000",
58632 => "0111111111000000",
58633 => "0111111111000000",
58634 => "0111111111000000",
58635 => "0111111111000000",
58636 => "0111111111000000",
58637 => "0111111111000000",
58638 => "0111111111000000",
58639 => "0111111111000000",
58640 => "0111111111000000",
58641 => "0111111111000000",
58642 => "0111111111000000",
58643 => "0111111111000000",
58644 => "0111111111000000",
58645 => "0111111111000000",
58646 => "0111111111000000",
58647 => "0111111111000000",
58648 => "0111111111000000",
58649 => "0111111111000000",
58650 => "0111111111000000",
58651 => "0111111111000000",
58652 => "0111111111000000",
58653 => "0111111111000000",
58654 => "0111111111000000",
58655 => "0111111111000000",
58656 => "0111111111000000",
58657 => "0111111111000000",
58658 => "0111111111000000",
58659 => "0111111111000000",
58660 => "0111111111000000",
58661 => "0111111111000000",
58662 => "0111111111000000",
58663 => "0111111111000000",
58664 => "0111111111000000",
58665 => "0111111111000000",
58666 => "0111111111000000",
58667 => "0111111111000000",
58668 => "0111111111000000",
58669 => "0111111111000000",
58670 => "0111111111000000",
58671 => "0111111111000000",
58672 => "0111111111000000",
58673 => "0111111111000000",
58674 => "0111111111000000",
58675 => "0111111111000000",
58676 => "0111111111000000",
58677 => "0111111111000000",
58678 => "0111111111000000",
58679 => "0111111111000000",
58680 => "0111111111000000",
58681 => "0111111111000000",
58682 => "0111111111000000",
58683 => "0111111111000000",
58684 => "0111111111000000",
58685 => "0111111111000000",
58686 => "0111111111000000",
58687 => "0111111111000000",
58688 => "0111111111000000",
58689 => "0111111111000000",
58690 => "0111111111000000",
58691 => "0111111111000000",
58692 => "0111111111000000",
58693 => "0111111111000000",
58694 => "0111111111000000",
58695 => "0111111111000000",
58696 => "0111111111000000",
58697 => "0111111111000000",
58698 => "0111111111000000",
58699 => "0111111111000000",
58700 => "0111111111000000",
58701 => "0111111111000000",
58702 => "0111111111000000",
58703 => "0111111111000000",
58704 => "0111111111000000",
58705 => "0111111111000000",
58706 => "0111111111000000",
58707 => "0111111111000000",
58708 => "0111111111000000",
58709 => "0111111111000000",
58710 => "0111111111000000",
58711 => "0111111111000000",
58712 => "0111111111000000",
58713 => "0111111111000000",
58714 => "0111111111000000",
58715 => "0111111111000000",
58716 => "0111111111000000",
58717 => "0111111111000000",
58718 => "0111111111000000",
58719 => "0111111111000000",
58720 => "0111111111000000",
58721 => "0111111111000000",
58722 => "0111111111000000",
58723 => "0111111111000000",
58724 => "0111111111000000",
58725 => "0111111111000000",
58726 => "0111111111000000",
58727 => "0111111111000000",
58728 => "0111111111000000",
58729 => "0111111111000000",
58730 => "0111111111000000",
58731 => "0111111111000000",
58732 => "0111111111000000",
58733 => "0111111111000000",
58734 => "0111111111000000",
58735 => "0111111111000000",
58736 => "0111111111000000",
58737 => "0111111111000000",
58738 => "0111111111000000",
58739 => "0111111111000000",
58740 => "0111111111000000",
58741 => "0111111111000000",
58742 => "0111111111000000",
58743 => "0111111111000000",
58744 => "0111111111000000",
58745 => "0111111111000000",
58746 => "0111111111000000",
58747 => "0111111111000000",
58748 => "0111111111000000",
58749 => "0111111111000000",
58750 => "0111111111000000",
58751 => "0111111111000000",
58752 => "0111111111000000",
58753 => "0111111111000000",
58754 => "0111111111000000",
58755 => "0111111111000000",
58756 => "0111111111000000",
58757 => "0111111111000000",
58758 => "0111111111000000",
58759 => "0111111111000000",
58760 => "0111111111000000",
58761 => "0111111111000000",
58762 => "0111111111000000",
58763 => "0111111111000000",
58764 => "0111111111000000",
58765 => "0111111111000000",
58766 => "0111111111000000",
58767 => "0111111111000000",
58768 => "0111111111000000",
58769 => "0111111111000000",
58770 => "0111111111000000",
58771 => "0111111111000000",
58772 => "0111111111000000",
58773 => "0111111111000000",
58774 => "0111111111000000",
58775 => "0111111111000000",
58776 => "0111111111000000",
58777 => "0111111111000000",
58778 => "0111111111000000",
58779 => "0111111111000000",
58780 => "0111111111000000",
58781 => "0111111111000000",
58782 => "0111111111000000",
58783 => "0111111111000000",
58784 => "0111111111000000",
58785 => "0111111111000000",
58786 => "0111111111000000",
58787 => "0111111111000000",
58788 => "0111111111000000",
58789 => "0111111111000000",
58790 => "0111111111000000",
58791 => "0111111111000000",
58792 => "0111111111000000",
58793 => "0111111111000000",
58794 => "0111111111000000",
58795 => "0111111111000000",
58796 => "0111111111000000",
58797 => "0111111111000000",
58798 => "0111111111000000",
58799 => "0111111111000000",
58800 => "0111111111000000",
58801 => "0111111111000000",
58802 => "0111111111000000",
58803 => "0111111111000000",
58804 => "0111111111000000",
58805 => "0111111111000000",
58806 => "0111111111000000",
58807 => "0111111111000000",
58808 => "0111111111000000",
58809 => "0111111111000000",
58810 => "0111111111000000",
58811 => "0111111111000000",
58812 => "0111111111000000",
58813 => "0111111111000000",
58814 => "0111111111000000",
58815 => "0111111111000000",
58816 => "0111111111000000",
58817 => "0111111111000000",
58818 => "0111111111000000",
58819 => "0111111111000000",
58820 => "0111111111000000",
58821 => "0111111111000000",
58822 => "0111111111000000",
58823 => "0111111111000000",
58824 => "0111111111000000",
58825 => "0111111111000000",
58826 => "0111111111000000",
58827 => "0111111111000000",
58828 => "0111111111000000",
58829 => "0111111111000000",
58830 => "0111111111000000",
58831 => "0111111111000000",
58832 => "0111111111000000",
58833 => "0111111111000000",
58834 => "0111111111000000",
58835 => "0111111111000000",
58836 => "0111111111000000",
58837 => "0111111111000000",
58838 => "0111111111000000",
58839 => "0111111111000000",
58840 => "0111111111000000",
58841 => "0111111111000000",
58842 => "0111111111000000",
58843 => "0111111111000000",
58844 => "0111111111000000",
58845 => "0111111111000000",
58846 => "0111111111000000",
58847 => "0111111111000000",
58848 => "0111111111000000",
58849 => "0111111111000000",
58850 => "0111111111000000",
58851 => "0111111111000000",
58852 => "0111111111000000",
58853 => "0111111111000000",
58854 => "0111111111000000",
58855 => "0111111111000000",
58856 => "0111111111000000",
58857 => "0111111111000000",
58858 => "0111111111000000",
58859 => "0111111111000000",
58860 => "0111111111010000",
58861 => "0111111111010000",
58862 => "0111111111010000",
58863 => "0111111111010000",
58864 => "0111111111010000",
58865 => "0111111111010000",
58866 => "0111111111010000",
58867 => "0111111111010000",
58868 => "0111111111010000",
58869 => "0111111111010000",
58870 => "0111111111010000",
58871 => "0111111111010000",
58872 => "0111111111010000",
58873 => "0111111111010000",
58874 => "0111111111010000",
58875 => "0111111111010000",
58876 => "0111111111010000",
58877 => "0111111111010000",
58878 => "0111111111010000",
58879 => "0111111111010000",
58880 => "0111111111010000",
58881 => "0111111111010000",
58882 => "0111111111010000",
58883 => "0111111111010000",
58884 => "0111111111010000",
58885 => "0111111111010000",
58886 => "0111111111010000",
58887 => "0111111111010000",
58888 => "0111111111010000",
58889 => "0111111111010000",
58890 => "0111111111010000",
58891 => "0111111111010000",
58892 => "0111111111010000",
58893 => "0111111111010000",
58894 => "0111111111010000",
58895 => "0111111111010000",
58896 => "0111111111010000",
58897 => "0111111111010000",
58898 => "0111111111010000",
58899 => "0111111111010000",
58900 => "0111111111010000",
58901 => "0111111111010000",
58902 => "0111111111010000",
58903 => "0111111111010000",
58904 => "0111111111010000",
58905 => "0111111111010000",
58906 => "0111111111010000",
58907 => "0111111111010000",
58908 => "0111111111010000",
58909 => "0111111111010000",
58910 => "0111111111010000",
58911 => "0111111111010000",
58912 => "0111111111010000",
58913 => "0111111111010000",
58914 => "0111111111010000",
58915 => "0111111111010000",
58916 => "0111111111010000",
58917 => "0111111111010000",
58918 => "0111111111010000",
58919 => "0111111111010000",
58920 => "0111111111010000",
58921 => "0111111111010000",
58922 => "0111111111010000",
58923 => "0111111111010000",
58924 => "0111111111010000",
58925 => "0111111111010000",
58926 => "0111111111010000",
58927 => "0111111111010000",
58928 => "0111111111010000",
58929 => "0111111111010000",
58930 => "0111111111010000",
58931 => "0111111111010000",
58932 => "0111111111010000",
58933 => "0111111111010000",
58934 => "0111111111010000",
58935 => "0111111111010000",
58936 => "0111111111010000",
58937 => "0111111111010000",
58938 => "0111111111010000",
58939 => "0111111111010000",
58940 => "0111111111010000",
58941 => "0111111111010000",
58942 => "0111111111010000",
58943 => "0111111111010000",
58944 => "0111111111010000",
58945 => "0111111111010000",
58946 => "0111111111010000",
58947 => "0111111111010000",
58948 => "0111111111010000",
58949 => "0111111111010000",
58950 => "0111111111010000",
58951 => "0111111111010000",
58952 => "0111111111010000",
58953 => "0111111111010000",
58954 => "0111111111010000",
58955 => "0111111111010000",
58956 => "0111111111010000",
58957 => "0111111111010000",
58958 => "0111111111010000",
58959 => "0111111111010000",
58960 => "0111111111010000",
58961 => "0111111111010000",
58962 => "0111111111010000",
58963 => "0111111111010000",
58964 => "0111111111010000",
58965 => "0111111111010000",
58966 => "0111111111010000",
58967 => "0111111111010000",
58968 => "0111111111010000",
58969 => "0111111111010000",
58970 => "0111111111010000",
58971 => "0111111111010000",
58972 => "0111111111010000",
58973 => "0111111111010000",
58974 => "0111111111010000",
58975 => "0111111111010000",
58976 => "0111111111010000",
58977 => "0111111111010000",
58978 => "0111111111010000",
58979 => "0111111111010000",
58980 => "0111111111010000",
58981 => "0111111111010000",
58982 => "0111111111010000",
58983 => "0111111111010000",
58984 => "0111111111010000",
58985 => "0111111111010000",
58986 => "0111111111010000",
58987 => "0111111111010000",
58988 => "0111111111010000",
58989 => "0111111111010000",
58990 => "0111111111010000",
58991 => "0111111111010000",
58992 => "0111111111010000",
58993 => "0111111111010000",
58994 => "0111111111010000",
58995 => "0111111111010000",
58996 => "0111111111010000",
58997 => "0111111111010000",
58998 => "0111111111010000",
58999 => "0111111111010000",
59000 => "0111111111010000",
59001 => "0111111111010000",
59002 => "0111111111010000",
59003 => "0111111111010000",
59004 => "0111111111010000",
59005 => "0111111111010000",
59006 => "0111111111010000",
59007 => "0111111111010000",
59008 => "0111111111010000",
59009 => "0111111111010000",
59010 => "0111111111010000",
59011 => "0111111111010000",
59012 => "0111111111010000",
59013 => "0111111111010000",
59014 => "0111111111010000",
59015 => "0111111111010000",
59016 => "0111111111010000",
59017 => "0111111111010000",
59018 => "0111111111010000",
59019 => "0111111111010000",
59020 => "0111111111010000",
59021 => "0111111111010000",
59022 => "0111111111010000",
59023 => "0111111111010000",
59024 => "0111111111010000",
59025 => "0111111111010000",
59026 => "0111111111010000",
59027 => "0111111111010000",
59028 => "0111111111010000",
59029 => "0111111111010000",
59030 => "0111111111010000",
59031 => "0111111111010000",
59032 => "0111111111010000",
59033 => "0111111111010000",
59034 => "0111111111010000",
59035 => "0111111111010000",
59036 => "0111111111010000",
59037 => "0111111111010000",
59038 => "0111111111010000",
59039 => "0111111111010000",
59040 => "0111111111010000",
59041 => "0111111111010000",
59042 => "0111111111010000",
59043 => "0111111111010000",
59044 => "0111111111010000",
59045 => "0111111111010000",
59046 => "0111111111010000",
59047 => "0111111111010000",
59048 => "0111111111010000",
59049 => "0111111111010000",
59050 => "0111111111010000",
59051 => "0111111111010000",
59052 => "0111111111010000",
59053 => "0111111111010000",
59054 => "0111111111010000",
59055 => "0111111111010000",
59056 => "0111111111010000",
59057 => "0111111111010000",
59058 => "0111111111010000",
59059 => "0111111111010000",
59060 => "0111111111010000",
59061 => "0111111111010000",
59062 => "0111111111010000",
59063 => "0111111111010000",
59064 => "0111111111010000",
59065 => "0111111111010000",
59066 => "0111111111010000",
59067 => "0111111111010000",
59068 => "0111111111010000",
59069 => "0111111111010000",
59070 => "0111111111010000",
59071 => "0111111111010000",
59072 => "0111111111010000",
59073 => "0111111111010000",
59074 => "0111111111010000",
59075 => "0111111111010000",
59076 => "0111111111010000",
59077 => "0111111111010000",
59078 => "0111111111010000",
59079 => "0111111111010000",
59080 => "0111111111010000",
59081 => "0111111111010000",
59082 => "0111111111010000",
59083 => "0111111111010000",
59084 => "0111111111010000",
59085 => "0111111111010000",
59086 => "0111111111010000",
59087 => "0111111111010000",
59088 => "0111111111010000",
59089 => "0111111111010000",
59090 => "0111111111010000",
59091 => "0111111111010000",
59092 => "0111111111010000",
59093 => "0111111111010000",
59094 => "0111111111010000",
59095 => "0111111111010000",
59096 => "0111111111010000",
59097 => "0111111111010000",
59098 => "0111111111010000",
59099 => "0111111111010000",
59100 => "0111111111010000",
59101 => "0111111111010000",
59102 => "0111111111010000",
59103 => "0111111111010000",
59104 => "0111111111010000",
59105 => "0111111111010000",
59106 => "0111111111010000",
59107 => "0111111111010000",
59108 => "0111111111010000",
59109 => "0111111111010000",
59110 => "0111111111010000",
59111 => "0111111111010000",
59112 => "0111111111010000",
59113 => "0111111111010000",
59114 => "0111111111010000",
59115 => "0111111111010000",
59116 => "0111111111010000",
59117 => "0111111111010000",
59118 => "0111111111010000",
59119 => "0111111111010000",
59120 => "0111111111010000",
59121 => "0111111111010000",
59122 => "0111111111010000",
59123 => "0111111111010000",
59124 => "0111111111010000",
59125 => "0111111111010000",
59126 => "0111111111010000",
59127 => "0111111111010000",
59128 => "0111111111010000",
59129 => "0111111111010000",
59130 => "0111111111010000",
59131 => "0111111111010000",
59132 => "0111111111010000",
59133 => "0111111111010000",
59134 => "0111111111010000",
59135 => "0111111111010000",
59136 => "0111111111010000",
59137 => "0111111111010000",
59138 => "0111111111010000",
59139 => "0111111111010000",
59140 => "0111111111010000",
59141 => "0111111111010000",
59142 => "0111111111010000",
59143 => "0111111111010000",
59144 => "0111111111010000",
59145 => "0111111111010000",
59146 => "0111111111010000",
59147 => "0111111111010000",
59148 => "0111111111010000",
59149 => "0111111111010000",
59150 => "0111111111010000",
59151 => "0111111111010000",
59152 => "0111111111010000",
59153 => "0111111111010000",
59154 => "0111111111010000",
59155 => "0111111111010000",
59156 => "0111111111010000",
59157 => "0111111111010000",
59158 => "0111111111010000",
59159 => "0111111111010000",
59160 => "0111111111010000",
59161 => "0111111111010000",
59162 => "0111111111010000",
59163 => "0111111111010000",
59164 => "0111111111010000",
59165 => "0111111111010000",
59166 => "0111111111010000",
59167 => "0111111111010000",
59168 => "0111111111010000",
59169 => "0111111111010000",
59170 => "0111111111010000",
59171 => "0111111111010000",
59172 => "0111111111010000",
59173 => "0111111111010000",
59174 => "0111111111010000",
59175 => "0111111111010000",
59176 => "0111111111010000",
59177 => "0111111111010000",
59178 => "0111111111010000",
59179 => "0111111111010000",
59180 => "0111111111010000",
59181 => "0111111111010000",
59182 => "0111111111010000",
59183 => "0111111111010000",
59184 => "0111111111010000",
59185 => "0111111111010000",
59186 => "0111111111010000",
59187 => "0111111111010000",
59188 => "0111111111010000",
59189 => "0111111111010000",
59190 => "0111111111010000",
59191 => "0111111111010000",
59192 => "0111111111010000",
59193 => "0111111111010000",
59194 => "0111111111010000",
59195 => "0111111111010000",
59196 => "0111111111010000",
59197 => "0111111111010000",
59198 => "0111111111010000",
59199 => "0111111111010000",
59200 => "0111111111010000",
59201 => "0111111111010000",
59202 => "0111111111010000",
59203 => "0111111111010000",
59204 => "0111111111010000",
59205 => "0111111111010000",
59206 => "0111111111010000",
59207 => "0111111111010000",
59208 => "0111111111010000",
59209 => "0111111111010000",
59210 => "0111111111010000",
59211 => "0111111111010000",
59212 => "0111111111010000",
59213 => "0111111111010000",
59214 => "0111111111010000",
59215 => "0111111111010000",
59216 => "0111111111010000",
59217 => "0111111111010000",
59218 => "0111111111010000",
59219 => "0111111111010000",
59220 => "0111111111010000",
59221 => "0111111111010000",
59222 => "0111111111010000",
59223 => "0111111111010000",
59224 => "0111111111010000",
59225 => "0111111111010000",
59226 => "0111111111010000",
59227 => "0111111111010000",
59228 => "0111111111010000",
59229 => "0111111111010000",
59230 => "0111111111010000",
59231 => "0111111111010000",
59232 => "0111111111010000",
59233 => "0111111111010000",
59234 => "0111111111010000",
59235 => "0111111111010000",
59236 => "0111111111010000",
59237 => "0111111111010000",
59238 => "0111111111010000",
59239 => "0111111111010000",
59240 => "0111111111010000",
59241 => "0111111111010000",
59242 => "0111111111010000",
59243 => "0111111111010000",
59244 => "0111111111010000",
59245 => "0111111111010000",
59246 => "0111111111010000",
59247 => "0111111111010000",
59248 => "0111111111010000",
59249 => "0111111111010000",
59250 => "0111111111010000",
59251 => "0111111111010000",
59252 => "0111111111010000",
59253 => "0111111111010000",
59254 => "0111111111010000",
59255 => "0111111111010000",
59256 => "0111111111010000",
59257 => "0111111111010000",
59258 => "0111111111010000",
59259 => "0111111111010000",
59260 => "0111111111010000",
59261 => "0111111111010000",
59262 => "0111111111010000",
59263 => "0111111111010000",
59264 => "0111111111010000",
59265 => "0111111111010000",
59266 => "0111111111010000",
59267 => "0111111111010000",
59268 => "0111111111010000",
59269 => "0111111111010000",
59270 => "0111111111010000",
59271 => "0111111111010000",
59272 => "0111111111010000",
59273 => "0111111111010000",
59274 => "0111111111010000",
59275 => "0111111111010000",
59276 => "0111111111010000",
59277 => "0111111111010000",
59278 => "0111111111010000",
59279 => "0111111111010000",
59280 => "0111111111010000",
59281 => "0111111111010000",
59282 => "0111111111010000",
59283 => "0111111111010000",
59284 => "0111111111010000",
59285 => "0111111111010000",
59286 => "0111111111010000",
59287 => "0111111111010000",
59288 => "0111111111010000",
59289 => "0111111111010000",
59290 => "0111111111010000",
59291 => "0111111111010000",
59292 => "0111111111010000",
59293 => "0111111111010000",
59294 => "0111111111010000",
59295 => "0111111111010000",
59296 => "0111111111010000",
59297 => "0111111111010000",
59298 => "0111111111010000",
59299 => "0111111111010000",
59300 => "0111111111010000",
59301 => "0111111111010000",
59302 => "0111111111010000",
59303 => "0111111111010000",
59304 => "0111111111010000",
59305 => "0111111111010000",
59306 => "0111111111010000",
59307 => "0111111111010000",
59308 => "0111111111010000",
59309 => "0111111111010000",
59310 => "0111111111010000",
59311 => "0111111111010000",
59312 => "0111111111010000",
59313 => "0111111111010000",
59314 => "0111111111010000",
59315 => "0111111111010000",
59316 => "0111111111010000",
59317 => "0111111111010000",
59318 => "0111111111010000",
59319 => "0111111111010000",
59320 => "0111111111010000",
59321 => "0111111111010000",
59322 => "0111111111010000",
59323 => "0111111111010000",
59324 => "0111111111010000",
59325 => "0111111111010000",
59326 => "0111111111010000",
59327 => "0111111111010000",
59328 => "0111111111010000",
59329 => "0111111111010000",
59330 => "0111111111010000",
59331 => "0111111111010000",
59332 => "0111111111010000",
59333 => "0111111111010000",
59334 => "0111111111010000",
59335 => "0111111111010000",
59336 => "0111111111010000",
59337 => "0111111111010000",
59338 => "0111111111010000",
59339 => "0111111111010000",
59340 => "0111111111010000",
59341 => "0111111111010000",
59342 => "0111111111010000",
59343 => "0111111111010000",
59344 => "0111111111010000",
59345 => "0111111111010000",
59346 => "0111111111010000",
59347 => "0111111111010000",
59348 => "0111111111010000",
59349 => "0111111111010000",
59350 => "0111111111010000",
59351 => "0111111111010000",
59352 => "0111111111010000",
59353 => "0111111111010000",
59354 => "0111111111010000",
59355 => "0111111111010000",
59356 => "0111111111010000",
59357 => "0111111111010000",
59358 => "0111111111010000",
59359 => "0111111111010000",
59360 => "0111111111010000",
59361 => "0111111111010000",
59362 => "0111111111010000",
59363 => "0111111111010000",
59364 => "0111111111010000",
59365 => "0111111111010000",
59366 => "0111111111010000",
59367 => "0111111111010000",
59368 => "0111111111010000",
59369 => "0111111111010000",
59370 => "0111111111010000",
59371 => "0111111111010000",
59372 => "0111111111010000",
59373 => "0111111111010000",
59374 => "0111111111010000",
59375 => "0111111111010000",
59376 => "0111111111010000",
59377 => "0111111111010000",
59378 => "0111111111010000",
59379 => "0111111111010000",
59380 => "0111111111010000",
59381 => "0111111111010000",
59382 => "0111111111010000",
59383 => "0111111111010000",
59384 => "0111111111010000",
59385 => "0111111111010000",
59386 => "0111111111010000",
59387 => "0111111111010000",
59388 => "0111111111010000",
59389 => "0111111111010000",
59390 => "0111111111010000",
59391 => "0111111111010000",
59392 => "0111111111010000",
59393 => "0111111111010000",
59394 => "0111111111010000",
59395 => "0111111111010000",
59396 => "0111111111010000",
59397 => "0111111111010000",
59398 => "0111111111010000",
59399 => "0111111111010000",
59400 => "0111111111010000",
59401 => "0111111111010000",
59402 => "0111111111010000",
59403 => "0111111111010000",
59404 => "0111111111010000",
59405 => "0111111111010000",
59406 => "0111111111010000",
59407 => "0111111111010000",
59408 => "0111111111010000",
59409 => "0111111111010000",
59410 => "0111111111010000",
59411 => "0111111111010000",
59412 => "0111111111010000",
59413 => "0111111111010000",
59414 => "0111111111010000",
59415 => "0111111111010000",
59416 => "0111111111010000",
59417 => "0111111111010000",
59418 => "0111111111010000",
59419 => "0111111111010000",
59420 => "0111111111010000",
59421 => "0111111111010000",
59422 => "0111111111010000",
59423 => "0111111111010000",
59424 => "0111111111010000",
59425 => "0111111111010000",
59426 => "0111111111010000",
59427 => "0111111111010000",
59428 => "0111111111010000",
59429 => "0111111111010000",
59430 => "0111111111010000",
59431 => "0111111111010000",
59432 => "0111111111010000",
59433 => "0111111111010000",
59434 => "0111111111010000",
59435 => "0111111111010000",
59436 => "0111111111010000",
59437 => "0111111111010000",
59438 => "0111111111010000",
59439 => "0111111111010000",
59440 => "0111111111010000",
59441 => "0111111111010000",
59442 => "0111111111010000",
59443 => "0111111111010000",
59444 => "0111111111010000",
59445 => "0111111111010000",
59446 => "0111111111010000",
59447 => "0111111111010000",
59448 => "0111111111010000",
59449 => "0111111111010000",
59450 => "0111111111010000",
59451 => "0111111111010000",
59452 => "0111111111010000",
59453 => "0111111111010000",
59454 => "0111111111010000",
59455 => "0111111111010000",
59456 => "0111111111010000",
59457 => "0111111111010000",
59458 => "0111111111010000",
59459 => "0111111111010000",
59460 => "0111111111010000",
59461 => "0111111111010000",
59462 => "0111111111010000",
59463 => "0111111111010000",
59464 => "0111111111010000",
59465 => "0111111111010000",
59466 => "0111111111010000",
59467 => "0111111111010000",
59468 => "0111111111010000",
59469 => "0111111111010000",
59470 => "0111111111010000",
59471 => "0111111111010000",
59472 => "0111111111010000",
59473 => "0111111111010000",
59474 => "0111111111010000",
59475 => "0111111111010000",
59476 => "0111111111010000",
59477 => "0111111111010000",
59478 => "0111111111010000",
59479 => "0111111111010000",
59480 => "0111111111010000",
59481 => "0111111111010000",
59482 => "0111111111010000",
59483 => "0111111111010000",
59484 => "0111111111010000",
59485 => "0111111111010000",
59486 => "0111111111010000",
59487 => "0111111111010000",
59488 => "0111111111010000",
59489 => "0111111111010000",
59490 => "0111111111010000",
59491 => "0111111111010000",
59492 => "0111111111010000",
59493 => "0111111111010000",
59494 => "0111111111010000",
59495 => "0111111111010000",
59496 => "0111111111010000",
59497 => "0111111111010000",
59498 => "0111111111010000",
59499 => "0111111111010000",
59500 => "0111111111010000",
59501 => "0111111111010000",
59502 => "0111111111010000",
59503 => "0111111111010000",
59504 => "0111111111010000",
59505 => "0111111111010000",
59506 => "0111111111010000",
59507 => "0111111111010000",
59508 => "0111111111010000",
59509 => "0111111111010000",
59510 => "0111111111010000",
59511 => "0111111111010000",
59512 => "0111111111010000",
59513 => "0111111111010000",
59514 => "0111111111010000",
59515 => "0111111111010000",
59516 => "0111111111010000",
59517 => "0111111111010000",
59518 => "0111111111010000",
59519 => "0111111111010000",
59520 => "0111111111010000",
59521 => "0111111111010000",
59522 => "0111111111010000",
59523 => "0111111111010000",
59524 => "0111111111010000",
59525 => "0111111111010000",
59526 => "0111111111010000",
59527 => "0111111111010000",
59528 => "0111111111010000",
59529 => "0111111111010000",
59530 => "0111111111010000",
59531 => "0111111111010000",
59532 => "0111111111010000",
59533 => "0111111111010000",
59534 => "0111111111010000",
59535 => "0111111111010000",
59536 => "0111111111010000",
59537 => "0111111111010000",
59538 => "0111111111010000",
59539 => "0111111111010000",
59540 => "0111111111010000",
59541 => "0111111111010000",
59542 => "0111111111010000",
59543 => "0111111111010000",
59544 => "0111111111010000",
59545 => "0111111111010000",
59546 => "0111111111010000",
59547 => "0111111111010000",
59548 => "0111111111010000",
59549 => "0111111111010000",
59550 => "0111111111010000",
59551 => "0111111111010000",
59552 => "0111111111010000",
59553 => "0111111111010000",
59554 => "0111111111010000",
59555 => "0111111111010000",
59556 => "0111111111010000",
59557 => "0111111111010000",
59558 => "0111111111010000",
59559 => "0111111111010000",
59560 => "0111111111010000",
59561 => "0111111111010000",
59562 => "0111111111010000",
59563 => "0111111111010000",
59564 => "0111111111010000",
59565 => "0111111111010000",
59566 => "0111111111010000",
59567 => "0111111111010000",
59568 => "0111111111010000",
59569 => "0111111111010000",
59570 => "0111111111010000",
59571 => "0111111111010000",
59572 => "0111111111010000",
59573 => "0111111111010000",
59574 => "0111111111010000",
59575 => "0111111111010000",
59576 => "0111111111010000",
59577 => "0111111111010000",
59578 => "0111111111010000",
59579 => "0111111111010000",
59580 => "0111111111010000",
59581 => "0111111111010000",
59582 => "0111111111010000",
59583 => "0111111111010000",
59584 => "0111111111010000",
59585 => "0111111111010000",
59586 => "0111111111010000",
59587 => "0111111111010000",
59588 => "0111111111010000",
59589 => "0111111111010000",
59590 => "0111111111010000",
59591 => "0111111111010000",
59592 => "0111111111010000",
59593 => "0111111111010000",
59594 => "0111111111010000",
59595 => "0111111111010000",
59596 => "0111111111010000",
59597 => "0111111111010000",
59598 => "0111111111010000",
59599 => "0111111111010000",
59600 => "0111111111010000",
59601 => "0111111111010000",
59602 => "0111111111010000",
59603 => "0111111111010000",
59604 => "0111111111010000",
59605 => "0111111111010000",
59606 => "0111111111010000",
59607 => "0111111111010000",
59608 => "0111111111010000",
59609 => "0111111111010000",
59610 => "0111111111010000",
59611 => "0111111111010000",
59612 => "0111111111010000",
59613 => "0111111111010000",
59614 => "0111111111010000",
59615 => "0111111111010000",
59616 => "0111111111010000",
59617 => "0111111111010000",
59618 => "0111111111010000",
59619 => "0111111111010000",
59620 => "0111111111010000",
59621 => "0111111111010000",
59622 => "0111111111010000",
59623 => "0111111111010000",
59624 => "0111111111010000",
59625 => "0111111111010000",
59626 => "0111111111010000",
59627 => "0111111111010000",
59628 => "0111111111010000",
59629 => "0111111111010000",
59630 => "0111111111010000",
59631 => "0111111111010000",
59632 => "0111111111010000",
59633 => "0111111111010000",
59634 => "0111111111010000",
59635 => "0111111111010000",
59636 => "0111111111010000",
59637 => "0111111111010000",
59638 => "0111111111010000",
59639 => "0111111111010000",
59640 => "0111111111010000",
59641 => "0111111111010000",
59642 => "0111111111010000",
59643 => "0111111111010000",
59644 => "0111111111010000",
59645 => "0111111111010000",
59646 => "0111111111010000",
59647 => "0111111111010000",
59648 => "0111111111010000",
59649 => "0111111111010000",
59650 => "0111111111010000",
59651 => "0111111111010000",
59652 => "0111111111010000",
59653 => "0111111111010000",
59654 => "0111111111010000",
59655 => "0111111111010000",
59656 => "0111111111010000",
59657 => "0111111111010000",
59658 => "0111111111010000",
59659 => "0111111111010000",
59660 => "0111111111010000",
59661 => "0111111111010000",
59662 => "0111111111010000",
59663 => "0111111111010000",
59664 => "0111111111010000",
59665 => "0111111111010000",
59666 => "0111111111010000",
59667 => "0111111111010000",
59668 => "0111111111010000",
59669 => "0111111111010000",
59670 => "0111111111010000",
59671 => "0111111111010000",
59672 => "0111111111010000",
59673 => "0111111111010000",
59674 => "0111111111010000",
59675 => "0111111111010000",
59676 => "0111111111010000",
59677 => "0111111111010000",
59678 => "0111111111010000",
59679 => "0111111111010000",
59680 => "0111111111010000",
59681 => "0111111111010000",
59682 => "0111111111010000",
59683 => "0111111111010000",
59684 => "0111111111010000",
59685 => "0111111111010000",
59686 => "0111111111010000",
59687 => "0111111111010000",
59688 => "0111111111010000",
59689 => "0111111111010000",
59690 => "0111111111010000",
59691 => "0111111111010000",
59692 => "0111111111010000",
59693 => "0111111111010000",
59694 => "0111111111010000",
59695 => "0111111111010000",
59696 => "0111111111010000",
59697 => "0111111111010000",
59698 => "0111111111010000",
59699 => "0111111111010000",
59700 => "0111111111010000",
59701 => "0111111111010000",
59702 => "0111111111010000",
59703 => "0111111111010000",
59704 => "0111111111010000",
59705 => "0111111111010000",
59706 => "0111111111010000",
59707 => "0111111111010000",
59708 => "0111111111010000",
59709 => "0111111111010000",
59710 => "0111111111010000",
59711 => "0111111111010000",
59712 => "0111111111010000",
59713 => "0111111111010000",
59714 => "0111111111010000",
59715 => "0111111111010000",
59716 => "0111111111010000",
59717 => "0111111111010000",
59718 => "0111111111010000",
59719 => "0111111111010000",
59720 => "0111111111010000",
59721 => "0111111111010000",
59722 => "0111111111010000",
59723 => "0111111111010000",
59724 => "0111111111010000",
59725 => "0111111111010000",
59726 => "0111111111010000",
59727 => "0111111111010000",
59728 => "0111111111010000",
59729 => "0111111111010000",
59730 => "0111111111010000",
59731 => "0111111111010000",
59732 => "0111111111010000",
59733 => "0111111111010000",
59734 => "0111111111010000",
59735 => "0111111111010000",
59736 => "0111111111010000",
59737 => "0111111111010000",
59738 => "0111111111010000",
59739 => "0111111111010000",
59740 => "0111111111010000",
59741 => "0111111111010000",
59742 => "0111111111010000",
59743 => "0111111111010000",
59744 => "0111111111010000",
59745 => "0111111111010000",
59746 => "0111111111010000",
59747 => "0111111111010000",
59748 => "0111111111010000",
59749 => "0111111111010000",
59750 => "0111111111010000",
59751 => "0111111111010000",
59752 => "0111111111010000",
59753 => "0111111111010000",
59754 => "0111111111010000",
59755 => "0111111111010000",
59756 => "0111111111010000",
59757 => "0111111111010000",
59758 => "0111111111010000",
59759 => "0111111111010000",
59760 => "0111111111010000",
59761 => "0111111111010000",
59762 => "0111111111010000",
59763 => "0111111111010000",
59764 => "0111111111010000",
59765 => "0111111111010000",
59766 => "0111111111010000",
59767 => "0111111111010000",
59768 => "0111111111010000",
59769 => "0111111111010000",
59770 => "0111111111010000",
59771 => "0111111111010000",
59772 => "0111111111010000",
59773 => "0111111111010000",
59774 => "0111111111010000",
59775 => "0111111111010000",
59776 => "0111111111010000",
59777 => "0111111111010000",
59778 => "0111111111010000",
59779 => "0111111111010000",
59780 => "0111111111010000",
59781 => "0111111111010000",
59782 => "0111111111010000",
59783 => "0111111111010000",
59784 => "0111111111010000",
59785 => "0111111111010000",
59786 => "0111111111010000",
59787 => "0111111111010000",
59788 => "0111111111010000",
59789 => "0111111111010000",
59790 => "0111111111010000",
59791 => "0111111111010000",
59792 => "0111111111010000",
59793 => "0111111111010000",
59794 => "0111111111010000",
59795 => "0111111111010000",
59796 => "0111111111010000",
59797 => "0111111111010000",
59798 => "0111111111010000",
59799 => "0111111111010000",
59800 => "0111111111010000",
59801 => "0111111111010000",
59802 => "0111111111010000",
59803 => "0111111111010000",
59804 => "0111111111010000",
59805 => "0111111111010000",
59806 => "0111111111010000",
59807 => "0111111111010000",
59808 => "0111111111010000",
59809 => "0111111111010000",
59810 => "0111111111010000",
59811 => "0111111111010000",
59812 => "0111111111010000",
59813 => "0111111111010000",
59814 => "0111111111010000",
59815 => "0111111111010000",
59816 => "0111111111010000",
59817 => "0111111111010000",
59818 => "0111111111010000",
59819 => "0111111111010000",
59820 => "0111111111010000",
59821 => "0111111111010000",
59822 => "0111111111010000",
59823 => "0111111111010000",
59824 => "0111111111010000",
59825 => "0111111111010000",
59826 => "0111111111010000",
59827 => "0111111111010000",
59828 => "0111111111010000",
59829 => "0111111111010000",
59830 => "0111111111010000",
59831 => "0111111111010000",
59832 => "0111111111010000",
59833 => "0111111111010000",
59834 => "0111111111010000",
59835 => "0111111111010000",
59836 => "0111111111010000",
59837 => "0111111111010000",
59838 => "0111111111010000",
59839 => "0111111111010000",
59840 => "0111111111010000",
59841 => "0111111111010000",
59842 => "0111111111010000",
59843 => "0111111111010000",
59844 => "0111111111010000",
59845 => "0111111111010000",
59846 => "0111111111010000",
59847 => "0111111111010000",
59848 => "0111111111010000",
59849 => "0111111111010000",
59850 => "0111111111010000",
59851 => "0111111111010000",
59852 => "0111111111010000",
59853 => "0111111111010000",
59854 => "0111111111010000",
59855 => "0111111111010000",
59856 => "0111111111010000",
59857 => "0111111111010000",
59858 => "0111111111010000",
59859 => "0111111111010000",
59860 => "0111111111010000",
59861 => "0111111111010000",
59862 => "0111111111010000",
59863 => "0111111111010000",
59864 => "0111111111010000",
59865 => "0111111111010000",
59866 => "0111111111010000",
59867 => "0111111111010000",
59868 => "0111111111010000",
59869 => "0111111111010000",
59870 => "0111111111010000",
59871 => "0111111111010000",
59872 => "0111111111010000",
59873 => "0111111111010000",
59874 => "0111111111010000",
59875 => "0111111111010000",
59876 => "0111111111010000",
59877 => "0111111111010000",
59878 => "0111111111010000",
59879 => "0111111111010000",
59880 => "0111111111010000",
59881 => "0111111111010000",
59882 => "0111111111010000",
59883 => "0111111111010000",
59884 => "0111111111010000",
59885 => "0111111111010000",
59886 => "0111111111010000",
59887 => "0111111111010000",
59888 => "0111111111010000",
59889 => "0111111111010000",
59890 => "0111111111010000",
59891 => "0111111111010000",
59892 => "0111111111010000",
59893 => "0111111111010000",
59894 => "0111111111010000",
59895 => "0111111111010000",
59896 => "0111111111010000",
59897 => "0111111111010000",
59898 => "0111111111010000",
59899 => "0111111111010000",
59900 => "0111111111010000",
59901 => "0111111111010000",
59902 => "0111111111010000",
59903 => "0111111111010000",
59904 => "0111111111010000",
59905 => "0111111111010000",
59906 => "0111111111010000",
59907 => "0111111111010000",
59908 => "0111111111010000",
59909 => "0111111111010000",
59910 => "0111111111010000",
59911 => "0111111111010000",
59912 => "0111111111010000",
59913 => "0111111111010000",
59914 => "0111111111010000",
59915 => "0111111111010000",
59916 => "0111111111010000",
59917 => "0111111111010000",
59918 => "0111111111010000",
59919 => "0111111111010000",
59920 => "0111111111010000",
59921 => "0111111111010000",
59922 => "0111111111010000",
59923 => "0111111111010000",
59924 => "0111111111010000",
59925 => "0111111111010000",
59926 => "0111111111010000",
59927 => "0111111111010000",
59928 => "0111111111010000",
59929 => "0111111111010000",
59930 => "0111111111010000",
59931 => "0111111111010000",
59932 => "0111111111010000",
59933 => "0111111111010000",
59934 => "0111111111010000",
59935 => "0111111111010000",
59936 => "0111111111010000",
59937 => "0111111111010000",
59938 => "0111111111010000",
59939 => "0111111111010000",
59940 => "0111111111010000",
59941 => "0111111111010000",
59942 => "0111111111010000",
59943 => "0111111111010000",
59944 => "0111111111010000",
59945 => "0111111111010000",
59946 => "0111111111010000",
59947 => "0111111111010000",
59948 => "0111111111010000",
59949 => "0111111111010000",
59950 => "0111111111010000",
59951 => "0111111111010000",
59952 => "0111111111010000",
59953 => "0111111111010000",
59954 => "0111111111010000",
59955 => "0111111111010000",
59956 => "0111111111010000",
59957 => "0111111111010000",
59958 => "0111111111010000",
59959 => "0111111111010000",
59960 => "0111111111010000",
59961 => "0111111111010000",
59962 => "0111111111010000",
59963 => "0111111111010000",
59964 => "0111111111010000",
59965 => "0111111111010000",
59966 => "0111111111010000",
59967 => "0111111111010000",
59968 => "0111111111010000",
59969 => "0111111111010000",
59970 => "0111111111010000",
59971 => "0111111111010000",
59972 => "0111111111010000",
59973 => "0111111111010000",
59974 => "0111111111010000",
59975 => "0111111111010000",
59976 => "0111111111010000",
59977 => "0111111111010000",
59978 => "0111111111010000",
59979 => "0111111111010000",
59980 => "0111111111010000",
59981 => "0111111111010000",
59982 => "0111111111010000",
59983 => "0111111111010000",
59984 => "0111111111010000",
59985 => "0111111111010000",
59986 => "0111111111010000",
59987 => "0111111111010000",
59988 => "0111111111010000",
59989 => "0111111111010000",
59990 => "0111111111010000",
59991 => "0111111111010000",
59992 => "0111111111010000",
59993 => "0111111111010000",
59994 => "0111111111010000",
59995 => "0111111111010000",
59996 => "0111111111010000",
59997 => "0111111111010000",
59998 => "0111111111010000",
59999 => "0111111111010000",
60000 => "0111111111010000",
60001 => "0111111111010000",
60002 => "0111111111010000",
60003 => "0111111111010000",
60004 => "0111111111010000",
60005 => "0111111111010000",
60006 => "0111111111010000",
60007 => "0111111111010000",
60008 => "0111111111010000",
60009 => "0111111111010000",
60010 => "0111111111010000",
60011 => "0111111111010000",
60012 => "0111111111010000",
60013 => "0111111111010000",
60014 => "0111111111010000",
60015 => "0111111111010000",
60016 => "0111111111010000",
60017 => "0111111111010000",
60018 => "0111111111010000",
60019 => "0111111111010000",
60020 => "0111111111010000",
60021 => "0111111111010000",
60022 => "0111111111010000",
60023 => "0111111111010000",
60024 => "0111111111010000",
60025 => "0111111111010000",
60026 => "0111111111010000",
60027 => "0111111111010000",
60028 => "0111111111010000",
60029 => "0111111111010000",
60030 => "0111111111010000",
60031 => "0111111111010000",
60032 => "0111111111010000",
60033 => "0111111111010000",
60034 => "0111111111010000",
60035 => "0111111111010000",
60036 => "0111111111010000",
60037 => "0111111111010000",
60038 => "0111111111010000",
60039 => "0111111111010000",
60040 => "0111111111010000",
60041 => "0111111111010000",
60042 => "0111111111010000",
60043 => "0111111111010000",
60044 => "0111111111010000",
60045 => "0111111111010000",
60046 => "0111111111010000",
60047 => "0111111111010000",
60048 => "0111111111010000",
60049 => "0111111111010000",
60050 => "0111111111010000",
60051 => "0111111111010000",
60052 => "0111111111010000",
60053 => "0111111111010000",
60054 => "0111111111010000",
60055 => "0111111111010000",
60056 => "0111111111010000",
60057 => "0111111111010000",
60058 => "0111111111010000",
60059 => "0111111111010000",
60060 => "0111111111010000",
60061 => "0111111111010000",
60062 => "0111111111010000",
60063 => "0111111111010000",
60064 => "0111111111010000",
60065 => "0111111111010000",
60066 => "0111111111010000",
60067 => "0111111111010000",
60068 => "0111111111010000",
60069 => "0111111111010000",
60070 => "0111111111010000",
60071 => "0111111111010000",
60072 => "0111111111010000",
60073 => "0111111111010000",
60074 => "0111111111010000",
60075 => "0111111111010000",
60076 => "0111111111010000",
60077 => "0111111111010000",
60078 => "0111111111010000",
60079 => "0111111111010000",
60080 => "0111111111010000",
60081 => "0111111111010000",
60082 => "0111111111010000",
60083 => "0111111111010000",
60084 => "0111111111010000",
60085 => "0111111111010000",
60086 => "0111111111010000",
60087 => "0111111111010000",
60088 => "0111111111010000",
60089 => "0111111111010000",
60090 => "0111111111010000",
60091 => "0111111111010000",
60092 => "0111111111010000",
60093 => "0111111111010000",
60094 => "0111111111010000",
60095 => "0111111111010000",
60096 => "0111111111010000",
60097 => "0111111111010000",
60098 => "0111111111010000",
60099 => "0111111111010000",
60100 => "0111111111010000",
60101 => "0111111111010000",
60102 => "0111111111010000",
60103 => "0111111111010000",
60104 => "0111111111010000",
60105 => "0111111111010000",
60106 => "0111111111010000",
60107 => "0111111111010000",
60108 => "0111111111010000",
60109 => "0111111111010000",
60110 => "0111111111010000",
60111 => "0111111111010000",
60112 => "0111111111010000",
60113 => "0111111111010000",
60114 => "0111111111010000",
60115 => "0111111111010000",
60116 => "0111111111010000",
60117 => "0111111111010000",
60118 => "0111111111010000",
60119 => "0111111111010000",
60120 => "0111111111010000",
60121 => "0111111111010000",
60122 => "0111111111010000",
60123 => "0111111111010000",
60124 => "0111111111010000",
60125 => "0111111111010000",
60126 => "0111111111010000",
60127 => "0111111111010000",
60128 => "0111111111010000",
60129 => "0111111111010000",
60130 => "0111111111010000",
60131 => "0111111111010000",
60132 => "0111111111010000",
60133 => "0111111111010000",
60134 => "0111111111010000",
60135 => "0111111111010000",
60136 => "0111111111010000",
60137 => "0111111111010000",
60138 => "0111111111010000",
60139 => "0111111111010000",
60140 => "0111111111010000",
60141 => "0111111111010000",
60142 => "0111111111010000",
60143 => "0111111111010000",
60144 => "0111111111010000",
60145 => "0111111111010000",
60146 => "0111111111010000",
60147 => "0111111111010000",
60148 => "0111111111010000",
60149 => "0111111111010000",
60150 => "0111111111010000",
60151 => "0111111111010000",
60152 => "0111111111010000",
60153 => "0111111111010000",
60154 => "0111111111010000",
60155 => "0111111111010000",
60156 => "0111111111010000",
60157 => "0111111111010000",
60158 => "0111111111010000",
60159 => "0111111111010000",
60160 => "0111111111010000",
60161 => "0111111111010000",
60162 => "0111111111010000",
60163 => "0111111111010000",
60164 => "0111111111010000",
60165 => "0111111111010000",
60166 => "0111111111010000",
60167 => "0111111111010000",
60168 => "0111111111010000",
60169 => "0111111111010000",
60170 => "0111111111010000",
60171 => "0111111111010000",
60172 => "0111111111010000",
60173 => "0111111111010000",
60174 => "0111111111010000",
60175 => "0111111111010000",
60176 => "0111111111010000",
60177 => "0111111111010000",
60178 => "0111111111010000",
60179 => "0111111111010000",
60180 => "0111111111010000",
60181 => "0111111111010000",
60182 => "0111111111010000",
60183 => "0111111111010000",
60184 => "0111111111010000",
60185 => "0111111111010000",
60186 => "0111111111010000",
60187 => "0111111111010000",
60188 => "0111111111010000",
60189 => "0111111111010000",
60190 => "0111111111010000",
60191 => "0111111111010000",
60192 => "0111111111010000",
60193 => "0111111111010000",
60194 => "0111111111010000",
60195 => "0111111111010000",
60196 => "0111111111010000",
60197 => "0111111111010000",
60198 => "0111111111010000",
60199 => "0111111111010000",
60200 => "0111111111010000",
60201 => "0111111111010000",
60202 => "0111111111010000",
60203 => "0111111111010000",
60204 => "0111111111010000",
60205 => "0111111111010000",
60206 => "0111111111010000",
60207 => "0111111111010000",
60208 => "0111111111010000",
60209 => "0111111111010000",
60210 => "0111111111010000",
60211 => "0111111111010000",
60212 => "0111111111010000",
60213 => "0111111111010000",
60214 => "0111111111010000",
60215 => "0111111111010000",
60216 => "0111111111010000",
60217 => "0111111111010000",
60218 => "0111111111010000",
60219 => "0111111111010000",
60220 => "0111111111010000",
60221 => "0111111111010000",
60222 => "0111111111010000",
60223 => "0111111111010000",
60224 => "0111111111010000",
60225 => "0111111111010000",
60226 => "0111111111010000",
60227 => "0111111111010000",
60228 => "0111111111010000",
60229 => "0111111111010000",
60230 => "0111111111010000",
60231 => "0111111111010000",
60232 => "0111111111010000",
60233 => "0111111111010000",
60234 => "0111111111010000",
60235 => "0111111111010000",
60236 => "0111111111010000",
60237 => "0111111111010000",
60238 => "0111111111010000",
60239 => "0111111111010000",
60240 => "0111111111100000",
60241 => "0111111111100000",
60242 => "0111111111100000",
60243 => "0111111111100000",
60244 => "0111111111100000",
60245 => "0111111111100000",
60246 => "0111111111100000",
60247 => "0111111111100000",
60248 => "0111111111100000",
60249 => "0111111111100000",
60250 => "0111111111100000",
60251 => "0111111111100000",
60252 => "0111111111100000",
60253 => "0111111111100000",
60254 => "0111111111100000",
60255 => "0111111111100000",
60256 => "0111111111100000",
60257 => "0111111111100000",
60258 => "0111111111100000",
60259 => "0111111111100000",
60260 => "0111111111100000",
60261 => "0111111111100000",
60262 => "0111111111100000",
60263 => "0111111111100000",
60264 => "0111111111100000",
60265 => "0111111111100000",
60266 => "0111111111100000",
60267 => "0111111111100000",
60268 => "0111111111100000",
60269 => "0111111111100000",
60270 => "0111111111100000",
60271 => "0111111111100000",
60272 => "0111111111100000",
60273 => "0111111111100000",
60274 => "0111111111100000",
60275 => "0111111111100000",
60276 => "0111111111100000",
60277 => "0111111111100000",
60278 => "0111111111100000",
60279 => "0111111111100000",
60280 => "0111111111100000",
60281 => "0111111111100000",
60282 => "0111111111100000",
60283 => "0111111111100000",
60284 => "0111111111100000",
60285 => "0111111111100000",
60286 => "0111111111100000",
60287 => "0111111111100000",
60288 => "0111111111100000",
60289 => "0111111111100000",
60290 => "0111111111100000",
60291 => "0111111111100000",
60292 => "0111111111100000",
60293 => "0111111111100000",
60294 => "0111111111100000",
60295 => "0111111111100000",
60296 => "0111111111100000",
60297 => "0111111111100000",
60298 => "0111111111100000",
60299 => "0111111111100000",
60300 => "0111111111100000",
60301 => "0111111111100000",
60302 => "0111111111100000",
60303 => "0111111111100000",
60304 => "0111111111100000",
60305 => "0111111111100000",
60306 => "0111111111100000",
60307 => "0111111111100000",
60308 => "0111111111100000",
60309 => "0111111111100000",
60310 => "0111111111100000",
60311 => "0111111111100000",
60312 => "0111111111100000",
60313 => "0111111111100000",
60314 => "0111111111100000",
60315 => "0111111111100000",
60316 => "0111111111100000",
60317 => "0111111111100000",
60318 => "0111111111100000",
60319 => "0111111111100000",
60320 => "0111111111100000",
60321 => "0111111111100000",
60322 => "0111111111100000",
60323 => "0111111111100000",
60324 => "0111111111100000",
60325 => "0111111111100000",
60326 => "0111111111100000",
60327 => "0111111111100000",
60328 => "0111111111100000",
60329 => "0111111111100000",
60330 => "0111111111100000",
60331 => "0111111111100000",
60332 => "0111111111100000",
60333 => "0111111111100000",
60334 => "0111111111100000",
60335 => "0111111111100000",
60336 => "0111111111100000",
60337 => "0111111111100000",
60338 => "0111111111100000",
60339 => "0111111111100000",
60340 => "0111111111100000",
60341 => "0111111111100000",
60342 => "0111111111100000",
60343 => "0111111111100000",
60344 => "0111111111100000",
60345 => "0111111111100000",
60346 => "0111111111100000",
60347 => "0111111111100000",
60348 => "0111111111100000",
60349 => "0111111111100000",
60350 => "0111111111100000",
60351 => "0111111111100000",
60352 => "0111111111100000",
60353 => "0111111111100000",
60354 => "0111111111100000",
60355 => "0111111111100000",
60356 => "0111111111100000",
60357 => "0111111111100000",
60358 => "0111111111100000",
60359 => "0111111111100000",
60360 => "0111111111100000",
60361 => "0111111111100000",
60362 => "0111111111100000",
60363 => "0111111111100000",
60364 => "0111111111100000",
60365 => "0111111111100000",
60366 => "0111111111100000",
60367 => "0111111111100000",
60368 => "0111111111100000",
60369 => "0111111111100000",
60370 => "0111111111100000",
60371 => "0111111111100000",
60372 => "0111111111100000",
60373 => "0111111111100000",
60374 => "0111111111100000",
60375 => "0111111111100000",
60376 => "0111111111100000",
60377 => "0111111111100000",
60378 => "0111111111100000",
60379 => "0111111111100000",
60380 => "0111111111100000",
60381 => "0111111111100000",
60382 => "0111111111100000",
60383 => "0111111111100000",
60384 => "0111111111100000",
60385 => "0111111111100000",
60386 => "0111111111100000",
60387 => "0111111111100000",
60388 => "0111111111100000",
60389 => "0111111111100000",
60390 => "0111111111100000",
60391 => "0111111111100000",
60392 => "0111111111100000",
60393 => "0111111111100000",
60394 => "0111111111100000",
60395 => "0111111111100000",
60396 => "0111111111100000",
60397 => "0111111111100000",
60398 => "0111111111100000",
60399 => "0111111111100000",
60400 => "0111111111100000",
60401 => "0111111111100000",
60402 => "0111111111100000",
60403 => "0111111111100000",
60404 => "0111111111100000",
60405 => "0111111111100000",
60406 => "0111111111100000",
60407 => "0111111111100000",
60408 => "0111111111100000",
60409 => "0111111111100000",
60410 => "0111111111100000",
60411 => "0111111111100000",
60412 => "0111111111100000",
60413 => "0111111111100000",
60414 => "0111111111100000",
60415 => "0111111111100000",
60416 => "0111111111100000",
60417 => "0111111111100000",
60418 => "0111111111100000",
60419 => "0111111111100000",
60420 => "0111111111100000",
60421 => "0111111111100000",
60422 => "0111111111100000",
60423 => "0111111111100000",
60424 => "0111111111100000",
60425 => "0111111111100000",
60426 => "0111111111100000",
60427 => "0111111111100000",
60428 => "0111111111100000",
60429 => "0111111111100000",
60430 => "0111111111100000",
60431 => "0111111111100000",
60432 => "0111111111100000",
60433 => "0111111111100000",
60434 => "0111111111100000",
60435 => "0111111111100000",
60436 => "0111111111100000",
60437 => "0111111111100000",
60438 => "0111111111100000",
60439 => "0111111111100000",
60440 => "0111111111100000",
60441 => "0111111111100000",
60442 => "0111111111100000",
60443 => "0111111111100000",
60444 => "0111111111100000",
60445 => "0111111111100000",
60446 => "0111111111100000",
60447 => "0111111111100000",
60448 => "0111111111100000",
60449 => "0111111111100000",
60450 => "0111111111100000",
60451 => "0111111111100000",
60452 => "0111111111100000",
60453 => "0111111111100000",
60454 => "0111111111100000",
60455 => "0111111111100000",
60456 => "0111111111100000",
60457 => "0111111111100000",
60458 => "0111111111100000",
60459 => "0111111111100000",
60460 => "0111111111100000",
60461 => "0111111111100000",
60462 => "0111111111100000",
60463 => "0111111111100000",
60464 => "0111111111100000",
60465 => "0111111111100000",
60466 => "0111111111100000",
60467 => "0111111111100000",
60468 => "0111111111100000",
60469 => "0111111111100000",
60470 => "0111111111100000",
60471 => "0111111111100000",
60472 => "0111111111100000",
60473 => "0111111111100000",
60474 => "0111111111100000",
60475 => "0111111111100000",
60476 => "0111111111100000",
60477 => "0111111111100000",
60478 => "0111111111100000",
60479 => "0111111111100000",
60480 => "0111111111100000",
60481 => "0111111111100000",
60482 => "0111111111100000",
60483 => "0111111111100000",
60484 => "0111111111100000",
60485 => "0111111111100000",
60486 => "0111111111100000",
60487 => "0111111111100000",
60488 => "0111111111100000",
60489 => "0111111111100000",
60490 => "0111111111100000",
60491 => "0111111111100000",
60492 => "0111111111100000",
60493 => "0111111111100000",
60494 => "0111111111100000",
60495 => "0111111111100000",
60496 => "0111111111100000",
60497 => "0111111111100000",
60498 => "0111111111100000",
60499 => "0111111111100000",
60500 => "0111111111100000",
60501 => "0111111111100000",
60502 => "0111111111100000",
60503 => "0111111111100000",
60504 => "0111111111100000",
60505 => "0111111111100000",
60506 => "0111111111100000",
60507 => "0111111111100000",
60508 => "0111111111100000",
60509 => "0111111111100000",
60510 => "0111111111100000",
60511 => "0111111111100000",
60512 => "0111111111100000",
60513 => "0111111111100000",
60514 => "0111111111100000",
60515 => "0111111111100000",
60516 => "0111111111100000",
60517 => "0111111111100000",
60518 => "0111111111100000",
60519 => "0111111111100000",
60520 => "0111111111100000",
60521 => "0111111111100000",
60522 => "0111111111100000",
60523 => "0111111111100000",
60524 => "0111111111100000",
60525 => "0111111111100000",
60526 => "0111111111100000",
60527 => "0111111111100000",
60528 => "0111111111100000",
60529 => "0111111111100000",
60530 => "0111111111100000",
60531 => "0111111111100000",
60532 => "0111111111100000",
60533 => "0111111111100000",
60534 => "0111111111100000",
60535 => "0111111111100000",
60536 => "0111111111100000",
60537 => "0111111111100000",
60538 => "0111111111100000",
60539 => "0111111111100000",
60540 => "0111111111100000",
60541 => "0111111111100000",
60542 => "0111111111100000",
60543 => "0111111111100000",
60544 => "0111111111100000",
60545 => "0111111111100000",
60546 => "0111111111100000",
60547 => "0111111111100000",
60548 => "0111111111100000",
60549 => "0111111111100000",
60550 => "0111111111100000",
60551 => "0111111111100000",
60552 => "0111111111100000",
60553 => "0111111111100000",
60554 => "0111111111100000",
60555 => "0111111111100000",
60556 => "0111111111100000",
60557 => "0111111111100000",
60558 => "0111111111100000",
60559 => "0111111111100000",
60560 => "0111111111100000",
60561 => "0111111111100000",
60562 => "0111111111100000",
60563 => "0111111111100000",
60564 => "0111111111100000",
60565 => "0111111111100000",
60566 => "0111111111100000",
60567 => "0111111111100000",
60568 => "0111111111100000",
60569 => "0111111111100000",
60570 => "0111111111100000",
60571 => "0111111111100000",
60572 => "0111111111100000",
60573 => "0111111111100000",
60574 => "0111111111100000",
60575 => "0111111111100000",
60576 => "0111111111100000",
60577 => "0111111111100000",
60578 => "0111111111100000",
60579 => "0111111111100000",
60580 => "0111111111100000",
60581 => "0111111111100000",
60582 => "0111111111100000",
60583 => "0111111111100000",
60584 => "0111111111100000",
60585 => "0111111111100000",
60586 => "0111111111100000",
60587 => "0111111111100000",
60588 => "0111111111100000",
60589 => "0111111111100000",
60590 => "0111111111100000",
60591 => "0111111111100000",
60592 => "0111111111100000",
60593 => "0111111111100000",
60594 => "0111111111100000",
60595 => "0111111111100000",
60596 => "0111111111100000",
60597 => "0111111111100000",
60598 => "0111111111100000",
60599 => "0111111111100000",
60600 => "0111111111100000",
60601 => "0111111111100000",
60602 => "0111111111100000",
60603 => "0111111111100000",
60604 => "0111111111100000",
60605 => "0111111111100000",
60606 => "0111111111100000",
60607 => "0111111111100000",
60608 => "0111111111100000",
60609 => "0111111111100000",
60610 => "0111111111100000",
60611 => "0111111111100000",
60612 => "0111111111100000",
60613 => "0111111111100000",
60614 => "0111111111100000",
60615 => "0111111111100000",
60616 => "0111111111100000",
60617 => "0111111111100000",
60618 => "0111111111100000",
60619 => "0111111111100000",
60620 => "0111111111100000",
60621 => "0111111111100000",
60622 => "0111111111100000",
60623 => "0111111111100000",
60624 => "0111111111100000",
60625 => "0111111111100000",
60626 => "0111111111100000",
60627 => "0111111111100000",
60628 => "0111111111100000",
60629 => "0111111111100000",
60630 => "0111111111100000",
60631 => "0111111111100000",
60632 => "0111111111100000",
60633 => "0111111111100000",
60634 => "0111111111100000",
60635 => "0111111111100000",
60636 => "0111111111100000",
60637 => "0111111111100000",
60638 => "0111111111100000",
60639 => "0111111111100000",
60640 => "0111111111100000",
60641 => "0111111111100000",
60642 => "0111111111100000",
60643 => "0111111111100000",
60644 => "0111111111100000",
60645 => "0111111111100000",
60646 => "0111111111100000",
60647 => "0111111111100000",
60648 => "0111111111100000",
60649 => "0111111111100000",
60650 => "0111111111100000",
60651 => "0111111111100000",
60652 => "0111111111100000",
60653 => "0111111111100000",
60654 => "0111111111100000",
60655 => "0111111111100000",
60656 => "0111111111100000",
60657 => "0111111111100000",
60658 => "0111111111100000",
60659 => "0111111111100000",
60660 => "0111111111100000",
60661 => "0111111111100000",
60662 => "0111111111100000",
60663 => "0111111111100000",
60664 => "0111111111100000",
60665 => "0111111111100000",
60666 => "0111111111100000",
60667 => "0111111111100000",
60668 => "0111111111100000",
60669 => "0111111111100000",
60670 => "0111111111100000",
60671 => "0111111111100000",
60672 => "0111111111100000",
60673 => "0111111111100000",
60674 => "0111111111100000",
60675 => "0111111111100000",
60676 => "0111111111100000",
60677 => "0111111111100000",
60678 => "0111111111100000",
60679 => "0111111111100000",
60680 => "0111111111100000",
60681 => "0111111111100000",
60682 => "0111111111100000",
60683 => "0111111111100000",
60684 => "0111111111100000",
60685 => "0111111111100000",
60686 => "0111111111100000",
60687 => "0111111111100000",
60688 => "0111111111100000",
60689 => "0111111111100000",
60690 => "0111111111100000",
60691 => "0111111111100000",
60692 => "0111111111100000",
60693 => "0111111111100000",
60694 => "0111111111100000",
60695 => "0111111111100000",
60696 => "0111111111100000",
60697 => "0111111111100000",
60698 => "0111111111100000",
60699 => "0111111111100000",
60700 => "0111111111100000",
60701 => "0111111111100000",
60702 => "0111111111100000",
60703 => "0111111111100000",
60704 => "0111111111100000",
60705 => "0111111111100000",
60706 => "0111111111100000",
60707 => "0111111111100000",
60708 => "0111111111100000",
60709 => "0111111111100000",
60710 => "0111111111100000",
60711 => "0111111111100000",
60712 => "0111111111100000",
60713 => "0111111111100000",
60714 => "0111111111100000",
60715 => "0111111111100000",
60716 => "0111111111100000",
60717 => "0111111111100000",
60718 => "0111111111100000",
60719 => "0111111111100000",
60720 => "0111111111100000",
60721 => "0111111111100000",
60722 => "0111111111100000",
60723 => "0111111111100000",
60724 => "0111111111100000",
60725 => "0111111111100000",
60726 => "0111111111100000",
60727 => "0111111111100000",
60728 => "0111111111100000",
60729 => "0111111111100000",
60730 => "0111111111100000",
60731 => "0111111111100000",
60732 => "0111111111100000",
60733 => "0111111111100000",
60734 => "0111111111100000",
60735 => "0111111111100000",
60736 => "0111111111100000",
60737 => "0111111111100000",
60738 => "0111111111100000",
60739 => "0111111111100000",
60740 => "0111111111100000",
60741 => "0111111111100000",
60742 => "0111111111100000",
60743 => "0111111111100000",
60744 => "0111111111100000",
60745 => "0111111111100000",
60746 => "0111111111100000",
60747 => "0111111111100000",
60748 => "0111111111100000",
60749 => "0111111111100000",
60750 => "0111111111100000",
60751 => "0111111111100000",
60752 => "0111111111100000",
60753 => "0111111111100000",
60754 => "0111111111100000",
60755 => "0111111111100000",
60756 => "0111111111100000",
60757 => "0111111111100000",
60758 => "0111111111100000",
60759 => "0111111111100000",
60760 => "0111111111100000",
60761 => "0111111111100000",
60762 => "0111111111100000",
60763 => "0111111111100000",
60764 => "0111111111100000",
60765 => "0111111111100000",
60766 => "0111111111100000",
60767 => "0111111111100000",
60768 => "0111111111100000",
60769 => "0111111111100000",
60770 => "0111111111100000",
60771 => "0111111111100000",
60772 => "0111111111100000",
60773 => "0111111111100000",
60774 => "0111111111100000",
60775 => "0111111111100000",
60776 => "0111111111100000",
60777 => "0111111111100000",
60778 => "0111111111100000",
60779 => "0111111111100000",
60780 => "0111111111100000",
60781 => "0111111111100000",
60782 => "0111111111100000",
60783 => "0111111111100000",
60784 => "0111111111100000",
60785 => "0111111111100000",
60786 => "0111111111100000",
60787 => "0111111111100000",
60788 => "0111111111100000",
60789 => "0111111111100000",
60790 => "0111111111100000",
60791 => "0111111111100000",
60792 => "0111111111100000",
60793 => "0111111111100000",
60794 => "0111111111100000",
60795 => "0111111111100000",
60796 => "0111111111100000",
60797 => "0111111111100000",
60798 => "0111111111100000",
60799 => "0111111111100000",
60800 => "0111111111100000",
60801 => "0111111111100000",
60802 => "0111111111100000",
60803 => "0111111111100000",
60804 => "0111111111100000",
60805 => "0111111111100000",
60806 => "0111111111100000",
60807 => "0111111111100000",
60808 => "0111111111100000",
60809 => "0111111111100000",
60810 => "0111111111100000",
60811 => "0111111111100000",
60812 => "0111111111100000",
60813 => "0111111111100000",
60814 => "0111111111100000",
60815 => "0111111111100000",
60816 => "0111111111100000",
60817 => "0111111111100000",
60818 => "0111111111100000",
60819 => "0111111111100000",
60820 => "0111111111100000",
60821 => "0111111111100000",
60822 => "0111111111100000",
60823 => "0111111111100000",
60824 => "0111111111100000",
60825 => "0111111111100000",
60826 => "0111111111100000",
60827 => "0111111111100000",
60828 => "0111111111100000",
60829 => "0111111111100000",
60830 => "0111111111100000",
60831 => "0111111111100000",
60832 => "0111111111100000",
60833 => "0111111111100000",
60834 => "0111111111100000",
60835 => "0111111111100000",
60836 => "0111111111100000",
60837 => "0111111111100000",
60838 => "0111111111100000",
60839 => "0111111111100000",
60840 => "0111111111100000",
60841 => "0111111111100000",
60842 => "0111111111100000",
60843 => "0111111111100000",
60844 => "0111111111100000",
60845 => "0111111111100000",
60846 => "0111111111100000",
60847 => "0111111111100000",
60848 => "0111111111100000",
60849 => "0111111111100000",
60850 => "0111111111100000",
60851 => "0111111111100000",
60852 => "0111111111100000",
60853 => "0111111111100000",
60854 => "0111111111100000",
60855 => "0111111111100000",
60856 => "0111111111100000",
60857 => "0111111111100000",
60858 => "0111111111100000",
60859 => "0111111111100000",
60860 => "0111111111100000",
60861 => "0111111111100000",
60862 => "0111111111100000",
60863 => "0111111111100000",
60864 => "0111111111100000",
60865 => "0111111111100000",
60866 => "0111111111100000",
60867 => "0111111111100000",
60868 => "0111111111100000",
60869 => "0111111111100000",
60870 => "0111111111100000",
60871 => "0111111111100000",
60872 => "0111111111100000",
60873 => "0111111111100000",
60874 => "0111111111100000",
60875 => "0111111111100000",
60876 => "0111111111100000",
60877 => "0111111111100000",
60878 => "0111111111100000",
60879 => "0111111111100000",
60880 => "0111111111100000",
60881 => "0111111111100000",
60882 => "0111111111100000",
60883 => "0111111111100000",
60884 => "0111111111100000",
60885 => "0111111111100000",
60886 => "0111111111100000",
60887 => "0111111111100000",
60888 => "0111111111100000",
60889 => "0111111111100000",
60890 => "0111111111100000",
60891 => "0111111111100000",
60892 => "0111111111100000",
60893 => "0111111111100000",
60894 => "0111111111100000",
60895 => "0111111111100000",
60896 => "0111111111100000",
60897 => "0111111111100000",
60898 => "0111111111100000",
60899 => "0111111111100000",
60900 => "0111111111100000",
60901 => "0111111111100000",
60902 => "0111111111100000",
60903 => "0111111111100000",
60904 => "0111111111100000",
60905 => "0111111111100000",
60906 => "0111111111100000",
60907 => "0111111111100000",
60908 => "0111111111100000",
60909 => "0111111111100000",
60910 => "0111111111100000",
60911 => "0111111111100000",
60912 => "0111111111100000",
60913 => "0111111111100000",
60914 => "0111111111100000",
60915 => "0111111111100000",
60916 => "0111111111100000",
60917 => "0111111111100000",
60918 => "0111111111100000",
60919 => "0111111111100000",
60920 => "0111111111100000",
60921 => "0111111111100000",
60922 => "0111111111100000",
60923 => "0111111111100000",
60924 => "0111111111100000",
60925 => "0111111111100000",
60926 => "0111111111100000",
60927 => "0111111111100000",
60928 => "0111111111100000",
60929 => "0111111111100000",
60930 => "0111111111100000",
60931 => "0111111111100000",
60932 => "0111111111100000",
60933 => "0111111111100000",
60934 => "0111111111100000",
60935 => "0111111111100000",
60936 => "0111111111100000",
60937 => "0111111111100000",
60938 => "0111111111100000",
60939 => "0111111111100000",
60940 => "0111111111100000",
60941 => "0111111111100000",
60942 => "0111111111100000",
60943 => "0111111111100000",
60944 => "0111111111100000",
60945 => "0111111111100000",
60946 => "0111111111100000",
60947 => "0111111111100000",
60948 => "0111111111100000",
60949 => "0111111111100000",
60950 => "0111111111100000",
60951 => "0111111111100000",
60952 => "0111111111100000",
60953 => "0111111111100000",
60954 => "0111111111100000",
60955 => "0111111111100000",
60956 => "0111111111100000",
60957 => "0111111111100000",
60958 => "0111111111100000",
60959 => "0111111111100000",
60960 => "0111111111100000",
60961 => "0111111111100000",
60962 => "0111111111100000",
60963 => "0111111111100000",
60964 => "0111111111100000",
60965 => "0111111111100000",
60966 => "0111111111100000",
60967 => "0111111111100000",
60968 => "0111111111100000",
60969 => "0111111111100000",
60970 => "0111111111100000",
60971 => "0111111111100000",
60972 => "0111111111100000",
60973 => "0111111111100000",
60974 => "0111111111100000",
60975 => "0111111111100000",
60976 => "0111111111100000",
60977 => "0111111111100000",
60978 => "0111111111100000",
60979 => "0111111111100000",
60980 => "0111111111100000",
60981 => "0111111111100000",
60982 => "0111111111100000",
60983 => "0111111111100000",
60984 => "0111111111100000",
60985 => "0111111111100000",
60986 => "0111111111100000",
60987 => "0111111111100000",
60988 => "0111111111100000",
60989 => "0111111111100000",
60990 => "0111111111100000",
60991 => "0111111111100000",
60992 => "0111111111100000",
60993 => "0111111111100000",
60994 => "0111111111100000",
60995 => "0111111111100000",
60996 => "0111111111100000",
60997 => "0111111111100000",
60998 => "0111111111100000",
60999 => "0111111111100000",
61000 => "0111111111100000",
61001 => "0111111111100000",
61002 => "0111111111100000",
61003 => "0111111111100000",
61004 => "0111111111100000",
61005 => "0111111111100000",
61006 => "0111111111100000",
61007 => "0111111111100000",
61008 => "0111111111100000",
61009 => "0111111111100000",
61010 => "0111111111100000",
61011 => "0111111111100000",
61012 => "0111111111100000",
61013 => "0111111111100000",
61014 => "0111111111100000",
61015 => "0111111111100000",
61016 => "0111111111100000",
61017 => "0111111111100000",
61018 => "0111111111100000",
61019 => "0111111111100000",
61020 => "0111111111100000",
61021 => "0111111111100000",
61022 => "0111111111100000",
61023 => "0111111111100000",
61024 => "0111111111100000",
61025 => "0111111111100000",
61026 => "0111111111100000",
61027 => "0111111111100000",
61028 => "0111111111100000",
61029 => "0111111111100000",
61030 => "0111111111100000",
61031 => "0111111111100000",
61032 => "0111111111100000",
61033 => "0111111111100000",
61034 => "0111111111100000",
61035 => "0111111111100000",
61036 => "0111111111100000",
61037 => "0111111111100000",
61038 => "0111111111100000",
61039 => "0111111111100000",
61040 => "0111111111100000",
61041 => "0111111111100000",
61042 => "0111111111100000",
61043 => "0111111111100000",
61044 => "0111111111100000",
61045 => "0111111111100000",
61046 => "0111111111100000",
61047 => "0111111111100000",
61048 => "0111111111100000",
61049 => "0111111111100000",
61050 => "0111111111100000",
61051 => "0111111111100000",
61052 => "0111111111100000",
61053 => "0111111111100000",
61054 => "0111111111100000",
61055 => "0111111111100000",
61056 => "0111111111100000",
61057 => "0111111111100000",
61058 => "0111111111100000",
61059 => "0111111111100000",
61060 => "0111111111100000",
61061 => "0111111111100000",
61062 => "0111111111100000",
61063 => "0111111111100000",
61064 => "0111111111100000",
61065 => "0111111111100000",
61066 => "0111111111100000",
61067 => "0111111111100000",
61068 => "0111111111100000",
61069 => "0111111111100000",
61070 => "0111111111100000",
61071 => "0111111111100000",
61072 => "0111111111100000",
61073 => "0111111111100000",
61074 => "0111111111100000",
61075 => "0111111111100000",
61076 => "0111111111100000",
61077 => "0111111111100000",
61078 => "0111111111100000",
61079 => "0111111111100000",
61080 => "0111111111100000",
61081 => "0111111111100000",
61082 => "0111111111100000",
61083 => "0111111111100000",
61084 => "0111111111100000",
61085 => "0111111111100000",
61086 => "0111111111100000",
61087 => "0111111111100000",
61088 => "0111111111100000",
61089 => "0111111111100000",
61090 => "0111111111100000",
61091 => "0111111111100000",
61092 => "0111111111100000",
61093 => "0111111111100000",
61094 => "0111111111100000",
61095 => "0111111111100000",
61096 => "0111111111100000",
61097 => "0111111111100000",
61098 => "0111111111100000",
61099 => "0111111111100000",
61100 => "0111111111100000",
61101 => "0111111111100000",
61102 => "0111111111100000",
61103 => "0111111111100000",
61104 => "0111111111100000",
61105 => "0111111111100000",
61106 => "0111111111100000",
61107 => "0111111111100000",
61108 => "0111111111100000",
61109 => "0111111111100000",
61110 => "0111111111100000",
61111 => "0111111111100000",
61112 => "0111111111100000",
61113 => "0111111111100000",
61114 => "0111111111100000",
61115 => "0111111111100000",
61116 => "0111111111100000",
61117 => "0111111111100000",
61118 => "0111111111100000",
61119 => "0111111111100000",
61120 => "0111111111100000",
61121 => "0111111111100000",
61122 => "0111111111100000",
61123 => "0111111111100000",
61124 => "0111111111100000",
61125 => "0111111111100000",
61126 => "0111111111100000",
61127 => "0111111111100000",
61128 => "0111111111100000",
61129 => "0111111111100000",
61130 => "0111111111100000",
61131 => "0111111111100000",
61132 => "0111111111100000",
61133 => "0111111111100000",
61134 => "0111111111100000",
61135 => "0111111111100000",
61136 => "0111111111100000",
61137 => "0111111111100000",
61138 => "0111111111100000",
61139 => "0111111111100000",
61140 => "0111111111100000",
61141 => "0111111111100000",
61142 => "0111111111100000",
61143 => "0111111111100000",
61144 => "0111111111100000",
61145 => "0111111111100000",
61146 => "0111111111100000",
61147 => "0111111111100000",
61148 => "0111111111100000",
61149 => "0111111111100000",
61150 => "0111111111100000",
61151 => "0111111111100000",
61152 => "0111111111100000",
61153 => "0111111111100000",
61154 => "0111111111100000",
61155 => "0111111111100000",
61156 => "0111111111100000",
61157 => "0111111111100000",
61158 => "0111111111100000",
61159 => "0111111111100000",
61160 => "0111111111100000",
61161 => "0111111111100000",
61162 => "0111111111100000",
61163 => "0111111111100000",
61164 => "0111111111100000",
61165 => "0111111111100000",
61166 => "0111111111100000",
61167 => "0111111111100000",
61168 => "0111111111100000",
61169 => "0111111111100000",
61170 => "0111111111100000",
61171 => "0111111111100000",
61172 => "0111111111100000",
61173 => "0111111111100000",
61174 => "0111111111100000",
61175 => "0111111111100000",
61176 => "0111111111100000",
61177 => "0111111111100000",
61178 => "0111111111100000",
61179 => "0111111111100000",
61180 => "0111111111100000",
61181 => "0111111111100000",
61182 => "0111111111100000",
61183 => "0111111111100000",
61184 => "0111111111100000",
61185 => "0111111111100000",
61186 => "0111111111100000",
61187 => "0111111111100000",
61188 => "0111111111100000",
61189 => "0111111111100000",
61190 => "0111111111100000",
61191 => "0111111111100000",
61192 => "0111111111100000",
61193 => "0111111111100000",
61194 => "0111111111100000",
61195 => "0111111111100000",
61196 => "0111111111100000",
61197 => "0111111111100000",
61198 => "0111111111100000",
61199 => "0111111111100000",
61200 => "0111111111100000",
61201 => "0111111111100000",
61202 => "0111111111100000",
61203 => "0111111111100000",
61204 => "0111111111100000",
61205 => "0111111111100000",
61206 => "0111111111100000",
61207 => "0111111111100000",
61208 => "0111111111100000",
61209 => "0111111111100000",
61210 => "0111111111100000",
61211 => "0111111111100000",
61212 => "0111111111100000",
61213 => "0111111111100000",
61214 => "0111111111100000",
61215 => "0111111111100000",
61216 => "0111111111100000",
61217 => "0111111111100000",
61218 => "0111111111100000",
61219 => "0111111111100000",
61220 => "0111111111100000",
61221 => "0111111111100000",
61222 => "0111111111100000",
61223 => "0111111111100000",
61224 => "0111111111100000",
61225 => "0111111111100000",
61226 => "0111111111100000",
61227 => "0111111111100000",
61228 => "0111111111100000",
61229 => "0111111111100000",
61230 => "0111111111100000",
61231 => "0111111111100000",
61232 => "0111111111100000",
61233 => "0111111111100000",
61234 => "0111111111100000",
61235 => "0111111111100000",
61236 => "0111111111100000",
61237 => "0111111111100000",
61238 => "0111111111100000",
61239 => "0111111111100000",
61240 => "0111111111100000",
61241 => "0111111111100000",
61242 => "0111111111100000",
61243 => "0111111111100000",
61244 => "0111111111100000",
61245 => "0111111111100000",
61246 => "0111111111100000",
61247 => "0111111111100000",
61248 => "0111111111100000",
61249 => "0111111111100000",
61250 => "0111111111100000",
61251 => "0111111111100000",
61252 => "0111111111100000",
61253 => "0111111111100000",
61254 => "0111111111100000",
61255 => "0111111111100000",
61256 => "0111111111100000",
61257 => "0111111111100000",
61258 => "0111111111100000",
61259 => "0111111111100000",
61260 => "0111111111100000",
61261 => "0111111111100000",
61262 => "0111111111100000",
61263 => "0111111111100000",
61264 => "0111111111100000",
61265 => "0111111111100000",
61266 => "0111111111100000",
61267 => "0111111111100000",
61268 => "0111111111100000",
61269 => "0111111111100000",
61270 => "0111111111100000",
61271 => "0111111111100000",
61272 => "0111111111100000",
61273 => "0111111111100000",
61274 => "0111111111100000",
61275 => "0111111111100000",
61276 => "0111111111100000",
61277 => "0111111111100000",
61278 => "0111111111100000",
61279 => "0111111111100000",
61280 => "0111111111100000",
61281 => "0111111111100000",
61282 => "0111111111100000",
61283 => "0111111111100000",
61284 => "0111111111100000",
61285 => "0111111111100000",
61286 => "0111111111100000",
61287 => "0111111111100000",
61288 => "0111111111100000",
61289 => "0111111111100000",
61290 => "0111111111100000",
61291 => "0111111111100000",
61292 => "0111111111100000",
61293 => "0111111111100000",
61294 => "0111111111100000",
61295 => "0111111111100000",
61296 => "0111111111100000",
61297 => "0111111111100000",
61298 => "0111111111100000",
61299 => "0111111111100000",
61300 => "0111111111100000",
61301 => "0111111111100000",
61302 => "0111111111100000",
61303 => "0111111111100000",
61304 => "0111111111100000",
61305 => "0111111111100000",
61306 => "0111111111100000",
61307 => "0111111111100000",
61308 => "0111111111100000",
61309 => "0111111111100000",
61310 => "0111111111100000",
61311 => "0111111111100000",
61312 => "0111111111100000",
61313 => "0111111111100000",
61314 => "0111111111100000",
61315 => "0111111111100000",
61316 => "0111111111100000",
61317 => "0111111111100000",
61318 => "0111111111100000",
61319 => "0111111111100000",
61320 => "0111111111100000",
61321 => "0111111111100000",
61322 => "0111111111100000",
61323 => "0111111111100000",
61324 => "0111111111100000",
61325 => "0111111111100000",
61326 => "0111111111100000",
61327 => "0111111111100000",
61328 => "0111111111100000",
61329 => "0111111111100000",
61330 => "0111111111100000",
61331 => "0111111111100000",
61332 => "0111111111100000",
61333 => "0111111111100000",
61334 => "0111111111100000",
61335 => "0111111111100000",
61336 => "0111111111100000",
61337 => "0111111111100000",
61338 => "0111111111100000",
61339 => "0111111111100000",
61340 => "0111111111100000",
61341 => "0111111111100000",
61342 => "0111111111100000",
61343 => "0111111111100000",
61344 => "0111111111100000",
61345 => "0111111111100000",
61346 => "0111111111100000",
61347 => "0111111111100000",
61348 => "0111111111100000",
61349 => "0111111111100000",
61350 => "0111111111100000",
61351 => "0111111111100000",
61352 => "0111111111100000",
61353 => "0111111111100000",
61354 => "0111111111100000",
61355 => "0111111111100000",
61356 => "0111111111100000",
61357 => "0111111111100000",
61358 => "0111111111100000",
61359 => "0111111111100000",
61360 => "0111111111100000",
61361 => "0111111111100000",
61362 => "0111111111100000",
61363 => "0111111111100000",
61364 => "0111111111100000",
61365 => "0111111111100000",
61366 => "0111111111100000",
61367 => "0111111111100000",
61368 => "0111111111100000",
61369 => "0111111111100000",
61370 => "0111111111100000",
61371 => "0111111111100000",
61372 => "0111111111100000",
61373 => "0111111111100000",
61374 => "0111111111100000",
61375 => "0111111111100000",
61376 => "0111111111100000",
61377 => "0111111111100000",
61378 => "0111111111100000",
61379 => "0111111111100000",
61380 => "0111111111100000",
61381 => "0111111111100000",
61382 => "0111111111100000",
61383 => "0111111111100000",
61384 => "0111111111100000",
61385 => "0111111111100000",
61386 => "0111111111100000",
61387 => "0111111111100000",
61388 => "0111111111100000",
61389 => "0111111111100000",
61390 => "0111111111100000",
61391 => "0111111111100000",
61392 => "0111111111100000",
61393 => "0111111111100000",
61394 => "0111111111100000",
61395 => "0111111111100000",
61396 => "0111111111100000",
61397 => "0111111111100000",
61398 => "0111111111100000",
61399 => "0111111111100000",
61400 => "0111111111100000",
61401 => "0111111111100000",
61402 => "0111111111100000",
61403 => "0111111111100000",
61404 => "0111111111100000",
61405 => "0111111111100000",
61406 => "0111111111100000",
61407 => "0111111111100000",
61408 => "0111111111100000",
61409 => "0111111111100000",
61410 => "0111111111100000",
61411 => "0111111111100000",
61412 => "0111111111100000",
61413 => "0111111111100000",
61414 => "0111111111100000",
61415 => "0111111111100000",
61416 => "0111111111100000",
61417 => "0111111111100000",
61418 => "0111111111100000",
61419 => "0111111111100000",
61420 => "0111111111100000",
61421 => "0111111111100000",
61422 => "0111111111100000",
61423 => "0111111111100000",
61424 => "0111111111100000",
61425 => "0111111111100000",
61426 => "0111111111100000",
61427 => "0111111111100000",
61428 => "0111111111100000",
61429 => "0111111111100000",
61430 => "0111111111100000",
61431 => "0111111111100000",
61432 => "0111111111100000",
61433 => "0111111111100000",
61434 => "0111111111100000",
61435 => "0111111111100000",
61436 => "0111111111100000",
61437 => "0111111111100000",
61438 => "0111111111100000",
61439 => "0111111111100000",
61440 => "0111111111100000",
61441 => "0111111111100000",
61442 => "0111111111100000",
61443 => "0111111111100000",
61444 => "0111111111100000",
61445 => "0111111111100000",
61446 => "0111111111100000",
61447 => "0111111111100000",
61448 => "0111111111100000",
61449 => "0111111111100000",
61450 => "0111111111100000",
61451 => "0111111111100000",
61452 => "0111111111100000",
61453 => "0111111111100000",
61454 => "0111111111100000",
61455 => "0111111111100000",
61456 => "0111111111100000",
61457 => "0111111111100000",
61458 => "0111111111100000",
61459 => "0111111111100000",
61460 => "0111111111100000",
61461 => "0111111111100000",
61462 => "0111111111100000",
61463 => "0111111111100000",
61464 => "0111111111100000",
61465 => "0111111111100000",
61466 => "0111111111100000",
61467 => "0111111111100000",
61468 => "0111111111100000",
61469 => "0111111111100000",
61470 => "0111111111100000",
61471 => "0111111111100000",
61472 => "0111111111100000",
61473 => "0111111111100000",
61474 => "0111111111100000",
61475 => "0111111111100000",
61476 => "0111111111100000",
61477 => "0111111111100000",
61478 => "0111111111100000",
61479 => "0111111111100000",
61480 => "0111111111100000",
61481 => "0111111111100000",
61482 => "0111111111100000",
61483 => "0111111111100000",
61484 => "0111111111100000",
61485 => "0111111111100000",
61486 => "0111111111100000",
61487 => "0111111111100000",
61488 => "0111111111100000",
61489 => "0111111111100000",
61490 => "0111111111100000",
61491 => "0111111111100000",
61492 => "0111111111100000",
61493 => "0111111111100000",
61494 => "0111111111100000",
61495 => "0111111111100000",
61496 => "0111111111100000",
61497 => "0111111111100000",
61498 => "0111111111100000",
61499 => "0111111111100000",
61500 => "0111111111100000",
61501 => "0111111111100000",
61502 => "0111111111100000",
61503 => "0111111111100000",
61504 => "0111111111100000",
61505 => "0111111111100000",
61506 => "0111111111100000",
61507 => "0111111111100000",
61508 => "0111111111100000",
61509 => "0111111111100000",
61510 => "0111111111100000",
61511 => "0111111111100000",
61512 => "0111111111100000",
61513 => "0111111111100000",
61514 => "0111111111100000",
61515 => "0111111111100000",
61516 => "0111111111100000",
61517 => "0111111111100000",
61518 => "0111111111100000",
61519 => "0111111111100000",
61520 => "0111111111100000",
61521 => "0111111111100000",
61522 => "0111111111100000",
61523 => "0111111111100000",
61524 => "0111111111100000",
61525 => "0111111111100000",
61526 => "0111111111100000",
61527 => "0111111111100000",
61528 => "0111111111100000",
61529 => "0111111111100000",
61530 => "0111111111100000",
61531 => "0111111111100000",
61532 => "0111111111100000",
61533 => "0111111111100000",
61534 => "0111111111100000",
61535 => "0111111111100000",
61536 => "0111111111100000",
61537 => "0111111111100000",
61538 => "0111111111100000",
61539 => "0111111111100000",
61540 => "0111111111100000",
61541 => "0111111111100000",
61542 => "0111111111100000",
61543 => "0111111111100000",
61544 => "0111111111100000",
61545 => "0111111111100000",
61546 => "0111111111100000",
61547 => "0111111111100000",
61548 => "0111111111100000",
61549 => "0111111111100000",
61550 => "0111111111100000",
61551 => "0111111111100000",
61552 => "0111111111100000",
61553 => "0111111111100000",
61554 => "0111111111100000",
61555 => "0111111111100000",
61556 => "0111111111100000",
61557 => "0111111111100000",
61558 => "0111111111100000",
61559 => "0111111111100000",
61560 => "0111111111100000",
61561 => "0111111111100000",
61562 => "0111111111100000",
61563 => "0111111111100000",
61564 => "0111111111100000",
61565 => "0111111111100000",
61566 => "0111111111100000",
61567 => "0111111111100000",
61568 => "0111111111100000",
61569 => "0111111111100000",
61570 => "0111111111100000",
61571 => "0111111111100000",
61572 => "0111111111100000",
61573 => "0111111111100000",
61574 => "0111111111100000",
61575 => "0111111111100000",
61576 => "0111111111100000",
61577 => "0111111111100000",
61578 => "0111111111100000",
61579 => "0111111111100000",
61580 => "0111111111100000",
61581 => "0111111111100000",
61582 => "0111111111100000",
61583 => "0111111111100000",
61584 => "0111111111100000",
61585 => "0111111111100000",
61586 => "0111111111100000",
61587 => "0111111111100000",
61588 => "0111111111100000",
61589 => "0111111111100000",
61590 => "0111111111100000",
61591 => "0111111111100000",
61592 => "0111111111100000",
61593 => "0111111111100000",
61594 => "0111111111100000",
61595 => "0111111111100000",
61596 => "0111111111100000",
61597 => "0111111111100000",
61598 => "0111111111100000",
61599 => "0111111111100000",
61600 => "0111111111100000",
61601 => "0111111111100000",
61602 => "0111111111100000",
61603 => "0111111111100000",
61604 => "0111111111100000",
61605 => "0111111111100000",
61606 => "0111111111100000",
61607 => "0111111111100000",
61608 => "0111111111100000",
61609 => "0111111111100000",
61610 => "0111111111100000",
61611 => "0111111111100000",
61612 => "0111111111100000",
61613 => "0111111111100000",
61614 => "0111111111100000",
61615 => "0111111111100000",
61616 => "0111111111100000",
61617 => "0111111111100000",
61618 => "0111111111100000",
61619 => "0111111111100000",
61620 => "0111111111100000",
61621 => "0111111111100000",
61622 => "0111111111100000",
61623 => "0111111111100000",
61624 => "0111111111100000",
61625 => "0111111111100000",
61626 => "0111111111100000",
61627 => "0111111111100000",
61628 => "0111111111100000",
61629 => "0111111111100000",
61630 => "0111111111100000",
61631 => "0111111111100000",
61632 => "0111111111100000",
61633 => "0111111111100000",
61634 => "0111111111100000",
61635 => "0111111111100000",
61636 => "0111111111100000",
61637 => "0111111111100000",
61638 => "0111111111100000",
61639 => "0111111111100000",
61640 => "0111111111100000",
61641 => "0111111111100000",
61642 => "0111111111100000",
61643 => "0111111111100000",
61644 => "0111111111100000",
61645 => "0111111111100000",
61646 => "0111111111100000",
61647 => "0111111111100000",
61648 => "0111111111100000",
61649 => "0111111111100000",
61650 => "0111111111100000",
61651 => "0111111111100000",
61652 => "0111111111100000",
61653 => "0111111111100000",
61654 => "0111111111100000",
61655 => "0111111111100000",
61656 => "0111111111100000",
61657 => "0111111111100000",
61658 => "0111111111100000",
61659 => "0111111111100000",
61660 => "0111111111100000",
61661 => "0111111111100000",
61662 => "0111111111100000",
61663 => "0111111111100000",
61664 => "0111111111100000",
61665 => "0111111111100000",
61666 => "0111111111100000",
61667 => "0111111111100000",
61668 => "0111111111100000",
61669 => "0111111111100000",
61670 => "0111111111100000",
61671 => "0111111111100000",
61672 => "0111111111100000",
61673 => "0111111111100000",
61674 => "0111111111100000",
61675 => "0111111111100000",
61676 => "0111111111100000",
61677 => "0111111111100000",
61678 => "0111111111100000",
61679 => "0111111111100000",
61680 => "0111111111100000",
61681 => "0111111111100000",
61682 => "0111111111100000",
61683 => "0111111111100000",
61684 => "0111111111100000",
61685 => "0111111111100000",
61686 => "0111111111100000",
61687 => "0111111111100000",
61688 => "0111111111100000",
61689 => "0111111111100000",
61690 => "0111111111100000",
61691 => "0111111111100000",
61692 => "0111111111100000",
61693 => "0111111111100000",
61694 => "0111111111100000",
61695 => "0111111111100000",
61696 => "0111111111100000",
61697 => "0111111111100000",
61698 => "0111111111100000",
61699 => "0111111111100000",
61700 => "0111111111100000",
61701 => "0111111111100000",
61702 => "0111111111100000",
61703 => "0111111111100000",
61704 => "0111111111100000",
61705 => "0111111111100000",
61706 => "0111111111100000",
61707 => "0111111111100000",
61708 => "0111111111100000",
61709 => "0111111111100000",
61710 => "0111111111100000",
61711 => "0111111111100000",
61712 => "0111111111100000",
61713 => "0111111111100000",
61714 => "0111111111100000",
61715 => "0111111111100000",
61716 => "0111111111100000",
61717 => "0111111111100000",
61718 => "0111111111100000",
61719 => "0111111111100000",
61720 => "0111111111100000",
61721 => "0111111111100000",
61722 => "0111111111100000",
61723 => "0111111111100000",
61724 => "0111111111100000",
61725 => "0111111111100000",
61726 => "0111111111100000",
61727 => "0111111111100000",
61728 => "0111111111100000",
61729 => "0111111111100000",
61730 => "0111111111100000",
61731 => "0111111111100000",
61732 => "0111111111100000",
61733 => "0111111111100000",
61734 => "0111111111100000",
61735 => "0111111111100000",
61736 => "0111111111100000",
61737 => "0111111111100000",
61738 => "0111111111100000",
61739 => "0111111111100000",
61740 => "0111111111100000",
61741 => "0111111111100000",
61742 => "0111111111100000",
61743 => "0111111111100000",
61744 => "0111111111100000",
61745 => "0111111111100000",
61746 => "0111111111100000",
61747 => "0111111111100000",
61748 => "0111111111100000",
61749 => "0111111111100000",
61750 => "0111111111100000",
61751 => "0111111111100000",
61752 => "0111111111100000",
61753 => "0111111111100000",
61754 => "0111111111100000",
61755 => "0111111111100000",
61756 => "0111111111100000",
61757 => "0111111111100000",
61758 => "0111111111100000",
61759 => "0111111111100000",
61760 => "0111111111100000",
61761 => "0111111111100000",
61762 => "0111111111100000",
61763 => "0111111111100000",
61764 => "0111111111100000",
61765 => "0111111111100000",
61766 => "0111111111100000",
61767 => "0111111111100000",
61768 => "0111111111100000",
61769 => "0111111111100000",
61770 => "0111111111100000",
61771 => "0111111111100000",
61772 => "0111111111100000",
61773 => "0111111111100000",
61774 => "0111111111100000",
61775 => "0111111111100000",
61776 => "0111111111100000",
61777 => "0111111111100000",
61778 => "0111111111100000",
61779 => "0111111111100000",
61780 => "0111111111100000",
61781 => "0111111111100000",
61782 => "0111111111100000",
61783 => "0111111111100000",
61784 => "0111111111100000",
61785 => "0111111111100000",
61786 => "0111111111100000",
61787 => "0111111111100000",
61788 => "0111111111100000",
61789 => "0111111111100000",
61790 => "0111111111100000",
61791 => "0111111111100000",
61792 => "0111111111100000",
61793 => "0111111111100000",
61794 => "0111111111100000",
61795 => "0111111111100000",
61796 => "0111111111100000",
61797 => "0111111111100000",
61798 => "0111111111100000",
61799 => "0111111111100000",
61800 => "0111111111100000",
61801 => "0111111111100000",
61802 => "0111111111100000",
61803 => "0111111111100000",
61804 => "0111111111100000",
61805 => "0111111111100000",
61806 => "0111111111100000",
61807 => "0111111111100000",
61808 => "0111111111100000",
61809 => "0111111111100000",
61810 => "0111111111100000",
61811 => "0111111111100000",
61812 => "0111111111100000",
61813 => "0111111111100000",
61814 => "0111111111100000",
61815 => "0111111111100000",
61816 => "0111111111100000",
61817 => "0111111111100000",
61818 => "0111111111100000",
61819 => "0111111111100000",
61820 => "0111111111100000",
61821 => "0111111111100000",
61822 => "0111111111100000",
61823 => "0111111111100000",
61824 => "0111111111100000",
61825 => "0111111111100000",
61826 => "0111111111100000",
61827 => "0111111111100000",
61828 => "0111111111100000",
61829 => "0111111111100000",
61830 => "0111111111100000",
61831 => "0111111111100000",
61832 => "0111111111100000",
61833 => "0111111111100000",
61834 => "0111111111100000",
61835 => "0111111111100000",
61836 => "0111111111100000",
61837 => "0111111111100000",
61838 => "0111111111100000",
61839 => "0111111111100000",
61840 => "0111111111100000",
61841 => "0111111111100000",
61842 => "0111111111100000",
61843 => "0111111111100000",
61844 => "0111111111100000",
61845 => "0111111111100000",
61846 => "0111111111100000",
61847 => "0111111111100000",
61848 => "0111111111100000",
61849 => "0111111111100000",
61850 => "0111111111100000",
61851 => "0111111111100000",
61852 => "0111111111100000",
61853 => "0111111111100000",
61854 => "0111111111100000",
61855 => "0111111111100000",
61856 => "0111111111100000",
61857 => "0111111111100000",
61858 => "0111111111100000",
61859 => "0111111111100000",
61860 => "0111111111100000",
61861 => "0111111111100000",
61862 => "0111111111100000",
61863 => "0111111111100000",
61864 => "0111111111100000",
61865 => "0111111111100000",
61866 => "0111111111100000",
61867 => "0111111111100000",
61868 => "0111111111100000",
61869 => "0111111111100000",
61870 => "0111111111100000",
61871 => "0111111111100000",
61872 => "0111111111100000",
61873 => "0111111111100000",
61874 => "0111111111100000",
61875 => "0111111111100000",
61876 => "0111111111100000",
61877 => "0111111111100000",
61878 => "0111111111100000",
61879 => "0111111111100000",
61880 => "0111111111100000",
61881 => "0111111111100000",
61882 => "0111111111100000",
61883 => "0111111111100000",
61884 => "0111111111100000",
61885 => "0111111111100000",
61886 => "0111111111100000",
61887 => "0111111111100000",
61888 => "0111111111100000",
61889 => "0111111111100000",
61890 => "0111111111100000",
61891 => "0111111111100000",
61892 => "0111111111100000",
61893 => "0111111111100000",
61894 => "0111111111100000",
61895 => "0111111111100000",
61896 => "0111111111100000",
61897 => "0111111111100000",
61898 => "0111111111100000",
61899 => "0111111111100000",
61900 => "0111111111100000",
61901 => "0111111111100000",
61902 => "0111111111100000",
61903 => "0111111111100000",
61904 => "0111111111100000",
61905 => "0111111111100000",
61906 => "0111111111100000",
61907 => "0111111111100000",
61908 => "0111111111100000",
61909 => "0111111111100000",
61910 => "0111111111100000",
61911 => "0111111111100000",
61912 => "0111111111100000",
61913 => "0111111111100000",
61914 => "0111111111100000",
61915 => "0111111111100000",
61916 => "0111111111100000",
61917 => "0111111111100000",
61918 => "0111111111100000",
61919 => "0111111111100000",
61920 => "0111111111100000",
61921 => "0111111111100000",
61922 => "0111111111100000",
61923 => "0111111111100000",
61924 => "0111111111100000",
61925 => "0111111111100000",
61926 => "0111111111100000",
61927 => "0111111111100000",
61928 => "0111111111100000",
61929 => "0111111111100000",
61930 => "0111111111100000",
61931 => "0111111111100000",
61932 => "0111111111100000",
61933 => "0111111111100000",
61934 => "0111111111100000",
61935 => "0111111111100000",
61936 => "0111111111100000",
61937 => "0111111111100000",
61938 => "0111111111100000",
61939 => "0111111111100000",
61940 => "0111111111100000",
61941 => "0111111111100000",
61942 => "0111111111100000",
61943 => "0111111111100000",
61944 => "0111111111100000",
61945 => "0111111111100000",
61946 => "0111111111100000",
61947 => "0111111111100000",
61948 => "0111111111100000",
61949 => "0111111111100000",
61950 => "0111111111100000",
61951 => "0111111111100000",
61952 => "0111111111100000",
61953 => "0111111111100000",
61954 => "0111111111100000",
61955 => "0111111111100000",
61956 => "0111111111100000",
61957 => "0111111111100000",
61958 => "0111111111100000",
61959 => "0111111111100000",
61960 => "0111111111100000",
61961 => "0111111111100000",
61962 => "0111111111100000",
61963 => "0111111111100000",
61964 => "0111111111100000",
61965 => "0111111111100000",
61966 => "0111111111100000",
61967 => "0111111111100000",
61968 => "0111111111100000",
61969 => "0111111111100000",
61970 => "0111111111100000",
61971 => "0111111111100000",
61972 => "0111111111100000",
61973 => "0111111111100000",
61974 => "0111111111100000",
61975 => "0111111111100000",
61976 => "0111111111100000",
61977 => "0111111111100000",
61978 => "0111111111100000",
61979 => "0111111111100000",
61980 => "0111111111100000",
61981 => "0111111111100000",
61982 => "0111111111100000",
61983 => "0111111111100000",
61984 => "0111111111100000",
61985 => "0111111111100000",
61986 => "0111111111100000",
61987 => "0111111111100000",
61988 => "0111111111100000",
61989 => "0111111111100000",
61990 => "0111111111100000",
61991 => "0111111111100000",
61992 => "0111111111100000",
61993 => "0111111111100000",
61994 => "0111111111100000",
61995 => "0111111111100000",
61996 => "0111111111100000",
61997 => "0111111111100000",
61998 => "0111111111100000",
61999 => "0111111111100000",
62000 => "0111111111100000",
62001 => "0111111111100000",
62002 => "0111111111100000",
62003 => "0111111111100000",
62004 => "0111111111100000",
62005 => "0111111111100000",
62006 => "0111111111100000",
62007 => "0111111111100000",
62008 => "0111111111100000",
62009 => "0111111111100000",
62010 => "0111111111100000",
62011 => "0111111111100000",
62012 => "0111111111100000",
62013 => "0111111111100000",
62014 => "0111111111100000",
62015 => "0111111111100000",
62016 => "0111111111100000",
62017 => "0111111111100000",
62018 => "0111111111100000",
62019 => "0111111111100000",
62020 => "0111111111100000",
62021 => "0111111111100000",
62022 => "0111111111100000",
62023 => "0111111111100000",
62024 => "0111111111100000",
62025 => "0111111111100000",
62026 => "0111111111100000",
62027 => "0111111111100000",
62028 => "0111111111100000",
62029 => "0111111111100000",
62030 => "0111111111100000",
62031 => "0111111111100000",
62032 => "0111111111100000",
62033 => "0111111111100000",
62034 => "0111111111100000",
62035 => "0111111111100000",
62036 => "0111111111100000",
62037 => "0111111111100000",
62038 => "0111111111100000",
62039 => "0111111111100000",
62040 => "0111111111100000",
62041 => "0111111111100000",
62042 => "0111111111100000",
62043 => "0111111111100000",
62044 => "0111111111100000",
62045 => "0111111111100000",
62046 => "0111111111100000",
62047 => "0111111111100000",
62048 => "0111111111100000",
62049 => "0111111111100000",
62050 => "0111111111100000",
62051 => "0111111111100000",
62052 => "0111111111100000",
62053 => "0111111111100000",
62054 => "0111111111100000",
62055 => "0111111111100000",
62056 => "0111111111100000",
62057 => "0111111111100000",
62058 => "0111111111100000",
62059 => "0111111111100000",
62060 => "0111111111100000",
62061 => "0111111111100000",
62062 => "0111111111100000",
62063 => "0111111111100000",
62064 => "0111111111100000",
62065 => "0111111111100000",
62066 => "0111111111100000",
62067 => "0111111111100000",
62068 => "0111111111100000",
62069 => "0111111111100000",
62070 => "0111111111100000",
62071 => "0111111111100000",
62072 => "0111111111100000",
62073 => "0111111111100000",
62074 => "0111111111100000",
62075 => "0111111111100000",
62076 => "0111111111100000",
62077 => "0111111111100000",
62078 => "0111111111100000",
62079 => "0111111111100000",
62080 => "0111111111100000",
62081 => "0111111111100000",
62082 => "0111111111100000",
62083 => "0111111111100000",
62084 => "0111111111100000",
62085 => "0111111111100000",
62086 => "0111111111100000",
62087 => "0111111111100000",
62088 => "0111111111100000",
62089 => "0111111111100000",
62090 => "0111111111100000",
62091 => "0111111111100000",
62092 => "0111111111100000",
62093 => "0111111111100000",
62094 => "0111111111100000",
62095 => "0111111111100000",
62096 => "0111111111100000",
62097 => "0111111111100000",
62098 => "0111111111100000",
62099 => "0111111111100000",
62100 => "0111111111100000",
62101 => "0111111111100000",
62102 => "0111111111100000",
62103 => "0111111111100000",
62104 => "0111111111100000",
62105 => "0111111111100000",
62106 => "0111111111100000",
62107 => "0111111111100000",
62108 => "0111111111100000",
62109 => "0111111111100000",
62110 => "0111111111100000",
62111 => "0111111111100000",
62112 => "0111111111100000",
62113 => "0111111111100000",
62114 => "0111111111100000",
62115 => "0111111111100000",
62116 => "0111111111100000",
62117 => "0111111111100000",
62118 => "0111111111100000",
62119 => "0111111111100000",
62120 => "0111111111100000",
62121 => "0111111111100000",
62122 => "0111111111100000",
62123 => "0111111111100000",
62124 => "0111111111100000",
62125 => "0111111111100000",
62126 => "0111111111100000",
62127 => "0111111111100000",
62128 => "0111111111100000",
62129 => "0111111111100000",
62130 => "0111111111100000",
62131 => "0111111111100000",
62132 => "0111111111100000",
62133 => "0111111111100000",
62134 => "0111111111100000",
62135 => "0111111111100000",
62136 => "0111111111100000",
62137 => "0111111111100000",
62138 => "0111111111100000",
62139 => "0111111111100000",
62140 => "0111111111100000",
62141 => "0111111111100000",
62142 => "0111111111100000",
62143 => "0111111111100000",
62144 => "0111111111100000",
62145 => "0111111111100000",
62146 => "0111111111100000",
62147 => "0111111111100000",
62148 => "0111111111100000",
62149 => "0111111111100000",
62150 => "0111111111100000",
62151 => "0111111111100000",
62152 => "0111111111100000",
62153 => "0111111111100000",
62154 => "0111111111100000",
62155 => "0111111111100000",
62156 => "0111111111100000",
62157 => "0111111111100000",
62158 => "0111111111100000",
62159 => "0111111111100000",
62160 => "0111111111100000",
62161 => "0111111111100000",
62162 => "0111111111100000",
62163 => "0111111111100000",
62164 => "0111111111100000",
62165 => "0111111111100000",
62166 => "0111111111100000",
62167 => "0111111111100000",
62168 => "0111111111100000",
62169 => "0111111111100000",
62170 => "0111111111100000",
62171 => "0111111111100000",
62172 => "0111111111100000",
62173 => "0111111111100000",
62174 => "0111111111100000",
62175 => "0111111111100000",
62176 => "0111111111100000",
62177 => "0111111111100000",
62178 => "0111111111100000",
62179 => "0111111111100000",
62180 => "0111111111100000",
62181 => "0111111111100000",
62182 => "0111111111100000",
62183 => "0111111111100000",
62184 => "0111111111100000",
62185 => "0111111111100000",
62186 => "0111111111100000",
62187 => "0111111111100000",
62188 => "0111111111100000",
62189 => "0111111111100000",
62190 => "0111111111100000",
62191 => "0111111111100000",
62192 => "0111111111100000",
62193 => "0111111111100000",
62194 => "0111111111100000",
62195 => "0111111111100000",
62196 => "0111111111100000",
62197 => "0111111111100000",
62198 => "0111111111100000",
62199 => "0111111111100000",
62200 => "0111111111100000",
62201 => "0111111111100000",
62202 => "0111111111100000",
62203 => "0111111111100000",
62204 => "0111111111100000",
62205 => "0111111111100000",
62206 => "0111111111100000",
62207 => "0111111111100000",
62208 => "0111111111100000",
62209 => "0111111111100000",
62210 => "0111111111100000",
62211 => "0111111111100000",
62212 => "0111111111100000",
62213 => "0111111111100000",
62214 => "0111111111100000",
62215 => "0111111111100000",
62216 => "0111111111100000",
62217 => "0111111111100000",
62218 => "0111111111100000",
62219 => "0111111111100000",
62220 => "0111111111100000",
62221 => "0111111111100000",
62222 => "0111111111100000",
62223 => "0111111111100000",
62224 => "0111111111100000",
62225 => "0111111111100000",
62226 => "0111111111100000",
62227 => "0111111111100000",
62228 => "0111111111100000",
62229 => "0111111111100000",
62230 => "0111111111100000",
62231 => "0111111111100000",
62232 => "0111111111100000",
62233 => "0111111111100000",
62234 => "0111111111100000",
62235 => "0111111111100000",
62236 => "0111111111100000",
62237 => "0111111111100000",
62238 => "0111111111100000",
62239 => "0111111111100000",
62240 => "0111111111100000",
62241 => "0111111111100000",
62242 => "0111111111100000",
62243 => "0111111111100000",
62244 => "0111111111100000",
62245 => "0111111111100000",
62246 => "0111111111100000",
62247 => "0111111111100000",
62248 => "0111111111100000",
62249 => "0111111111100000",
62250 => "0111111111100000",
62251 => "0111111111100000",
62252 => "0111111111100000",
62253 => "0111111111100000",
62254 => "0111111111100000",
62255 => "0111111111100000",
62256 => "0111111111100000",
62257 => "0111111111100000",
62258 => "0111111111100000",
62259 => "0111111111100000",
62260 => "0111111111100000",
62261 => "0111111111100000",
62262 => "0111111111100000",
62263 => "0111111111100000",
62264 => "0111111111100000",
62265 => "0111111111100000",
62266 => "0111111111100000",
62267 => "0111111111100000",
62268 => "0111111111100000",
62269 => "0111111111100000",
62270 => "0111111111100000",
62271 => "0111111111100000",
62272 => "0111111111100000",
62273 => "0111111111100000",
62274 => "0111111111100000",
62275 => "0111111111100000",
62276 => "0111111111100000",
62277 => "0111111111100000",
62278 => "0111111111100000",
62279 => "0111111111100000",
62280 => "0111111111100000",
62281 => "0111111111100000",
62282 => "0111111111100000",
62283 => "0111111111100000",
62284 => "0111111111100000",
62285 => "0111111111100000",
62286 => "0111111111100000",
62287 => "0111111111100000",
62288 => "0111111111100000",
62289 => "0111111111100000",
62290 => "0111111111100000",
62291 => "0111111111100000",
62292 => "0111111111100000",
62293 => "0111111111100000",
62294 => "0111111111100000",
62295 => "0111111111100000",
62296 => "0111111111100000",
62297 => "0111111111100000",
62298 => "0111111111100000",
62299 => "0111111111100000",
62300 => "0111111111100000",
62301 => "0111111111100000",
62302 => "0111111111100000",
62303 => "0111111111100000",
62304 => "0111111111100000",
62305 => "0111111111100000",
62306 => "0111111111100000",
62307 => "0111111111100000",
62308 => "0111111111100000",
62309 => "0111111111100000",
62310 => "0111111111100000",
62311 => "0111111111100000",
62312 => "0111111111100000",
62313 => "0111111111100000",
62314 => "0111111111100000",
62315 => "0111111111100000",
62316 => "0111111111100000",
62317 => "0111111111100000",
62318 => "0111111111100000",
62319 => "0111111111100000",
62320 => "0111111111100000",
62321 => "0111111111100000",
62322 => "0111111111100000",
62323 => "0111111111100000",
62324 => "0111111111100000",
62325 => "0111111111100000",
62326 => "0111111111100000",
62327 => "0111111111100000",
62328 => "0111111111100000",
62329 => "0111111111100000",
62330 => "0111111111100000",
62331 => "0111111111100000",
62332 => "0111111111100000",
62333 => "0111111111100000",
62334 => "0111111111110000",
62335 => "0111111111110000",
62336 => "0111111111110000",
62337 => "0111111111110000",
62338 => "0111111111110000",
62339 => "0111111111110000",
62340 => "0111111111110000",
62341 => "0111111111110000",
62342 => "0111111111110000",
62343 => "0111111111110000",
62344 => "0111111111110000",
62345 => "0111111111110000",
62346 => "0111111111110000",
62347 => "0111111111110000",
62348 => "0111111111110000",
62349 => "0111111111110000",
62350 => "0111111111110000",
62351 => "0111111111110000",
62352 => "0111111111110000",
62353 => "0111111111110000",
62354 => "0111111111110000",
62355 => "0111111111110000",
62356 => "0111111111110000",
62357 => "0111111111110000",
62358 => "0111111111110000",
62359 => "0111111111110000",
62360 => "0111111111110000",
62361 => "0111111111110000",
62362 => "0111111111110000",
62363 => "0111111111110000",
62364 => "0111111111110000",
62365 => "0111111111110000",
62366 => "0111111111110000",
62367 => "0111111111110000",
62368 => "0111111111110000",
62369 => "0111111111110000",
62370 => "0111111111110000",
62371 => "0111111111110000",
62372 => "0111111111110000",
62373 => "0111111111110000",
62374 => "0111111111110000",
62375 => "0111111111110000",
62376 => "0111111111110000",
62377 => "0111111111110000",
62378 => "0111111111110000",
62379 => "0111111111110000",
62380 => "0111111111110000",
62381 => "0111111111110000",
62382 => "0111111111110000",
62383 => "0111111111110000",
62384 => "0111111111110000",
62385 => "0111111111110000",
62386 => "0111111111110000",
62387 => "0111111111110000",
62388 => "0111111111110000",
62389 => "0111111111110000",
62390 => "0111111111110000",
62391 => "0111111111110000",
62392 => "0111111111110000",
62393 => "0111111111110000",
62394 => "0111111111110000",
62395 => "0111111111110000",
62396 => "0111111111110000",
62397 => "0111111111110000",
62398 => "0111111111110000",
62399 => "0111111111110000",
62400 => "0111111111110000",
62401 => "0111111111110000",
62402 => "0111111111110000",
62403 => "0111111111110000",
62404 => "0111111111110000",
62405 => "0111111111110000",
62406 => "0111111111110000",
62407 => "0111111111110000",
62408 => "0111111111110000",
62409 => "0111111111110000",
62410 => "0111111111110000",
62411 => "0111111111110000",
62412 => "0111111111110000",
62413 => "0111111111110000",
62414 => "0111111111110000",
62415 => "0111111111110000",
62416 => "0111111111110000",
62417 => "0111111111110000",
62418 => "0111111111110000",
62419 => "0111111111110000",
62420 => "0111111111110000",
62421 => "0111111111110000",
62422 => "0111111111110000",
62423 => "0111111111110000",
62424 => "0111111111110000",
62425 => "0111111111110000",
62426 => "0111111111110000",
62427 => "0111111111110000",
62428 => "0111111111110000",
62429 => "0111111111110000",
62430 => "0111111111110000",
62431 => "0111111111110000",
62432 => "0111111111110000",
62433 => "0111111111110000",
62434 => "0111111111110000",
62435 => "0111111111110000",
62436 => "0111111111110000",
62437 => "0111111111110000",
62438 => "0111111111110000",
62439 => "0111111111110000",
62440 => "0111111111110000",
62441 => "0111111111110000",
62442 => "0111111111110000",
62443 => "0111111111110000",
62444 => "0111111111110000",
62445 => "0111111111110000",
62446 => "0111111111110000",
62447 => "0111111111110000",
62448 => "0111111111110000",
62449 => "0111111111110000",
62450 => "0111111111110000",
62451 => "0111111111110000",
62452 => "0111111111110000",
62453 => "0111111111110000",
62454 => "0111111111110000",
62455 => "0111111111110000",
62456 => "0111111111110000",
62457 => "0111111111110000",
62458 => "0111111111110000",
62459 => "0111111111110000",
62460 => "0111111111110000",
62461 => "0111111111110000",
62462 => "0111111111110000",
62463 => "0111111111110000",
62464 => "0111111111110000",
62465 => "0111111111110000",
62466 => "0111111111110000",
62467 => "0111111111110000",
62468 => "0111111111110000",
62469 => "0111111111110000",
62470 => "0111111111110000",
62471 => "0111111111110000",
62472 => "0111111111110000",
62473 => "0111111111110000",
62474 => "0111111111110000",
62475 => "0111111111110000",
62476 => "0111111111110000",
62477 => "0111111111110000",
62478 => "0111111111110000",
62479 => "0111111111110000",
62480 => "0111111111110000",
62481 => "0111111111110000",
62482 => "0111111111110000",
62483 => "0111111111110000",
62484 => "0111111111110000",
62485 => "0111111111110000",
62486 => "0111111111110000",
62487 => "0111111111110000",
62488 => "0111111111110000",
62489 => "0111111111110000",
62490 => "0111111111110000",
62491 => "0111111111110000",
62492 => "0111111111110000",
62493 => "0111111111110000",
62494 => "0111111111110000",
62495 => "0111111111110000",
62496 => "0111111111110000",
62497 => "0111111111110000",
62498 => "0111111111110000",
62499 => "0111111111110000",
62500 => "0111111111110000",
62501 => "0111111111110000",
62502 => "0111111111110000",
62503 => "0111111111110000",
62504 => "0111111111110000",
62505 => "0111111111110000",
62506 => "0111111111110000",
62507 => "0111111111110000",
62508 => "0111111111110000",
62509 => "0111111111110000",
62510 => "0111111111110000",
62511 => "0111111111110000",
62512 => "0111111111110000",
62513 => "0111111111110000",
62514 => "0111111111110000",
62515 => "0111111111110000",
62516 => "0111111111110000",
62517 => "0111111111110000",
62518 => "0111111111110000",
62519 => "0111111111110000",
62520 => "0111111111110000",
62521 => "0111111111110000",
62522 => "0111111111110000",
62523 => "0111111111110000",
62524 => "0111111111110000",
62525 => "0111111111110000",
62526 => "0111111111110000",
62527 => "0111111111110000",
62528 => "0111111111110000",
62529 => "0111111111110000",
62530 => "0111111111110000",
62531 => "0111111111110000",
62532 => "0111111111110000",
62533 => "0111111111110000",
62534 => "0111111111110000",
62535 => "0111111111110000",
62536 => "0111111111110000",
62537 => "0111111111110000",
62538 => "0111111111110000",
62539 => "0111111111110000",
62540 => "0111111111110000",
62541 => "0111111111110000",
62542 => "0111111111110000",
62543 => "0111111111110000",
62544 => "0111111111110000",
62545 => "0111111111110000",
62546 => "0111111111110000",
62547 => "0111111111110000",
62548 => "0111111111110000",
62549 => "0111111111110000",
62550 => "0111111111110000",
62551 => "0111111111110000",
62552 => "0111111111110000",
62553 => "0111111111110000",
62554 => "0111111111110000",
62555 => "0111111111110000",
62556 => "0111111111110000",
62557 => "0111111111110000",
62558 => "0111111111110000",
62559 => "0111111111110000",
62560 => "0111111111110000",
62561 => "0111111111110000",
62562 => "0111111111110000",
62563 => "0111111111110000",
62564 => "0111111111110000",
62565 => "0111111111110000",
62566 => "0111111111110000",
62567 => "0111111111110000",
62568 => "0111111111110000",
62569 => "0111111111110000",
62570 => "0111111111110000",
62571 => "0111111111110000",
62572 => "0111111111110000",
62573 => "0111111111110000",
62574 => "0111111111110000",
62575 => "0111111111110000",
62576 => "0111111111110000",
62577 => "0111111111110000",
62578 => "0111111111110000",
62579 => "0111111111110000",
62580 => "0111111111110000",
62581 => "0111111111110000",
62582 => "0111111111110000",
62583 => "0111111111110000",
62584 => "0111111111110000",
62585 => "0111111111110000",
62586 => "0111111111110000",
62587 => "0111111111110000",
62588 => "0111111111110000",
62589 => "0111111111110000",
62590 => "0111111111110000",
62591 => "0111111111110000",
62592 => "0111111111110000",
62593 => "0111111111110000",
62594 => "0111111111110000",
62595 => "0111111111110000",
62596 => "0111111111110000",
62597 => "0111111111110000",
62598 => "0111111111110000",
62599 => "0111111111110000",
62600 => "0111111111110000",
62601 => "0111111111110000",
62602 => "0111111111110000",
62603 => "0111111111110000",
62604 => "0111111111110000",
62605 => "0111111111110000",
62606 => "0111111111110000",
62607 => "0111111111110000",
62608 => "0111111111110000",
62609 => "0111111111110000",
62610 => "0111111111110000",
62611 => "0111111111110000",
62612 => "0111111111110000",
62613 => "0111111111110000",
62614 => "0111111111110000",
62615 => "0111111111110000",
62616 => "0111111111110000",
62617 => "0111111111110000",
62618 => "0111111111110000",
62619 => "0111111111110000",
62620 => "0111111111110000",
62621 => "0111111111110000",
62622 => "0111111111110000",
62623 => "0111111111110000",
62624 => "0111111111110000",
62625 => "0111111111110000",
62626 => "0111111111110000",
62627 => "0111111111110000",
62628 => "0111111111110000",
62629 => "0111111111110000",
62630 => "0111111111110000",
62631 => "0111111111110000",
62632 => "0111111111110000",
62633 => "0111111111110000",
62634 => "0111111111110000",
62635 => "0111111111110000",
62636 => "0111111111110000",
62637 => "0111111111110000",
62638 => "0111111111110000",
62639 => "0111111111110000",
62640 => "0111111111110000",
62641 => "0111111111110000",
62642 => "0111111111110000",
62643 => "0111111111110000",
62644 => "0111111111110000",
62645 => "0111111111110000",
62646 => "0111111111110000",
62647 => "0111111111110000",
62648 => "0111111111110000",
62649 => "0111111111110000",
62650 => "0111111111110000",
62651 => "0111111111110000",
62652 => "0111111111110000",
62653 => "0111111111110000",
62654 => "0111111111110000",
62655 => "0111111111110000",
62656 => "0111111111110000",
62657 => "0111111111110000",
62658 => "0111111111110000",
62659 => "0111111111110000",
62660 => "0111111111110000",
62661 => "0111111111110000",
62662 => "0111111111110000",
62663 => "0111111111110000",
62664 => "0111111111110000",
62665 => "0111111111110000",
62666 => "0111111111110000",
62667 => "0111111111110000",
62668 => "0111111111110000",
62669 => "0111111111110000",
62670 => "0111111111110000",
62671 => "0111111111110000",
62672 => "0111111111110000",
62673 => "0111111111110000",
62674 => "0111111111110000",
62675 => "0111111111110000",
62676 => "0111111111110000",
62677 => "0111111111110000",
62678 => "0111111111110000",
62679 => "0111111111110000",
62680 => "0111111111110000",
62681 => "0111111111110000",
62682 => "0111111111110000",
62683 => "0111111111110000",
62684 => "0111111111110000",
62685 => "0111111111110000",
62686 => "0111111111110000",
62687 => "0111111111110000",
62688 => "0111111111110000",
62689 => "0111111111110000",
62690 => "0111111111110000",
62691 => "0111111111110000",
62692 => "0111111111110000",
62693 => "0111111111110000",
62694 => "0111111111110000",
62695 => "0111111111110000",
62696 => "0111111111110000",
62697 => "0111111111110000",
62698 => "0111111111110000",
62699 => "0111111111110000",
62700 => "0111111111110000",
62701 => "0111111111110000",
62702 => "0111111111110000",
62703 => "0111111111110000",
62704 => "0111111111110000",
62705 => "0111111111110000",
62706 => "0111111111110000",
62707 => "0111111111110000",
62708 => "0111111111110000",
62709 => "0111111111110000",
62710 => "0111111111110000",
62711 => "0111111111110000",
62712 => "0111111111110000",
62713 => "0111111111110000",
62714 => "0111111111110000",
62715 => "0111111111110000",
62716 => "0111111111110000",
62717 => "0111111111110000",
62718 => "0111111111110000",
62719 => "0111111111110000",
62720 => "0111111111110000",
62721 => "0111111111110000",
62722 => "0111111111110000",
62723 => "0111111111110000",
62724 => "0111111111110000",
62725 => "0111111111110000",
62726 => "0111111111110000",
62727 => "0111111111110000",
62728 => "0111111111110000",
62729 => "0111111111110000",
62730 => "0111111111110000",
62731 => "0111111111110000",
62732 => "0111111111110000",
62733 => "0111111111110000",
62734 => "0111111111110000",
62735 => "0111111111110000",
62736 => "0111111111110000",
62737 => "0111111111110000",
62738 => "0111111111110000",
62739 => "0111111111110000",
62740 => "0111111111110000",
62741 => "0111111111110000",
62742 => "0111111111110000",
62743 => "0111111111110000",
62744 => "0111111111110000",
62745 => "0111111111110000",
62746 => "0111111111110000",
62747 => "0111111111110000",
62748 => "0111111111110000",
62749 => "0111111111110000",
62750 => "0111111111110000",
62751 => "0111111111110000",
62752 => "0111111111110000",
62753 => "0111111111110000",
62754 => "0111111111110000",
62755 => "0111111111110000",
62756 => "0111111111110000",
62757 => "0111111111110000",
62758 => "0111111111110000",
62759 => "0111111111110000",
62760 => "0111111111110000",
62761 => "0111111111110000",
62762 => "0111111111110000",
62763 => "0111111111110000",
62764 => "0111111111110000",
62765 => "0111111111110000",
62766 => "0111111111110000",
62767 => "0111111111110000",
62768 => "0111111111110000",
62769 => "0111111111110000",
62770 => "0111111111110000",
62771 => "0111111111110000",
62772 => "0111111111110000",
62773 => "0111111111110000",
62774 => "0111111111110000",
62775 => "0111111111110000",
62776 => "0111111111110000",
62777 => "0111111111110000",
62778 => "0111111111110000",
62779 => "0111111111110000",
62780 => "0111111111110000",
62781 => "0111111111110000",
62782 => "0111111111110000",
62783 => "0111111111110000",
62784 => "0111111111110000",
62785 => "0111111111110000",
62786 => "0111111111110000",
62787 => "0111111111110000",
62788 => "0111111111110000",
62789 => "0111111111110000",
62790 => "0111111111110000",
62791 => "0111111111110000",
62792 => "0111111111110000",
62793 => "0111111111110000",
62794 => "0111111111110000",
62795 => "0111111111110000",
62796 => "0111111111110000",
62797 => "0111111111110000",
62798 => "0111111111110000",
62799 => "0111111111110000",
62800 => "0111111111110000",
62801 => "0111111111110000",
62802 => "0111111111110000",
62803 => "0111111111110000",
62804 => "0111111111110000",
62805 => "0111111111110000",
62806 => "0111111111110000",
62807 => "0111111111110000",
62808 => "0111111111110000",
62809 => "0111111111110000",
62810 => "0111111111110000",
62811 => "0111111111110000",
62812 => "0111111111110000",
62813 => "0111111111110000",
62814 => "0111111111110000",
62815 => "0111111111110000",
62816 => "0111111111110000",
62817 => "0111111111110000",
62818 => "0111111111110000",
62819 => "0111111111110000",
62820 => "0111111111110000",
62821 => "0111111111110000",
62822 => "0111111111110000",
62823 => "0111111111110000",
62824 => "0111111111110000",
62825 => "0111111111110000",
62826 => "0111111111110000",
62827 => "0111111111110000",
62828 => "0111111111110000",
62829 => "0111111111110000",
62830 => "0111111111110000",
62831 => "0111111111110000",
62832 => "0111111111110000",
62833 => "0111111111110000",
62834 => "0111111111110000",
62835 => "0111111111110000",
62836 => "0111111111110000",
62837 => "0111111111110000",
62838 => "0111111111110000",
62839 => "0111111111110000",
62840 => "0111111111110000",
62841 => "0111111111110000",
62842 => "0111111111110000",
62843 => "0111111111110000",
62844 => "0111111111110000",
62845 => "0111111111110000",
62846 => "0111111111110000",
62847 => "0111111111110000",
62848 => "0111111111110000",
62849 => "0111111111110000",
62850 => "0111111111110000",
62851 => "0111111111110000",
62852 => "0111111111110000",
62853 => "0111111111110000",
62854 => "0111111111110000",
62855 => "0111111111110000",
62856 => "0111111111110000",
62857 => "0111111111110000",
62858 => "0111111111110000",
62859 => "0111111111110000",
62860 => "0111111111110000",
62861 => "0111111111110000",
62862 => "0111111111110000",
62863 => "0111111111110000",
62864 => "0111111111110000",
62865 => "0111111111110000",
62866 => "0111111111110000",
62867 => "0111111111110000",
62868 => "0111111111110000",
62869 => "0111111111110000",
62870 => "0111111111110000",
62871 => "0111111111110000",
62872 => "0111111111110000",
62873 => "0111111111110000",
62874 => "0111111111110000",
62875 => "0111111111110000",
62876 => "0111111111110000",
62877 => "0111111111110000",
62878 => "0111111111110000",
62879 => "0111111111110000",
62880 => "0111111111110000",
62881 => "0111111111110000",
62882 => "0111111111110000",
62883 => "0111111111110000",
62884 => "0111111111110000",
62885 => "0111111111110000",
62886 => "0111111111110000",
62887 => "0111111111110000",
62888 => "0111111111110000",
62889 => "0111111111110000",
62890 => "0111111111110000",
62891 => "0111111111110000",
62892 => "0111111111110000",
62893 => "0111111111110000",
62894 => "0111111111110000",
62895 => "0111111111110000",
62896 => "0111111111110000",
62897 => "0111111111110000",
62898 => "0111111111110000",
62899 => "0111111111110000",
62900 => "0111111111110000",
62901 => "0111111111110000",
62902 => "0111111111110000",
62903 => "0111111111110000",
62904 => "0111111111110000",
62905 => "0111111111110000",
62906 => "0111111111110000",
62907 => "0111111111110000",
62908 => "0111111111110000",
62909 => "0111111111110000",
62910 => "0111111111110000",
62911 => "0111111111110000",
62912 => "0111111111110000",
62913 => "0111111111110000",
62914 => "0111111111110000",
62915 => "0111111111110000",
62916 => "0111111111110000",
62917 => "0111111111110000",
62918 => "0111111111110000",
62919 => "0111111111110000",
62920 => "0111111111110000",
62921 => "0111111111110000",
62922 => "0111111111110000",
62923 => "0111111111110000",
62924 => "0111111111110000",
62925 => "0111111111110000",
62926 => "0111111111110000",
62927 => "0111111111110000",
62928 => "0111111111110000",
62929 => "0111111111110000",
62930 => "0111111111110000",
62931 => "0111111111110000",
62932 => "0111111111110000",
62933 => "0111111111110000",
62934 => "0111111111110000",
62935 => "0111111111110000",
62936 => "0111111111110000",
62937 => "0111111111110000",
62938 => "0111111111110000",
62939 => "0111111111110000",
62940 => "0111111111110000",
62941 => "0111111111110000",
62942 => "0111111111110000",
62943 => "0111111111110000",
62944 => "0111111111110000",
62945 => "0111111111110000",
62946 => "0111111111110000",
62947 => "0111111111110000",
62948 => "0111111111110000",
62949 => "0111111111110000",
62950 => "0111111111110000",
62951 => "0111111111110000",
62952 => "0111111111110000",
62953 => "0111111111110000",
62954 => "0111111111110000",
62955 => "0111111111110000",
62956 => "0111111111110000",
62957 => "0111111111110000",
62958 => "0111111111110000",
62959 => "0111111111110000",
62960 => "0111111111110000",
62961 => "0111111111110000",
62962 => "0111111111110000",
62963 => "0111111111110000",
62964 => "0111111111110000",
62965 => "0111111111110000",
62966 => "0111111111110000",
62967 => "0111111111110000",
62968 => "0111111111110000",
62969 => "0111111111110000",
62970 => "0111111111110000",
62971 => "0111111111110000",
62972 => "0111111111110000",
62973 => "0111111111110000",
62974 => "0111111111110000",
62975 => "0111111111110000",
62976 => "0111111111110000",
62977 => "0111111111110000",
62978 => "0111111111110000",
62979 => "0111111111110000",
62980 => "0111111111110000",
62981 => "0111111111110000",
62982 => "0111111111110000",
62983 => "0111111111110000",
62984 => "0111111111110000",
62985 => "0111111111110000",
62986 => "0111111111110000",
62987 => "0111111111110000",
62988 => "0111111111110000",
62989 => "0111111111110000",
62990 => "0111111111110000",
62991 => "0111111111110000",
62992 => "0111111111110000",
62993 => "0111111111110000",
62994 => "0111111111110000",
62995 => "0111111111110000",
62996 => "0111111111110000",
62997 => "0111111111110000",
62998 => "0111111111110000",
62999 => "0111111111110000",
63000 => "0111111111110000",
63001 => "0111111111110000",
63002 => "0111111111110000",
63003 => "0111111111110000",
63004 => "0111111111110000",
63005 => "0111111111110000",
63006 => "0111111111110000",
63007 => "0111111111110000",
63008 => "0111111111110000",
63009 => "0111111111110000",
63010 => "0111111111110000",
63011 => "0111111111110000",
63012 => "0111111111110000",
63013 => "0111111111110000",
63014 => "0111111111110000",
63015 => "0111111111110000",
63016 => "0111111111110000",
63017 => "0111111111110000",
63018 => "0111111111110000",
63019 => "0111111111110000",
63020 => "0111111111110000",
63021 => "0111111111110000",
63022 => "0111111111110000",
63023 => "0111111111110000",
63024 => "0111111111110000",
63025 => "0111111111110000",
63026 => "0111111111110000",
63027 => "0111111111110000",
63028 => "0111111111110000",
63029 => "0111111111110000",
63030 => "0111111111110000",
63031 => "0111111111110000",
63032 => "0111111111110000",
63033 => "0111111111110000",
63034 => "0111111111110000",
63035 => "0111111111110000",
63036 => "0111111111110000",
63037 => "0111111111110000",
63038 => "0111111111110000",
63039 => "0111111111110000",
63040 => "0111111111110000",
63041 => "0111111111110000",
63042 => "0111111111110000",
63043 => "0111111111110000",
63044 => "0111111111110000",
63045 => "0111111111110000",
63046 => "0111111111110000",
63047 => "0111111111110000",
63048 => "0111111111110000",
63049 => "0111111111110000",
63050 => "0111111111110000",
63051 => "0111111111110000",
63052 => "0111111111110000",
63053 => "0111111111110000",
63054 => "0111111111110000",
63055 => "0111111111110000",
63056 => "0111111111110000",
63057 => "0111111111110000",
63058 => "0111111111110000",
63059 => "0111111111110000",
63060 => "0111111111110000",
63061 => "0111111111110000",
63062 => "0111111111110000",
63063 => "0111111111110000",
63064 => "0111111111110000",
63065 => "0111111111110000",
63066 => "0111111111110000",
63067 => "0111111111110000",
63068 => "0111111111110000",
63069 => "0111111111110000",
63070 => "0111111111110000",
63071 => "0111111111110000",
63072 => "0111111111110000",
63073 => "0111111111110000",
63074 => "0111111111110000",
63075 => "0111111111110000",
63076 => "0111111111110000",
63077 => "0111111111110000",
63078 => "0111111111110000",
63079 => "0111111111110000",
63080 => "0111111111110000",
63081 => "0111111111110000",
63082 => "0111111111110000",
63083 => "0111111111110000",
63084 => "0111111111110000",
63085 => "0111111111110000",
63086 => "0111111111110000",
63087 => "0111111111110000",
63088 => "0111111111110000",
63089 => "0111111111110000",
63090 => "0111111111110000",
63091 => "0111111111110000",
63092 => "0111111111110000",
63093 => "0111111111110000",
63094 => "0111111111110000",
63095 => "0111111111110000",
63096 => "0111111111110000",
63097 => "0111111111110000",
63098 => "0111111111110000",
63099 => "0111111111110000",
63100 => "0111111111110000",
63101 => "0111111111110000",
63102 => "0111111111110000",
63103 => "0111111111110000",
63104 => "0111111111110000",
63105 => "0111111111110000",
63106 => "0111111111110000",
63107 => "0111111111110000",
63108 => "0111111111110000",
63109 => "0111111111110000",
63110 => "0111111111110000",
63111 => "0111111111110000",
63112 => "0111111111110000",
63113 => "0111111111110000",
63114 => "0111111111110000",
63115 => "0111111111110000",
63116 => "0111111111110000",
63117 => "0111111111110000",
63118 => "0111111111110000",
63119 => "0111111111110000",
63120 => "0111111111110000",
63121 => "0111111111110000",
63122 => "0111111111110000",
63123 => "0111111111110000",
63124 => "0111111111110000",
63125 => "0111111111110000",
63126 => "0111111111110000",
63127 => "0111111111110000",
63128 => "0111111111110000",
63129 => "0111111111110000",
63130 => "0111111111110000",
63131 => "0111111111110000",
63132 => "0111111111110000",
63133 => "0111111111110000",
63134 => "0111111111110000",
63135 => "0111111111110000",
63136 => "0111111111110000",
63137 => "0111111111110000",
63138 => "0111111111110000",
63139 => "0111111111110000",
63140 => "0111111111110000",
63141 => "0111111111110000",
63142 => "0111111111110000",
63143 => "0111111111110000",
63144 => "0111111111110000",
63145 => "0111111111110000",
63146 => "0111111111110000",
63147 => "0111111111110000",
63148 => "0111111111110000",
63149 => "0111111111110000",
63150 => "0111111111110000",
63151 => "0111111111110000",
63152 => "0111111111110000",
63153 => "0111111111110000",
63154 => "0111111111110000",
63155 => "0111111111110000",
63156 => "0111111111110000",
63157 => "0111111111110000",
63158 => "0111111111110000",
63159 => "0111111111110000",
63160 => "0111111111110000",
63161 => "0111111111110000",
63162 => "0111111111110000",
63163 => "0111111111110000",
63164 => "0111111111110000",
63165 => "0111111111110000",
63166 => "0111111111110000",
63167 => "0111111111110000",
63168 => "0111111111110000",
63169 => "0111111111110000",
63170 => "0111111111110000",
63171 => "0111111111110000",
63172 => "0111111111110000",
63173 => "0111111111110000",
63174 => "0111111111110000",
63175 => "0111111111110000",
63176 => "0111111111110000",
63177 => "0111111111110000",
63178 => "0111111111110000",
63179 => "0111111111110000",
63180 => "0111111111110000",
63181 => "0111111111110000",
63182 => "0111111111110000",
63183 => "0111111111110000",
63184 => "0111111111110000",
63185 => "0111111111110000",
63186 => "0111111111110000",
63187 => "0111111111110000",
63188 => "0111111111110000",
63189 => "0111111111110000",
63190 => "0111111111110000",
63191 => "0111111111110000",
63192 => "0111111111110000",
63193 => "0111111111110000",
63194 => "0111111111110000",
63195 => "0111111111110000",
63196 => "0111111111110000",
63197 => "0111111111110000",
63198 => "0111111111110000",
63199 => "0111111111110000",
63200 => "0111111111110000",
63201 => "0111111111110000",
63202 => "0111111111110000",
63203 => "0111111111110000",
63204 => "0111111111110000",
63205 => "0111111111110000",
63206 => "0111111111110000",
63207 => "0111111111110000",
63208 => "0111111111110000",
63209 => "0111111111110000",
63210 => "0111111111110000",
63211 => "0111111111110000",
63212 => "0111111111110000",
63213 => "0111111111110000",
63214 => "0111111111110000",
63215 => "0111111111110000",
63216 => "0111111111110000",
63217 => "0111111111110000",
63218 => "0111111111110000",
63219 => "0111111111110000",
63220 => "0111111111110000",
63221 => "0111111111110000",
63222 => "0111111111110000",
63223 => "0111111111110000",
63224 => "0111111111110000",
63225 => "0111111111110000",
63226 => "0111111111110000",
63227 => "0111111111110000",
63228 => "0111111111110000",
63229 => "0111111111110000",
63230 => "0111111111110000",
63231 => "0111111111110000",
63232 => "0111111111110000",
63233 => "0111111111110000",
63234 => "0111111111110000",
63235 => "0111111111110000",
63236 => "0111111111110000",
63237 => "0111111111110000",
63238 => "0111111111110000",
63239 => "0111111111110000",
63240 => "0111111111110000",
63241 => "0111111111110000",
63242 => "0111111111110000",
63243 => "0111111111110000",
63244 => "0111111111110000",
63245 => "0111111111110000",
63246 => "0111111111110000",
63247 => "0111111111110000",
63248 => "0111111111110000",
63249 => "0111111111110000",
63250 => "0111111111110000",
63251 => "0111111111110000",
63252 => "0111111111110000",
63253 => "0111111111110000",
63254 => "0111111111110000",
63255 => "0111111111110000",
63256 => "0111111111110000",
63257 => "0111111111110000",
63258 => "0111111111110000",
63259 => "0111111111110000",
63260 => "0111111111110000",
63261 => "0111111111110000",
63262 => "0111111111110000",
63263 => "0111111111110000",
63264 => "0111111111110000",
63265 => "0111111111110000",
63266 => "0111111111110000",
63267 => "0111111111110000",
63268 => "0111111111110000",
63269 => "0111111111110000",
63270 => "0111111111110000",
63271 => "0111111111110000",
63272 => "0111111111110000",
63273 => "0111111111110000",
63274 => "0111111111110000",
63275 => "0111111111110000",
63276 => "0111111111110000",
63277 => "0111111111110000",
63278 => "0111111111110000",
63279 => "0111111111110000",
63280 => "0111111111110000",
63281 => "0111111111110000",
63282 => "0111111111110000",
63283 => "0111111111110000",
63284 => "0111111111110000",
63285 => "0111111111110000",
63286 => "0111111111110000",
63287 => "0111111111110000",
63288 => "0111111111110000",
63289 => "0111111111110000",
63290 => "0111111111110000",
63291 => "0111111111110000",
63292 => "0111111111110000",
63293 => "0111111111110000",
63294 => "0111111111110000",
63295 => "0111111111110000",
63296 => "0111111111110000",
63297 => "0111111111110000",
63298 => "0111111111110000",
63299 => "0111111111110000",
63300 => "0111111111110000",
63301 => "0111111111110000",
63302 => "0111111111110000",
63303 => "0111111111110000",
63304 => "0111111111110000",
63305 => "0111111111110000",
63306 => "0111111111110000",
63307 => "0111111111110000",
63308 => "0111111111110000",
63309 => "0111111111110000",
63310 => "0111111111110000",
63311 => "0111111111110000",
63312 => "0111111111110000",
63313 => "0111111111110000",
63314 => "0111111111110000",
63315 => "0111111111110000",
63316 => "0111111111110000",
63317 => "0111111111110000",
63318 => "0111111111110000",
63319 => "0111111111110000",
63320 => "0111111111110000",
63321 => "0111111111110000",
63322 => "0111111111110000",
63323 => "0111111111110000",
63324 => "0111111111110000",
63325 => "0111111111110000",
63326 => "0111111111110000",
63327 => "0111111111110000",
63328 => "0111111111110000",
63329 => "0111111111110000",
63330 => "0111111111110000",
63331 => "0111111111110000",
63332 => "0111111111110000",
63333 => "0111111111110000",
63334 => "0111111111110000",
63335 => "0111111111110000",
63336 => "0111111111110000",
63337 => "0111111111110000",
63338 => "0111111111110000",
63339 => "0111111111110000",
63340 => "0111111111110000",
63341 => "0111111111110000",
63342 => "0111111111110000",
63343 => "0111111111110000",
63344 => "0111111111110000",
63345 => "0111111111110000",
63346 => "0111111111110000",
63347 => "0111111111110000",
63348 => "0111111111110000",
63349 => "0111111111110000",
63350 => "0111111111110000",
63351 => "0111111111110000",
63352 => "0111111111110000",
63353 => "0111111111110000",
63354 => "0111111111110000",
63355 => "0111111111110000",
63356 => "0111111111110000",
63357 => "0111111111110000",
63358 => "0111111111110000",
63359 => "0111111111110000",
63360 => "0111111111110000",
63361 => "0111111111110000",
63362 => "0111111111110000",
63363 => "0111111111110000",
63364 => "0111111111110000",
63365 => "0111111111110000",
63366 => "0111111111110000",
63367 => "0111111111110000",
63368 => "0111111111110000",
63369 => "0111111111110000",
63370 => "0111111111110000",
63371 => "0111111111110000",
63372 => "0111111111110000",
63373 => "0111111111110000",
63374 => "0111111111110000",
63375 => "0111111111110000",
63376 => "0111111111110000",
63377 => "0111111111110000",
63378 => "0111111111110000",
63379 => "0111111111110000",
63380 => "0111111111110000",
63381 => "0111111111110000",
63382 => "0111111111110000",
63383 => "0111111111110000",
63384 => "0111111111110000",
63385 => "0111111111110000",
63386 => "0111111111110000",
63387 => "0111111111110000",
63388 => "0111111111110000",
63389 => "0111111111110000",
63390 => "0111111111110000",
63391 => "0111111111110000",
63392 => "0111111111110000",
63393 => "0111111111110000",
63394 => "0111111111110000",
63395 => "0111111111110000",
63396 => "0111111111110000",
63397 => "0111111111110000",
63398 => "0111111111110000",
63399 => "0111111111110000",
63400 => "0111111111110000",
63401 => "0111111111110000",
63402 => "0111111111110000",
63403 => "0111111111110000",
63404 => "0111111111110000",
63405 => "0111111111110000",
63406 => "0111111111110000",
63407 => "0111111111110000",
63408 => "0111111111110000",
63409 => "0111111111110000",
63410 => "0111111111110000",
63411 => "0111111111110000",
63412 => "0111111111110000",
63413 => "0111111111110000",
63414 => "0111111111110000",
63415 => "0111111111110000",
63416 => "0111111111110000",
63417 => "0111111111110000",
63418 => "0111111111110000",
63419 => "0111111111110000",
63420 => "0111111111110000",
63421 => "0111111111110000",
63422 => "0111111111110000",
63423 => "0111111111110000",
63424 => "0111111111110000",
63425 => "0111111111110000",
63426 => "0111111111110000",
63427 => "0111111111110000",
63428 => "0111111111110000",
63429 => "0111111111110000",
63430 => "0111111111110000",
63431 => "0111111111110000",
63432 => "0111111111110000",
63433 => "0111111111110000",
63434 => "0111111111110000",
63435 => "0111111111110000",
63436 => "0111111111110000",
63437 => "0111111111110000",
63438 => "0111111111110000",
63439 => "0111111111110000",
63440 => "0111111111110000",
63441 => "0111111111110000",
63442 => "0111111111110000",
63443 => "0111111111110000",
63444 => "0111111111110000",
63445 => "0111111111110000",
63446 => "0111111111110000",
63447 => "0111111111110000",
63448 => "0111111111110000",
63449 => "0111111111110000",
63450 => "0111111111110000",
63451 => "0111111111110000",
63452 => "0111111111110000",
63453 => "0111111111110000",
63454 => "0111111111110000",
63455 => "0111111111110000",
63456 => "0111111111110000",
63457 => "0111111111110000",
63458 => "0111111111110000",
63459 => "0111111111110000",
63460 => "0111111111110000",
63461 => "0111111111110000",
63462 => "0111111111110000",
63463 => "0111111111110000",
63464 => "0111111111110000",
63465 => "0111111111110000",
63466 => "0111111111110000",
63467 => "0111111111110000",
63468 => "0111111111110000",
63469 => "0111111111110000",
63470 => "0111111111110000",
63471 => "0111111111110000",
63472 => "0111111111110000",
63473 => "0111111111110000",
63474 => "0111111111110000",
63475 => "0111111111110000",
63476 => "0111111111110000",
63477 => "0111111111110000",
63478 => "0111111111110000",
63479 => "0111111111110000",
63480 => "0111111111110000",
63481 => "0111111111110000",
63482 => "0111111111110000",
63483 => "0111111111110000",
63484 => "0111111111110000",
63485 => "0111111111110000",
63486 => "0111111111110000",
63487 => "0111111111110000",
63488 => "0111111111110000",
63489 => "0111111111110000",
63490 => "0111111111110000",
63491 => "0111111111110000",
63492 => "0111111111110000",
63493 => "0111111111110000",
63494 => "0111111111110000",
63495 => "0111111111110000",
63496 => "0111111111110000",
63497 => "0111111111110000",
63498 => "0111111111110000",
63499 => "0111111111110000",
63500 => "0111111111110000",
63501 => "0111111111110000",
63502 => "0111111111110000",
63503 => "0111111111110000",
63504 => "0111111111110000",
63505 => "0111111111110000",
63506 => "0111111111110000",
63507 => "0111111111110000",
63508 => "0111111111110000",
63509 => "0111111111110000",
63510 => "0111111111110000",
63511 => "0111111111110000",
63512 => "0111111111110000",
63513 => "0111111111110000",
63514 => "0111111111110000",
63515 => "0111111111110000",
63516 => "0111111111110000",
63517 => "0111111111110000",
63518 => "0111111111110000",
63519 => "0111111111110000",
63520 => "0111111111110000",
63521 => "0111111111110000",
63522 => "0111111111110000",
63523 => "0111111111110000",
63524 => "0111111111110000",
63525 => "0111111111110000",
63526 => "0111111111110000",
63527 => "0111111111110000",
63528 => "0111111111110000",
63529 => "0111111111110000",
63530 => "0111111111110000",
63531 => "0111111111110000",
63532 => "0111111111110000",
63533 => "0111111111110000",
63534 => "0111111111110000",
63535 => "0111111111110000",
63536 => "0111111111110000",
63537 => "0111111111110000",
63538 => "0111111111110000",
63539 => "0111111111110000",
63540 => "0111111111110000",
63541 => "0111111111110000",
63542 => "0111111111110000",
63543 => "0111111111110000",
63544 => "0111111111110000",
63545 => "0111111111110000",
63546 => "0111111111110000",
63547 => "0111111111110000",
63548 => "0111111111110000",
63549 => "0111111111110000",
63550 => "0111111111110000",
63551 => "0111111111110000",
63552 => "0111111111110000",
63553 => "0111111111110000",
63554 => "0111111111110000",
63555 => "0111111111110000",
63556 => "0111111111110000",
63557 => "0111111111110000",
63558 => "0111111111110000",
63559 => "0111111111110000",
63560 => "0111111111110000",
63561 => "0111111111110000",
63562 => "0111111111110000",
63563 => "0111111111110000",
63564 => "0111111111110000",
63565 => "0111111111110000",
63566 => "0111111111110000",
63567 => "0111111111110000",
63568 => "0111111111110000",
63569 => "0111111111110000",
63570 => "0111111111110000",
63571 => "0111111111110000",
63572 => "0111111111110000",
63573 => "0111111111110000",
63574 => "0111111111110000",
63575 => "0111111111110000",
63576 => "0111111111110000",
63577 => "0111111111110000",
63578 => "0111111111110000",
63579 => "0111111111110000",
63580 => "0111111111110000",
63581 => "0111111111110000",
63582 => "0111111111110000",
63583 => "0111111111110000",
63584 => "0111111111110000",
63585 => "0111111111110000",
63586 => "0111111111110000",
63587 => "0111111111110000",
63588 => "0111111111110000",
63589 => "0111111111110000",
63590 => "0111111111110000",
63591 => "0111111111110000",
63592 => "0111111111110000",
63593 => "0111111111110000",
63594 => "0111111111110000",
63595 => "0111111111110000",
63596 => "0111111111110000",
63597 => "0111111111110000",
63598 => "0111111111110000",
63599 => "0111111111110000",
63600 => "0111111111110000",
63601 => "0111111111110000",
63602 => "0111111111110000",
63603 => "0111111111110000",
63604 => "0111111111110000",
63605 => "0111111111110000",
63606 => "0111111111110000",
63607 => "0111111111110000",
63608 => "0111111111110000",
63609 => "0111111111110000",
63610 => "0111111111110000",
63611 => "0111111111110000",
63612 => "0111111111110000",
63613 => "0111111111110000",
63614 => "0111111111110000",
63615 => "0111111111110000",
63616 => "0111111111110000",
63617 => "0111111111110000",
63618 => "0111111111110000",
63619 => "0111111111110000",
63620 => "0111111111110000",
63621 => "0111111111110000",
63622 => "0111111111110000",
63623 => "0111111111110000",
63624 => "0111111111110000",
63625 => "0111111111110000",
63626 => "0111111111110000",
63627 => "0111111111110000",
63628 => "0111111111110000",
63629 => "0111111111110000",
63630 => "0111111111110000",
63631 => "0111111111110000",
63632 => "0111111111110000",
63633 => "0111111111110000",
63634 => "0111111111110000",
63635 => "0111111111110000",
63636 => "0111111111110000",
63637 => "0111111111110000",
63638 => "0111111111110000",
63639 => "0111111111110000",
63640 => "0111111111110000",
63641 => "0111111111110000",
63642 => "0111111111110000",
63643 => "0111111111110000",
63644 => "0111111111110000",
63645 => "0111111111110000",
63646 => "0111111111110000",
63647 => "0111111111110000",
63648 => "0111111111110000",
63649 => "0111111111110000",
63650 => "0111111111110000",
63651 => "0111111111110000",
63652 => "0111111111110000",
63653 => "0111111111110000",
63654 => "0111111111110000",
63655 => "0111111111110000",
63656 => "0111111111110000",
63657 => "0111111111110000",
63658 => "0111111111110000",
63659 => "0111111111110000",
63660 => "0111111111110000",
63661 => "0111111111110000",
63662 => "0111111111110000",
63663 => "0111111111110000",
63664 => "0111111111110000",
63665 => "0111111111110000",
63666 => "0111111111110000",
63667 => "0111111111110000",
63668 => "0111111111110000",
63669 => "0111111111110000",
63670 => "0111111111110000",
63671 => "0111111111110000",
63672 => "0111111111110000",
63673 => "0111111111110000",
63674 => "0111111111110000",
63675 => "0111111111110000",
63676 => "0111111111110000",
63677 => "0111111111110000",
63678 => "0111111111110000",
63679 => "0111111111110000",
63680 => "0111111111110000",
63681 => "0111111111110000",
63682 => "0111111111110000",
63683 => "0111111111110000",
63684 => "0111111111110000",
63685 => "0111111111110000",
63686 => "0111111111110000",
63687 => "0111111111110000",
63688 => "0111111111110000",
63689 => "0111111111110000",
63690 => "0111111111110000",
63691 => "0111111111110000",
63692 => "0111111111110000",
63693 => "0111111111110000",
63694 => "0111111111110000",
63695 => "0111111111110000",
63696 => "0111111111110000",
63697 => "0111111111110000",
63698 => "0111111111110000",
63699 => "0111111111110000",
63700 => "0111111111110000",
63701 => "0111111111110000",
63702 => "0111111111110000",
63703 => "0111111111110000",
63704 => "0111111111110000",
63705 => "0111111111110000",
63706 => "0111111111110000",
63707 => "0111111111110000",
63708 => "0111111111110000",
63709 => "0111111111110000",
63710 => "0111111111110000",
63711 => "0111111111110000",
63712 => "0111111111110000",
63713 => "0111111111110000",
63714 => "0111111111110000",
63715 => "0111111111110000",
63716 => "0111111111110000",
63717 => "0111111111110000",
63718 => "0111111111110000",
63719 => "0111111111110000",
63720 => "0111111111110000",
63721 => "0111111111110000",
63722 => "0111111111110000",
63723 => "0111111111110000",
63724 => "0111111111110000",
63725 => "0111111111110000",
63726 => "0111111111110000",
63727 => "0111111111110000",
63728 => "0111111111110000",
63729 => "0111111111110000",
63730 => "0111111111110000",
63731 => "0111111111110000",
63732 => "0111111111110000",
63733 => "0111111111110000",
63734 => "0111111111110000",
63735 => "0111111111110000",
63736 => "0111111111110000",
63737 => "0111111111110000",
63738 => "0111111111110000",
63739 => "0111111111110000",
63740 => "0111111111110000",
63741 => "0111111111110000",
63742 => "0111111111110000",
63743 => "0111111111110000",
63744 => "0111111111110000",
63745 => "0111111111110000",
63746 => "0111111111110000",
63747 => "0111111111110000",
63748 => "0111111111110000",
63749 => "0111111111110000",
63750 => "0111111111110000",
63751 => "0111111111110000",
63752 => "0111111111110000",
63753 => "0111111111110000",
63754 => "0111111111110000",
63755 => "0111111111110000",
63756 => "0111111111110000",
63757 => "0111111111110000",
63758 => "0111111111110000",
63759 => "0111111111110000",
63760 => "0111111111110000",
63761 => "0111111111110000",
63762 => "0111111111110000",
63763 => "0111111111110000",
63764 => "0111111111110000",
63765 => "0111111111110000",
63766 => "0111111111110000",
63767 => "0111111111110000",
63768 => "0111111111110000",
63769 => "0111111111110000",
63770 => "0111111111110000",
63771 => "0111111111110000",
63772 => "0111111111110000",
63773 => "0111111111110000",
63774 => "0111111111110000",
63775 => "0111111111110000",
63776 => "0111111111110000",
63777 => "0111111111110000",
63778 => "0111111111110000",
63779 => "0111111111110000",
63780 => "0111111111110000",
63781 => "0111111111110000",
63782 => "0111111111110000",
63783 => "0111111111110000",
63784 => "0111111111110000",
63785 => "0111111111110000",
63786 => "0111111111110000",
63787 => "0111111111110000",
63788 => "0111111111110000",
63789 => "0111111111110000",
63790 => "0111111111110000",
63791 => "0111111111110000",
63792 => "0111111111110000",
63793 => "0111111111110000",
63794 => "0111111111110000",
63795 => "0111111111110000",
63796 => "0111111111110000",
63797 => "0111111111110000",
63798 => "0111111111110000",
63799 => "0111111111110000",
63800 => "0111111111110000",
63801 => "0111111111110000",
63802 => "0111111111110000",
63803 => "0111111111110000",
63804 => "0111111111110000",
63805 => "0111111111110000",
63806 => "0111111111110000",
63807 => "0111111111110000",
63808 => "0111111111110000",
63809 => "0111111111110000",
63810 => "0111111111110000",
63811 => "0111111111110000",
63812 => "0111111111110000",
63813 => "0111111111110000",
63814 => "0111111111110000",
63815 => "0111111111110000",
63816 => "0111111111110000",
63817 => "0111111111110000",
63818 => "0111111111110000",
63819 => "0111111111110000",
63820 => "0111111111110000",
63821 => "0111111111110000",
63822 => "0111111111110000",
63823 => "0111111111110000",
63824 => "0111111111110000",
63825 => "0111111111110000",
63826 => "0111111111110000",
63827 => "0111111111110000",
63828 => "0111111111110000",
63829 => "0111111111110000",
63830 => "0111111111110000",
63831 => "0111111111110000",
63832 => "0111111111110000",
63833 => "0111111111110000",
63834 => "0111111111110000",
63835 => "0111111111110000",
63836 => "0111111111110000",
63837 => "0111111111110000",
63838 => "0111111111110000",
63839 => "0111111111110000",
63840 => "0111111111110000",
63841 => "0111111111110000",
63842 => "0111111111110000",
63843 => "0111111111110000",
63844 => "0111111111110000",
63845 => "0111111111110000",
63846 => "0111111111110000",
63847 => "0111111111110000",
63848 => "0111111111110000",
63849 => "0111111111110000",
63850 => "0111111111110000",
63851 => "0111111111110000",
63852 => "0111111111110000",
63853 => "0111111111110000",
63854 => "0111111111110000",
63855 => "0111111111110000",
63856 => "0111111111110000",
63857 => "0111111111110000",
63858 => "0111111111110000",
63859 => "0111111111110000",
63860 => "0111111111110000",
63861 => "0111111111110000",
63862 => "0111111111110000",
63863 => "0111111111110000",
63864 => "0111111111110000",
63865 => "0111111111110000",
63866 => "0111111111110000",
63867 => "0111111111110000",
63868 => "0111111111110000",
63869 => "0111111111110000",
63870 => "0111111111110000",
63871 => "0111111111110000",
63872 => "0111111111110000",
63873 => "0111111111110000",
63874 => "0111111111110000",
63875 => "0111111111110000",
63876 => "0111111111110000",
63877 => "0111111111110000",
63878 => "0111111111110000",
63879 => "0111111111110000",
63880 => "0111111111110000",
63881 => "0111111111110000",
63882 => "0111111111110000",
63883 => "0111111111110000",
63884 => "0111111111110000",
63885 => "0111111111110000",
63886 => "0111111111110000",
63887 => "0111111111110000",
63888 => "0111111111110000",
63889 => "0111111111110000",
63890 => "0111111111110000",
63891 => "0111111111110000",
63892 => "0111111111110000",
63893 => "0111111111110000",
63894 => "0111111111110000",
63895 => "0111111111110000",
63896 => "0111111111110000",
63897 => "0111111111110000",
63898 => "0111111111110000",
63899 => "0111111111110000",
63900 => "0111111111110000",
63901 => "0111111111110000",
63902 => "0111111111110000",
63903 => "0111111111110000",
63904 => "0111111111110000",
63905 => "0111111111110000",
63906 => "0111111111110000",
63907 => "0111111111110000",
63908 => "0111111111110000",
63909 => "0111111111110000",
63910 => "0111111111110000",
63911 => "0111111111110000",
63912 => "0111111111110000",
63913 => "0111111111110000",
63914 => "0111111111110000",
63915 => "0111111111110000",
63916 => "0111111111110000",
63917 => "0111111111110000",
63918 => "0111111111110000",
63919 => "0111111111110000",
63920 => "0111111111110000",
63921 => "0111111111110000",
63922 => "0111111111110000",
63923 => "0111111111110000",
63924 => "0111111111110000",
63925 => "0111111111110000",
63926 => "0111111111110000",
63927 => "0111111111110000",
63928 => "0111111111110000",
63929 => "0111111111110000",
63930 => "0111111111110000",
63931 => "0111111111110000",
63932 => "0111111111110000",
63933 => "0111111111110000",
63934 => "0111111111110000",
63935 => "0111111111110000",
63936 => "0111111111110000",
63937 => "0111111111110000",
63938 => "0111111111110000",
63939 => "0111111111110000",
63940 => "0111111111110000",
63941 => "0111111111110000",
63942 => "0111111111110000",
63943 => "0111111111110000",
63944 => "0111111111110000",
63945 => "0111111111110000",
63946 => "0111111111110000",
63947 => "0111111111110000",
63948 => "0111111111110000",
63949 => "0111111111110000",
63950 => "0111111111110000",
63951 => "0111111111110000",
63952 => "0111111111110000",
63953 => "0111111111110000",
63954 => "0111111111110000",
63955 => "0111111111110000",
63956 => "0111111111110000",
63957 => "0111111111110000",
63958 => "0111111111110000",
63959 => "0111111111110000",
63960 => "0111111111110000",
63961 => "0111111111110000",
63962 => "0111111111110000",
63963 => "0111111111110000",
63964 => "0111111111110000",
63965 => "0111111111110000",
63966 => "0111111111110000",
63967 => "0111111111110000",
63968 => "0111111111110000",
63969 => "0111111111110000",
63970 => "0111111111110000",
63971 => "0111111111110000",
63972 => "0111111111110000",
63973 => "0111111111110000",
63974 => "0111111111110000",
63975 => "0111111111110000",
63976 => "0111111111110000",
63977 => "0111111111110000",
63978 => "0111111111110000",
63979 => "0111111111110000",
63980 => "0111111111110000",
63981 => "0111111111110000",
63982 => "0111111111110000",
63983 => "0111111111110000",
63984 => "0111111111110000",
63985 => "0111111111110000",
63986 => "0111111111110000",
63987 => "0111111111110000",
63988 => "0111111111110000",
63989 => "0111111111110000",
63990 => "0111111111110000",
63991 => "0111111111110000",
63992 => "0111111111110000",
63993 => "0111111111110000",
63994 => "0111111111110000",
63995 => "0111111111110000",
63996 => "0111111111110000",
63997 => "0111111111110000",
63998 => "0111111111110000",
63999 => "0111111111110000",
64000 => "0111111111110000",
64001 => "0111111111110000",
64002 => "0111111111110000",
64003 => "0111111111110000",
64004 => "0111111111110000",
64005 => "0111111111110000",
64006 => "0111111111110000",
64007 => "0111111111110000",
64008 => "0111111111110000",
64009 => "0111111111110000",
64010 => "0111111111110000",
64011 => "0111111111110000",
64012 => "0111111111110000",
64013 => "0111111111110000",
64014 => "0111111111110000",
64015 => "0111111111110000",
64016 => "0111111111110000",
64017 => "0111111111110000",
64018 => "0111111111110000",
64019 => "0111111111110000",
64020 => "0111111111110000",
64021 => "0111111111110000",
64022 => "0111111111110000",
64023 => "0111111111110000",
64024 => "0111111111110000",
64025 => "0111111111110000",
64026 => "0111111111110000",
64027 => "0111111111110000",
64028 => "0111111111110000",
64029 => "0111111111110000",
64030 => "0111111111110000",
64031 => "0111111111110000",
64032 => "0111111111110000",
64033 => "0111111111110000",
64034 => "0111111111110000",
64035 => "0111111111110000",
64036 => "0111111111110000",
64037 => "0111111111110000",
64038 => "0111111111110000",
64039 => "0111111111110000",
64040 => "0111111111110000",
64041 => "0111111111110000",
64042 => "0111111111110000",
64043 => "0111111111110000",
64044 => "0111111111110000",
64045 => "0111111111110000",
64046 => "0111111111110000",
64047 => "0111111111110000",
64048 => "0111111111110000",
64049 => "0111111111110000",
64050 => "0111111111110000",
64051 => "0111111111110000",
64052 => "0111111111110000",
64053 => "0111111111110000",
64054 => "0111111111110000",
64055 => "0111111111110000",
64056 => "0111111111110000",
64057 => "0111111111110000",
64058 => "0111111111110000",
64059 => "0111111111110000",
64060 => "0111111111110000",
64061 => "0111111111110000",
64062 => "0111111111110000",
64063 => "0111111111110000",
64064 => "0111111111110000",
64065 => "0111111111110000",
64066 => "0111111111110000",
64067 => "0111111111110000",
64068 => "0111111111110000",
64069 => "0111111111110000",
64070 => "0111111111110000",
64071 => "0111111111110000",
64072 => "0111111111110000",
64073 => "0111111111110000",
64074 => "0111111111110000",
64075 => "0111111111110000",
64076 => "0111111111110000",
64077 => "0111111111110000",
64078 => "0111111111110000",
64079 => "0111111111110000",
64080 => "0111111111110000",
64081 => "0111111111110000",
64082 => "0111111111110000",
64083 => "0111111111110000",
64084 => "0111111111110000",
64085 => "0111111111110000",
64086 => "0111111111110000",
64087 => "0111111111110000",
64088 => "0111111111110000",
64089 => "0111111111110000",
64090 => "0111111111110000",
64091 => "0111111111110000",
64092 => "0111111111110000",
64093 => "0111111111110000",
64094 => "0111111111110000",
64095 => "0111111111110000",
64096 => "0111111111110000",
64097 => "0111111111110000",
64098 => "0111111111110000",
64099 => "0111111111110000",
64100 => "0111111111110000",
64101 => "0111111111110000",
64102 => "0111111111110000",
64103 => "0111111111110000",
64104 => "0111111111110000",
64105 => "0111111111110000",
64106 => "0111111111110000",
64107 => "0111111111110000",
64108 => "0111111111110000",
64109 => "0111111111110000",
64110 => "0111111111110000",
64111 => "0111111111110000",
64112 => "0111111111110000",
64113 => "0111111111110000",
64114 => "0111111111110000",
64115 => "0111111111110000",
64116 => "0111111111110000",
64117 => "0111111111110000",
64118 => "0111111111110000",
64119 => "0111111111110000",
64120 => "0111111111110000",
64121 => "0111111111110000",
64122 => "0111111111110000",
64123 => "0111111111110000",
64124 => "0111111111110000",
64125 => "0111111111110000",
64126 => "0111111111110000",
64127 => "0111111111110000",
64128 => "0111111111110000",
64129 => "0111111111110000",
64130 => "0111111111110000",
64131 => "0111111111110000",
64132 => "0111111111110000",
64133 => "0111111111110000",
64134 => "0111111111110000",
64135 => "0111111111110000",
64136 => "0111111111110000",
64137 => "0111111111110000",
64138 => "0111111111110000",
64139 => "0111111111110000",
64140 => "0111111111110000",
64141 => "0111111111110000",
64142 => "0111111111110000",
64143 => "0111111111110000",
64144 => "0111111111110000",
64145 => "0111111111110000",
64146 => "0111111111110000",
64147 => "0111111111110000",
64148 => "0111111111110000",
64149 => "0111111111110000",
64150 => "0111111111110000",
64151 => "0111111111110000",
64152 => "0111111111110000",
64153 => "0111111111110000",
64154 => "0111111111110000",
64155 => "0111111111110000",
64156 => "0111111111110000",
64157 => "0111111111110000",
64158 => "0111111111110000",
64159 => "0111111111110000",
64160 => "0111111111110000",
64161 => "0111111111110000",
64162 => "0111111111110000",
64163 => "0111111111110000",
64164 => "0111111111110000",
64165 => "0111111111110000",
64166 => "0111111111110000",
64167 => "0111111111110000",
64168 => "0111111111110000",
64169 => "0111111111110000",
64170 => "0111111111110000",
64171 => "0111111111110000",
64172 => "0111111111110000",
64173 => "0111111111110000",
64174 => "0111111111110000",
64175 => "0111111111110000",
64176 => "0111111111110000",
64177 => "0111111111110000",
64178 => "0111111111110000",
64179 => "0111111111110000",
64180 => "0111111111110000",
64181 => "0111111111110000",
64182 => "0111111111110000",
64183 => "0111111111110000",
64184 => "0111111111110000",
64185 => "0111111111110000",
64186 => "0111111111110000",
64187 => "0111111111110000",
64188 => "0111111111110000",
64189 => "0111111111110000",
64190 => "0111111111110000",
64191 => "0111111111110000",
64192 => "0111111111110000",
64193 => "0111111111110000",
64194 => "0111111111110000",
64195 => "0111111111110000",
64196 => "0111111111110000",
64197 => "0111111111110000",
64198 => "0111111111110000",
64199 => "0111111111110000",
64200 => "0111111111110000",
64201 => "0111111111110000",
64202 => "0111111111110000",
64203 => "0111111111110000",
64204 => "0111111111110000",
64205 => "0111111111110000",
64206 => "0111111111110000",
64207 => "0111111111110000",
64208 => "0111111111110000",
64209 => "0111111111110000",
64210 => "0111111111110000",
64211 => "0111111111110000",
64212 => "0111111111110000",
64213 => "0111111111110000",
64214 => "0111111111110000",
64215 => "0111111111110000",
64216 => "0111111111110000",
64217 => "0111111111110000",
64218 => "0111111111110000",
64219 => "0111111111110000",
64220 => "0111111111110000",
64221 => "0111111111110000",
64222 => "0111111111110000",
64223 => "0111111111110000",
64224 => "0111111111110000",
64225 => "0111111111110000",
64226 => "0111111111110000",
64227 => "0111111111110000",
64228 => "0111111111110000",
64229 => "0111111111110000",
64230 => "0111111111110000",
64231 => "0111111111110000",
64232 => "0111111111110000",
64233 => "0111111111110000",
64234 => "0111111111110000",
64235 => "0111111111110000",
64236 => "0111111111110000",
64237 => "0111111111110000",
64238 => "0111111111110000",
64239 => "0111111111110000",
64240 => "0111111111110000",
64241 => "0111111111110000",
64242 => "0111111111110000",
64243 => "0111111111110000",
64244 => "0111111111110000",
64245 => "0111111111110000",
64246 => "0111111111110000",
64247 => "0111111111110000",
64248 => "0111111111110000",
64249 => "0111111111110000",
64250 => "0111111111110000",
64251 => "0111111111110000",
64252 => "0111111111110000",
64253 => "0111111111110000",
64254 => "0111111111110000",
64255 => "0111111111110000",
64256 => "0111111111110000",
64257 => "0111111111110000",
64258 => "0111111111110000",
64259 => "0111111111110000",
64260 => "0111111111110000",
64261 => "0111111111110000",
64262 => "0111111111110000",
64263 => "0111111111110000",
64264 => "0111111111110000",
64265 => "0111111111110000",
64266 => "0111111111110000",
64267 => "0111111111110000",
64268 => "0111111111110000",
64269 => "0111111111110000",
64270 => "0111111111110000",
64271 => "0111111111110000",
64272 => "0111111111110000",
64273 => "0111111111110000",
64274 => "0111111111110000",
64275 => "0111111111110000",
64276 => "0111111111110000",
64277 => "0111111111110000",
64278 => "0111111111110000",
64279 => "0111111111110000",
64280 => "0111111111110000",
64281 => "0111111111110000",
64282 => "0111111111110000",
64283 => "0111111111110000",
64284 => "0111111111110000",
64285 => "0111111111110000",
64286 => "0111111111110000",
64287 => "0111111111110000",
64288 => "0111111111110000",
64289 => "0111111111110000",
64290 => "0111111111110000",
64291 => "0111111111110000",
64292 => "0111111111110000",
64293 => "0111111111110000",
64294 => "0111111111110000",
64295 => "0111111111110000",
64296 => "0111111111110000",
64297 => "0111111111110000",
64298 => "0111111111110000",
64299 => "0111111111110000",
64300 => "0111111111110000",
64301 => "0111111111110000",
64302 => "0111111111110000",
64303 => "0111111111110000",
64304 => "0111111111110000",
64305 => "0111111111110000",
64306 => "0111111111110000",
64307 => "0111111111110000",
64308 => "0111111111110000",
64309 => "0111111111110000",
64310 => "0111111111110000",
64311 => "0111111111110000",
64312 => "0111111111110000",
64313 => "0111111111110000",
64314 => "0111111111110000",
64315 => "0111111111110000",
64316 => "0111111111110000",
64317 => "0111111111110000",
64318 => "0111111111110000",
64319 => "0111111111110000",
64320 => "0111111111110000",
64321 => "0111111111110000",
64322 => "0111111111110000",
64323 => "0111111111110000",
64324 => "0111111111110000",
64325 => "0111111111110000",
64326 => "0111111111110000",
64327 => "0111111111110000",
64328 => "0111111111110000",
64329 => "0111111111110000",
64330 => "0111111111110000",
64331 => "0111111111110000",
64332 => "0111111111110000",
64333 => "0111111111110000",
64334 => "0111111111110000",
64335 => "0111111111110000",
64336 => "0111111111110000",
64337 => "0111111111110000",
64338 => "0111111111110000",
64339 => "0111111111110000",
64340 => "0111111111110000",
64341 => "0111111111110000",
64342 => "0111111111110000",
64343 => "0111111111110000",
64344 => "0111111111110000",
64345 => "0111111111110000",
64346 => "0111111111110000",
64347 => "0111111111110000",
64348 => "0111111111110000",
64349 => "0111111111110000",
64350 => "0111111111110000",
64351 => "0111111111110000",
64352 => "0111111111110000",
64353 => "0111111111110000",
64354 => "0111111111110000",
64355 => "0111111111110000",
64356 => "0111111111110000",
64357 => "0111111111110000",
64358 => "0111111111110000",
64359 => "0111111111110000",
64360 => "0111111111110000",
64361 => "0111111111110000",
64362 => "0111111111110000",
64363 => "0111111111110000",
64364 => "0111111111110000",
64365 => "0111111111110000",
64366 => "0111111111110000",
64367 => "0111111111110000",
64368 => "0111111111110000",
64369 => "0111111111110000",
64370 => "0111111111110000",
64371 => "0111111111110000",
64372 => "0111111111110000",
64373 => "0111111111110000",
64374 => "0111111111110000",
64375 => "0111111111110000",
64376 => "0111111111110000",
64377 => "0111111111110000",
64378 => "0111111111110000",
64379 => "0111111111110000",
64380 => "0111111111110000",
64381 => "0111111111110000",
64382 => "0111111111110000",
64383 => "0111111111110000",
64384 => "0111111111110000",
64385 => "0111111111110000",
64386 => "0111111111110000",
64387 => "0111111111110000",
64388 => "0111111111110000",
64389 => "0111111111110000",
64390 => "0111111111110000",
64391 => "0111111111110000",
64392 => "0111111111110000",
64393 => "0111111111110000",
64394 => "0111111111110000",
64395 => "0111111111110000",
64396 => "0111111111110000",
64397 => "0111111111110000",
64398 => "0111111111110000",
64399 => "0111111111110000",
64400 => "0111111111110000",
64401 => "0111111111110000",
64402 => "0111111111110000",
64403 => "0111111111110000",
64404 => "0111111111110000",
64405 => "0111111111110000",
64406 => "0111111111110000",
64407 => "0111111111110000",
64408 => "0111111111110000",
64409 => "0111111111110000",
64410 => "0111111111110000",
64411 => "0111111111110000",
64412 => "0111111111110000",
64413 => "0111111111110000",
64414 => "0111111111110000",
64415 => "0111111111110000",
64416 => "0111111111110000",
64417 => "0111111111110000",
64418 => "0111111111110000",
64419 => "0111111111110000",
64420 => "0111111111110000",
64421 => "0111111111110000",
64422 => "0111111111110000",
64423 => "0111111111110000",
64424 => "0111111111110000",
64425 => "0111111111110000",
64426 => "0111111111110000",
64427 => "0111111111110000",
64428 => "0111111111110000",
64429 => "0111111111110000",
64430 => "0111111111110000",
64431 => "0111111111110000",
64432 => "0111111111110000",
64433 => "0111111111110000",
64434 => "0111111111110000",
64435 => "0111111111110000",
64436 => "0111111111110000",
64437 => "0111111111110000",
64438 => "0111111111110000",
64439 => "0111111111110000",
64440 => "0111111111110000",
64441 => "0111111111110000",
64442 => "0111111111110000",
64443 => "0111111111110000",
64444 => "0111111111110000",
64445 => "0111111111110000",
64446 => "0111111111110000",
64447 => "0111111111110000",
64448 => "0111111111110000",
64449 => "0111111111110000",
64450 => "0111111111110000",
64451 => "0111111111110000",
64452 => "0111111111110000",
64453 => "0111111111110000",
64454 => "0111111111110000",
64455 => "0111111111110000",
64456 => "0111111111110000",
64457 => "0111111111110000",
64458 => "0111111111110000",
64459 => "0111111111110000",
64460 => "0111111111110000",
64461 => "0111111111110000",
64462 => "0111111111110000",
64463 => "0111111111110000",
64464 => "0111111111110000",
64465 => "0111111111110000",
64466 => "0111111111110000",
64467 => "0111111111110000",
64468 => "0111111111110000",
64469 => "0111111111110000",
64470 => "0111111111110000",
64471 => "0111111111110000",
64472 => "0111111111110000",
64473 => "0111111111110000",
64474 => "0111111111110000",
64475 => "0111111111110000",
64476 => "0111111111110000",
64477 => "0111111111110000",
64478 => "0111111111110000",
64479 => "0111111111110000",
64480 => "0111111111110000",
64481 => "0111111111110000",
64482 => "0111111111110000",
64483 => "0111111111110000",
64484 => "0111111111110000",
64485 => "0111111111110000",
64486 => "0111111111110000",
64487 => "0111111111110000",
64488 => "0111111111110000",
64489 => "0111111111110000",
64490 => "0111111111110000",
64491 => "0111111111110000",
64492 => "0111111111110000",
64493 => "0111111111110000",
64494 => "0111111111110000",
64495 => "0111111111110000",
64496 => "0111111111110000",
64497 => "0111111111110000",
64498 => "0111111111110000",
64499 => "0111111111110000",
64500 => "0111111111110000",
64501 => "0111111111110000",
64502 => "0111111111110000",
64503 => "0111111111110000",
64504 => "0111111111110000",
64505 => "0111111111110000",
64506 => "0111111111110000",
64507 => "0111111111110000",
64508 => "0111111111110000",
64509 => "0111111111110000",
64510 => "0111111111110000",
64511 => "0111111111110000",
64512 => "0111111111110000",
64513 => "0111111111110000",
64514 => "0111111111110000",
64515 => "0111111111110000",
64516 => "0111111111110000",
64517 => "0111111111110000",
64518 => "0111111111110000",
64519 => "0111111111110000",
64520 => "0111111111110000",
64521 => "0111111111110000",
64522 => "0111111111110000",
64523 => "0111111111110000",
64524 => "0111111111110000",
64525 => "0111111111110000",
64526 => "0111111111110000",
64527 => "0111111111110000",
64528 => "0111111111110000",
64529 => "0111111111110000",
64530 => "0111111111110000",
64531 => "0111111111110000",
64532 => "0111111111110000",
64533 => "0111111111110000",
64534 => "0111111111110000",
64535 => "0111111111110000",
64536 => "0111111111110000",
64537 => "0111111111110000",
64538 => "0111111111110000",
64539 => "0111111111110000",
64540 => "0111111111110000",
64541 => "0111111111110000",
64542 => "0111111111110000",
64543 => "0111111111110000",
64544 => "0111111111110000",
64545 => "0111111111110000",
64546 => "0111111111110000",
64547 => "0111111111110000",
64548 => "0111111111110000",
64549 => "0111111111110000",
64550 => "0111111111110000",
64551 => "0111111111110000",
64552 => "0111111111110000",
64553 => "0111111111110000",
64554 => "0111111111110000",
64555 => "0111111111110000",
64556 => "0111111111110000",
64557 => "0111111111110000",
64558 => "0111111111110000",
64559 => "0111111111110000",
64560 => "0111111111110000",
64561 => "0111111111110000",
64562 => "0111111111110000",
64563 => "0111111111110000",
64564 => "0111111111110000",
64565 => "0111111111110000",
64566 => "0111111111110000",
64567 => "0111111111110000",
64568 => "0111111111110000",
64569 => "0111111111110000",
64570 => "0111111111110000",
64571 => "0111111111110000",
64572 => "0111111111110000",
64573 => "0111111111110000",
64574 => "0111111111110000",
64575 => "0111111111110000",
64576 => "0111111111110000",
64577 => "0111111111110000",
64578 => "0111111111110000",
64579 => "0111111111110000",
64580 => "0111111111110000",
64581 => "0111111111110000",
64582 => "0111111111110000",
64583 => "0111111111110000",
64584 => "0111111111110000",
64585 => "0111111111110000",
64586 => "0111111111110000",
64587 => "0111111111110000",
64588 => "0111111111110000",
64589 => "0111111111110000",
64590 => "0111111111110000",
64591 => "0111111111110000",
64592 => "0111111111110000",
64593 => "0111111111110000",
64594 => "0111111111110000",
64595 => "0111111111110000",
64596 => "0111111111110000",
64597 => "0111111111110000",
64598 => "0111111111110000",
64599 => "0111111111110000",
64600 => "0111111111110000",
64601 => "0111111111110000",
64602 => "0111111111110000",
64603 => "0111111111110000",
64604 => "0111111111110000",
64605 => "0111111111110000",
64606 => "0111111111110000",
64607 => "0111111111110000",
64608 => "0111111111110000",
64609 => "0111111111110000",
64610 => "0111111111110000",
64611 => "0111111111110000",
64612 => "0111111111110000",
64613 => "0111111111110000",
64614 => "0111111111110000",
64615 => "0111111111110000",
64616 => "0111111111110000",
64617 => "0111111111110000",
64618 => "0111111111110000",
64619 => "0111111111110000",
64620 => "0111111111110000",
64621 => "0111111111110000",
64622 => "0111111111110000",
64623 => "0111111111110000",
64624 => "0111111111110000",
64625 => "0111111111110000",
64626 => "0111111111110000",
64627 => "0111111111110000",
64628 => "0111111111110000",
64629 => "0111111111110000",
64630 => "0111111111110000",
64631 => "0111111111110000",
64632 => "0111111111110000",
64633 => "0111111111110000",
64634 => "0111111111110000",
64635 => "0111111111110000",
64636 => "0111111111110000",
64637 => "0111111111110000",
64638 => "0111111111110000",
64639 => "0111111111110000",
64640 => "0111111111110000",
64641 => "0111111111110000",
64642 => "0111111111110000",
64643 => "0111111111110000",
64644 => "0111111111110000",
64645 => "0111111111110000",
64646 => "0111111111110000",
64647 => "0111111111110000",
64648 => "0111111111110000",
64649 => "0111111111110000",
64650 => "0111111111110000",
64651 => "0111111111110000",
64652 => "0111111111110000",
64653 => "0111111111110000",
64654 => "0111111111110000",
64655 => "0111111111110000",
64656 => "0111111111110000",
64657 => "0111111111110000",
64658 => "0111111111110000",
64659 => "0111111111110000",
64660 => "0111111111110000",
64661 => "0111111111110000",
64662 => "0111111111110000",
64663 => "0111111111110000",
64664 => "0111111111110000",
64665 => "0111111111110000",
64666 => "0111111111110000",
64667 => "0111111111110000",
64668 => "0111111111110000",
64669 => "0111111111110000",
64670 => "0111111111110000",
64671 => "0111111111110000",
64672 => "0111111111110000",
64673 => "0111111111110000",
64674 => "0111111111110000",
64675 => "0111111111110000",
64676 => "0111111111110000",
64677 => "0111111111110000",
64678 => "0111111111110000",
64679 => "0111111111110000",
64680 => "0111111111110000",
64681 => "0111111111110000",
64682 => "0111111111110000",
64683 => "0111111111110000",
64684 => "0111111111110000",
64685 => "0111111111110000",
64686 => "0111111111110000",
64687 => "0111111111110000",
64688 => "0111111111110000",
64689 => "0111111111110000",
64690 => "0111111111110000",
64691 => "0111111111110000",
64692 => "0111111111110000",
64693 => "0111111111110000",
64694 => "0111111111110000",
64695 => "0111111111110000",
64696 => "0111111111110000",
64697 => "0111111111110000",
64698 => "0111111111110000",
64699 => "0111111111110000",
64700 => "0111111111110000",
64701 => "0111111111110000",
64702 => "0111111111110000",
64703 => "0111111111110000",
64704 => "0111111111110000",
64705 => "0111111111110000",
64706 => "0111111111110000",
64707 => "0111111111110000",
64708 => "0111111111110000",
64709 => "0111111111110000",
64710 => "0111111111110000",
64711 => "0111111111110000",
64712 => "0111111111110000",
64713 => "0111111111110000",
64714 => "0111111111110000",
64715 => "0111111111110000",
64716 => "0111111111110000",
64717 => "0111111111110000",
64718 => "0111111111110000",
64719 => "0111111111110000",
64720 => "0111111111110000",
64721 => "0111111111110000",
64722 => "0111111111110000",
64723 => "0111111111110000",
64724 => "0111111111110000",
64725 => "0111111111110000",
64726 => "0111111111110000",
64727 => "0111111111110000",
64728 => "0111111111110000",
64729 => "0111111111110000",
64730 => "0111111111110000",
64731 => "0111111111110000",
64732 => "0111111111110000",
64733 => "0111111111110000",
64734 => "0111111111110000",
64735 => "0111111111110000",
64736 => "0111111111110000",
64737 => "0111111111110000",
64738 => "0111111111110000",
64739 => "0111111111110000",
64740 => "0111111111110000",
64741 => "0111111111110000",
64742 => "0111111111110000",
64743 => "0111111111110000",
64744 => "0111111111110000",
64745 => "0111111111110000",
64746 => "0111111111110000",
64747 => "0111111111110000",
64748 => "0111111111110000",
64749 => "0111111111110000",
64750 => "0111111111110000",
64751 => "0111111111110000",
64752 => "0111111111110000",
64753 => "0111111111110000",
64754 => "0111111111110000",
64755 => "0111111111110000",
64756 => "0111111111110000",
64757 => "0111111111110000",
64758 => "0111111111110000",
64759 => "0111111111110000",
64760 => "0111111111110000",
64761 => "0111111111110000",
64762 => "0111111111110000",
64763 => "0111111111110000",
64764 => "0111111111110000",
64765 => "0111111111110000",
64766 => "0111111111110000",
64767 => "0111111111110000",
64768 => "0111111111110000",
64769 => "0111111111110000",
64770 => "0111111111110000",
64771 => "0111111111110000",
64772 => "0111111111110000",
64773 => "0111111111110000",
64774 => "0111111111110000",
64775 => "0111111111110000",
64776 => "0111111111110000",
64777 => "0111111111110000",
64778 => "0111111111110000",
64779 => "0111111111110000",
64780 => "0111111111110000",
64781 => "0111111111110000",
64782 => "0111111111110000",
64783 => "0111111111110000",
64784 => "0111111111110000",
64785 => "0111111111110000",
64786 => "0111111111110000",
64787 => "0111111111110000",
64788 => "0111111111110000",
64789 => "0111111111110000",
64790 => "0111111111110000",
64791 => "0111111111110000",
64792 => "0111111111110000",
64793 => "0111111111110000",
64794 => "0111111111110000",
64795 => "0111111111110000",
64796 => "0111111111110000",
64797 => "0111111111110000",
64798 => "0111111111110000",
64799 => "0111111111110000",
64800 => "0111111111110000",
64801 => "0111111111110000",
64802 => "0111111111110000",
64803 => "0111111111110000",
64804 => "0111111111110000",
64805 => "0111111111110000",
64806 => "0111111111110000",
64807 => "0111111111110000",
64808 => "0111111111110000",
64809 => "0111111111110000",
64810 => "0111111111110000",
64811 => "0111111111110000",
64812 => "0111111111110000",
64813 => "0111111111110000",
64814 => "0111111111110000",
64815 => "0111111111110000",
64816 => "0111111111110000",
64817 => "0111111111110000",
64818 => "0111111111110000",
64819 => "0111111111110000",
64820 => "0111111111110000",
64821 => "0111111111110000",
64822 => "0111111111110000",
64823 => "0111111111110000",
64824 => "0111111111110000",
64825 => "0111111111110000",
64826 => "0111111111110000",
64827 => "0111111111110000",
64828 => "0111111111110000",
64829 => "0111111111110000",
64830 => "0111111111110000",
64831 => "0111111111110000",
64832 => "0111111111110000",
64833 => "0111111111110000",
64834 => "0111111111110000",
64835 => "0111111111110000",
64836 => "0111111111110000",
64837 => "0111111111110000",
64838 => "0111111111110000",
64839 => "0111111111110000",
64840 => "0111111111110000",
64841 => "0111111111110000",
64842 => "0111111111110000",
64843 => "0111111111110000",
64844 => "0111111111110000",
64845 => "0111111111110000",
64846 => "0111111111110000",
64847 => "0111111111110000",
64848 => "0111111111110000",
64849 => "0111111111110000",
64850 => "0111111111110000",
64851 => "0111111111110000",
64852 => "0111111111110000",
64853 => "0111111111110000",
64854 => "0111111111110000",
64855 => "0111111111110000",
64856 => "0111111111110000",
64857 => "0111111111110000",
64858 => "0111111111110000",
64859 => "0111111111110000",
64860 => "0111111111110000",
64861 => "0111111111110000",
64862 => "0111111111110000",
64863 => "0111111111110000",
64864 => "0111111111110000",
64865 => "0111111111110000",
64866 => "0111111111110000",
64867 => "0111111111110000",
64868 => "0111111111110000",
64869 => "0111111111110000",
64870 => "0111111111110000",
64871 => "0111111111110000",
64872 => "0111111111110000",
64873 => "0111111111110000",
64874 => "0111111111110000",
64875 => "0111111111110000",
64876 => "0111111111110000",
64877 => "0111111111110000",
64878 => "0111111111110000",
64879 => "0111111111110000",
64880 => "0111111111110000",
64881 => "0111111111110000",
64882 => "0111111111110000",
64883 => "0111111111110000",
64884 => "0111111111110000",
64885 => "0111111111110000",
64886 => "0111111111110000",
64887 => "0111111111110000",
64888 => "0111111111110000",
64889 => "0111111111110000",
64890 => "0111111111110000",
64891 => "0111111111110000",
64892 => "0111111111110000",
64893 => "0111111111110000",
64894 => "0111111111110000",
64895 => "0111111111110000",
64896 => "0111111111110000",
64897 => "0111111111110000",
64898 => "0111111111110000",
64899 => "0111111111110000",
64900 => "0111111111110000",
64901 => "0111111111110000",
64902 => "0111111111110000",
64903 => "0111111111110000",
64904 => "0111111111110000",
64905 => "0111111111110000",
64906 => "0111111111110000",
64907 => "0111111111110000",
64908 => "0111111111110000",
64909 => "0111111111110000",
64910 => "0111111111110000",
64911 => "0111111111110000",
64912 => "0111111111110000",
64913 => "0111111111110000",
64914 => "0111111111110000",
64915 => "0111111111110000",
64916 => "0111111111110000",
64917 => "0111111111110000",
64918 => "0111111111110000",
64919 => "0111111111110000",
64920 => "0111111111110000",
64921 => "0111111111110000",
64922 => "0111111111110000",
64923 => "0111111111110000",
64924 => "0111111111110000",
64925 => "0111111111110000",
64926 => "0111111111110000",
64927 => "0111111111110000",
64928 => "0111111111110000",
64929 => "0111111111110000",
64930 => "0111111111110000",
64931 => "0111111111110000",
64932 => "0111111111110000",
64933 => "0111111111110000",
64934 => "0111111111110000",
64935 => "0111111111110000",
64936 => "0111111111110000",
64937 => "0111111111110000",
64938 => "0111111111110000",
64939 => "0111111111110000",
64940 => "0111111111110000",
64941 => "0111111111110000",
64942 => "0111111111110000",
64943 => "0111111111110000",
64944 => "0111111111110000",
64945 => "0111111111110000",
64946 => "0111111111110000",
64947 => "0111111111110000",
64948 => "0111111111110000",
64949 => "0111111111110000",
64950 => "0111111111110000",
64951 => "0111111111110000",
64952 => "0111111111110000",
64953 => "0111111111110000",
64954 => "0111111111110000",
64955 => "0111111111110000",
64956 => "0111111111110000",
64957 => "0111111111110000",
64958 => "0111111111110000",
64959 => "0111111111110000",
64960 => "0111111111110000",
64961 => "0111111111110000",
64962 => "0111111111110000",
64963 => "0111111111110000",
64964 => "0111111111110000",
64965 => "0111111111110000",
64966 => "0111111111110000",
64967 => "0111111111110000",
64968 => "0111111111110000",
64969 => "0111111111110000",
64970 => "0111111111110000",
64971 => "0111111111110000",
64972 => "0111111111110000",
64973 => "0111111111110000",
64974 => "0111111111110000",
64975 => "0111111111110000",
64976 => "0111111111110000",
64977 => "0111111111110000",
64978 => "0111111111110000",
64979 => "0111111111110000",
64980 => "0111111111110000",
64981 => "0111111111110000",
64982 => "0111111111110000",
64983 => "0111111111110000",
64984 => "0111111111110000",
64985 => "0111111111110000",
64986 => "0111111111110000",
64987 => "0111111111110000",
64988 => "0111111111110000",
64989 => "0111111111110000",
64990 => "0111111111110000",
64991 => "0111111111110000",
64992 => "0111111111110000",
64993 => "0111111111110000",
64994 => "0111111111110000",
64995 => "0111111111110000",
64996 => "0111111111110000",
64997 => "0111111111110000",
64998 => "0111111111110000",
64999 => "0111111111110000",
65000 => "0111111111110000",
65001 => "0111111111110000",
65002 => "0111111111110000",
65003 => "0111111111110000",
65004 => "0111111111110000",
65005 => "0111111111110000",
65006 => "0111111111110000",
65007 => "0111111111110000",
65008 => "0111111111110000",
65009 => "0111111111110000",
65010 => "0111111111110000",
65011 => "0111111111110000",
65012 => "0111111111110000",
65013 => "0111111111110000",
65014 => "0111111111110000",
65015 => "0111111111110000",
65016 => "0111111111110000",
65017 => "0111111111110000",
65018 => "0111111111110000",
65019 => "0111111111110000",
65020 => "0111111111110000",
65021 => "0111111111110000",
65022 => "0111111111110000",
65023 => "0111111111110000",
65024 => "0111111111110000",
65025 => "0111111111110000",
65026 => "0111111111110000",
65027 => "0111111111110000",
65028 => "0111111111110000",
65029 => "0111111111110000",
65030 => "0111111111110000",
65031 => "0111111111110000",
65032 => "0111111111110000",
65033 => "0111111111110000",
65034 => "0111111111110000",
65035 => "0111111111110000",
65036 => "0111111111110000",
65037 => "0111111111110000",
65038 => "0111111111110000",
65039 => "0111111111110000",
65040 => "0111111111110000",
65041 => "0111111111110000",
65042 => "0111111111110000",
65043 => "0111111111110000",
65044 => "0111111111110000",
65045 => "0111111111110000",
65046 => "0111111111110000",
65047 => "0111111111110000",
65048 => "0111111111110000",
65049 => "0111111111110000",
65050 => "0111111111110000",
65051 => "0111111111110000",
65052 => "0111111111110000",
65053 => "0111111111110000",
65054 => "0111111111110000",
65055 => "0111111111110000",
65056 => "0111111111110000",
65057 => "0111111111110000",
65058 => "0111111111110000",
65059 => "0111111111110000",
65060 => "0111111111110000",
65061 => "0111111111110000",
65062 => "0111111111110000",
65063 => "0111111111110000",
65064 => "0111111111110000",
65065 => "0111111111110000",
65066 => "0111111111110000",
65067 => "0111111111110000",
65068 => "0111111111110000",
65069 => "0111111111110000",
65070 => "0111111111110000",
65071 => "0111111111110000",
65072 => "0111111111110000",
65073 => "0111111111110000",
65074 => "0111111111110000",
65075 => "0111111111110000",
65076 => "0111111111110000",
65077 => "0111111111110000",
65078 => "0111111111110000",
65079 => "0111111111110000",
65080 => "0111111111110000",
65081 => "0111111111110000",
65082 => "0111111111110000",
65083 => "0111111111110000",
65084 => "0111111111110000",
65085 => "0111111111110000",
65086 => "0111111111110000",
65087 => "0111111111110000",
65088 => "0111111111110000",
65089 => "0111111111110000",
65090 => "0111111111110000",
65091 => "0111111111110000",
65092 => "0111111111110000",
65093 => "0111111111110000",
65094 => "0111111111110000",
65095 => "0111111111110000",
65096 => "0111111111110000",
65097 => "0111111111110000",
65098 => "0111111111110000",
65099 => "0111111111110000",
65100 => "0111111111110000",
65101 => "0111111111110000",
65102 => "0111111111110000",
65103 => "0111111111110000",
65104 => "0111111111110000",
65105 => "0111111111110000",
65106 => "0111111111110000",
65107 => "0111111111110000",
65108 => "0111111111110000",
65109 => "0111111111110000",
65110 => "0111111111110000",
65111 => "0111111111110000",
65112 => "0111111111110000",
65113 => "0111111111110000",
65114 => "0111111111110000",
65115 => "0111111111110000",
65116 => "0111111111110000",
65117 => "0111111111110000",
65118 => "0111111111110000",
65119 => "0111111111110000",
65120 => "0111111111110000",
65121 => "0111111111110000",
65122 => "0111111111110000",
65123 => "0111111111110000",
65124 => "0111111111110000",
65125 => "0111111111110000",
65126 => "0111111111110000",
65127 => "0111111111110000",
65128 => "0111111111110000",
65129 => "0111111111110000",
65130 => "0111111111110000",
65131 => "0111111111110000",
65132 => "0111111111110000",
65133 => "0111111111110000",
65134 => "0111111111110000",
65135 => "0111111111110000",
65136 => "0111111111110000",
65137 => "0111111111110000",
65138 => "0111111111110000",
65139 => "0111111111110000",
65140 => "0111111111110000",
65141 => "0111111111110000",
65142 => "0111111111110000",
65143 => "0111111111110000",
65144 => "0111111111110000",
65145 => "0111111111110000",
65146 => "0111111111110000",
65147 => "0111111111110000",
65148 => "0111111111110000",
65149 => "0111111111110000",
65150 => "0111111111110000",
65151 => "0111111111110000",
65152 => "0111111111110000",
65153 => "0111111111110000",
65154 => "0111111111110000",
65155 => "0111111111110000",
65156 => "0111111111110000",
65157 => "0111111111110000",
65158 => "0111111111110000",
65159 => "0111111111110000",
65160 => "0111111111110000",
65161 => "0111111111110000",
65162 => "0111111111110000",
65163 => "0111111111110000",
65164 => "0111111111110000",
65165 => "0111111111110000",
65166 => "0111111111110000",
65167 => "0111111111110000",
65168 => "0111111111110000",
65169 => "0111111111110000",
65170 => "0111111111110000",
65171 => "0111111111110000",
65172 => "0111111111110000",
65173 => "0111111111110000",
65174 => "0111111111110000",
65175 => "0111111111110000",
65176 => "0111111111110000",
65177 => "0111111111110000",
65178 => "0111111111110000",
65179 => "0111111111110000",
65180 => "0111111111110000",
65181 => "0111111111110000",
65182 => "0111111111110000",
65183 => "0111111111110000",
65184 => "0111111111110000",
65185 => "0111111111110000",
65186 => "0111111111110000",
65187 => "0111111111110000",
65188 => "0111111111110000",
65189 => "0111111111110000",
65190 => "0111111111110000",
65191 => "0111111111110000",
65192 => "0111111111110000",
65193 => "0111111111110000",
65194 => "0111111111110000",
65195 => "0111111111110000",
65196 => "0111111111110000",
65197 => "0111111111110000",
65198 => "0111111111110000",
65199 => "0111111111110000",
65200 => "0111111111110000",
65201 => "0111111111110000",
65202 => "0111111111110000",
65203 => "0111111111110000",
65204 => "0111111111110000",
65205 => "0111111111110000",
65206 => "0111111111110000",
65207 => "0111111111110000",
65208 => "0111111111110000",
65209 => "0111111111110000",
65210 => "0111111111110000",
65211 => "0111111111110000",
65212 => "0111111111110000",
65213 => "0111111111110000",
65214 => "0111111111110000",
65215 => "0111111111110000",
65216 => "0111111111110000",
65217 => "0111111111110000",
65218 => "0111111111110000",
65219 => "0111111111110000",
65220 => "0111111111110000",
65221 => "0111111111110000",
65222 => "0111111111110000",
65223 => "0111111111110000",
65224 => "0111111111110000",
65225 => "0111111111110000",
65226 => "0111111111110000",
65227 => "0111111111110000",
65228 => "0111111111110000",
65229 => "0111111111110000",
65230 => "0111111111110000",
65231 => "0111111111110000",
65232 => "0111111111110000",
65233 => "0111111111110000",
65234 => "0111111111110000",
65235 => "0111111111110000",
65236 => "0111111111110000",
65237 => "0111111111110000",
65238 => "0111111111110000",
65239 => "0111111111110000",
65240 => "0111111111110000",
65241 => "0111111111110000",
65242 => "0111111111110000",
65243 => "0111111111110000",
65244 => "0111111111110000",
65245 => "0111111111110000",
65246 => "0111111111110000",
65247 => "0111111111110000",
65248 => "0111111111110000",
65249 => "0111111111110000",
65250 => "0111111111110000",
65251 => "0111111111110000",
65252 => "0111111111110000",
65253 => "0111111111110000",
65254 => "0111111111110000",
65255 => "0111111111110000",
65256 => "0111111111110000",
65257 => "0111111111110000",
65258 => "0111111111110000",
65259 => "0111111111110000",
65260 => "0111111111110000",
65261 => "0111111111110000",
65262 => "0111111111110000",
65263 => "0111111111110000",
65264 => "0111111111110000",
65265 => "0111111111110000",
65266 => "0111111111110000",
65267 => "0111111111110000",
65268 => "0111111111110000",
65269 => "0111111111110000",
65270 => "0111111111110000",
65271 => "0111111111110000",
65272 => "0111111111110000",
65273 => "0111111111110000",
65274 => "0111111111110000",
65275 => "0111111111110000",
65276 => "0111111111110000",
65277 => "0111111111110000",
65278 => "0111111111110000",
65279 => "0111111111110000",
65280 => "0111111111110000",
65281 => "0111111111110000",
65282 => "0111111111110000",
65283 => "0111111111110000",
65284 => "0111111111110000",
65285 => "0111111111110000",
65286 => "0111111111110000",
65287 => "0111111111110000",
65288 => "0111111111110000",
65289 => "0111111111110000",
65290 => "0111111111110000",
65291 => "0111111111110000",
65292 => "0111111111110000",
65293 => "0111111111110000",
65294 => "0111111111110000",
65295 => "0111111111110000",
65296 => "0111111111110000",
65297 => "0111111111110000",
65298 => "0111111111110000",
65299 => "0111111111110000",
65300 => "0111111111110000",
65301 => "0111111111110000",
65302 => "0111111111110000",
65303 => "0111111111110000",
65304 => "0111111111110000",
65305 => "0111111111110000",
65306 => "0111111111110000",
65307 => "0111111111110000",
65308 => "0111111111110000",
65309 => "0111111111110000",
65310 => "0111111111110000",
65311 => "0111111111110000",
65312 => "0111111111110000",
65313 => "0111111111110000",
65314 => "0111111111110000",
65315 => "0111111111110000",
65316 => "0111111111110000",
65317 => "0111111111110000",
65318 => "0111111111110000",
65319 => "0111111111110000",
65320 => "0111111111110000",
65321 => "0111111111110000",
65322 => "0111111111110000",
65323 => "0111111111110000",
65324 => "0111111111110000",
65325 => "0111111111110000",
65326 => "0111111111110000",
65327 => "0111111111110000",
65328 => "0111111111110000",
65329 => "0111111111110000",
65330 => "0111111111110000",
65331 => "0111111111110000",
65332 => "0111111111110000",
65333 => "0111111111110000",
65334 => "0111111111110000",
65335 => "0111111111110000",
65336 => "0111111111110000",
65337 => "0111111111110000",
65338 => "0111111111110000",
65339 => "0111111111110000",
65340 => "0111111111110000",
65341 => "0111111111110000",
65342 => "0111111111110000",
65343 => "0111111111110000",
65344 => "0111111111110000",
65345 => "0111111111110000",
65346 => "0111111111110000",
65347 => "0111111111110000",
65348 => "0111111111110000",
65349 => "0111111111110000",
65350 => "0111111111110000",
65351 => "0111111111110000",
65352 => "0111111111110000",
65353 => "0111111111110000",
65354 => "0111111111110000",
65355 => "0111111111110000",
65356 => "0111111111110000",
65357 => "0111111111110000",
65358 => "0111111111110000",
65359 => "0111111111110000",
65360 => "0111111111110000",
65361 => "0111111111110000",
65362 => "0111111111110000",
65363 => "0111111111110000",
65364 => "0111111111110000",
65365 => "0111111111110000",
65366 => "0111111111110000",
65367 => "0111111111110000",
65368 => "0111111111110000",
65369 => "0111111111110000",
65370 => "0111111111110000",
65371 => "0111111111110000",
65372 => "0111111111110000",
65373 => "0111111111110000",
65374 => "0111111111110000",
65375 => "0111111111110000",
65376 => "0111111111110000",
65377 => "0111111111110000",
65378 => "0111111111110000",
65379 => "0111111111110000",
65380 => "0111111111110000",
65381 => "0111111111110000",
65382 => "0111111111110000",
65383 => "0111111111110000",
65384 => "0111111111110000",
65385 => "0111111111110000",
65386 => "0111111111110000",
65387 => "0111111111110000",
65388 => "0111111111110000",
65389 => "0111111111110000",
65390 => "0111111111110000",
65391 => "0111111111110000",
65392 => "0111111111110000",
65393 => "0111111111110000",
65394 => "0111111111110000",
65395 => "0111111111110000",
65396 => "0111111111110000",
65397 => "0111111111110000",
65398 => "0111111111110000",
65399 => "0111111111110000",
65400 => "0111111111110000",
65401 => "0111111111110000",
65402 => "0111111111110000",
65403 => "0111111111110000",
65404 => "0111111111110000",
65405 => "0111111111110000",
65406 => "0111111111110000",
65407 => "0111111111110000",
65408 => "0111111111110000",
65409 => "0111111111110000",
65410 => "0111111111110000",
65411 => "0111111111110000",
65412 => "0111111111110000",
65413 => "0111111111110000",
65414 => "0111111111110000",
65415 => "0111111111110000",
65416 => "0111111111110000",
65417 => "0111111111110000",
65418 => "0111111111110000",
65419 => "0111111111110000",
65420 => "0111111111110000",
65421 => "0111111111110000",
65422 => "0111111111110000",
65423 => "0111111111110000",
65424 => "0111111111110000",
65425 => "0111111111110000",
65426 => "0111111111110000",
65427 => "0111111111110000",
65428 => "0111111111110000",
65429 => "0111111111110000",
65430 => "0111111111110000",
65431 => "0111111111110000",
65432 => "0111111111110000",
65433 => "0111111111110000",
65434 => "0111111111110000",
65435 => "0111111111110000",
65436 => "0111111111110000",
65437 => "0111111111110000",
65438 => "0111111111110000",
65439 => "0111111111110000",
65440 => "0111111111110000",
65441 => "0111111111110000",
65442 => "0111111111110000",
65443 => "0111111111110000",
65444 => "0111111111110000",
65445 => "0111111111110000",
65446 => "0111111111110000",
65447 => "0111111111110000",
65448 => "0111111111110000",
65449 => "0111111111110000",
65450 => "0111111111110000",
65451 => "0111111111110000",
65452 => "0111111111110000",
65453 => "0111111111110000",
65454 => "0111111111110000",
65455 => "0111111111110000",
65456 => "0111111111110000",
65457 => "0111111111110000",
65458 => "0111111111110000",
65459 => "0111111111110000",
65460 => "0111111111110000",
65461 => "0111111111110000",
65462 => "0111111111110000",
65463 => "0111111111110000",
65464 => "0111111111110000",
65465 => "0111111111110000",
65466 => "0111111111110000",
65467 => "0111111111110000",
65468 => "0111111111110000",
65469 => "0111111111110000",
65470 => "0111111111110000",
65471 => "0111111111110000",
65472 => "0111111111110000",
65473 => "0111111111110000",
65474 => "0111111111110000",
65475 => "0111111111110000",
65476 => "0111111111110000",
65477 => "0111111111110000",
65478 => "0111111111110000",
65479 => "0111111111110000",
65480 => "0111111111110000",
65481 => "0111111111110000",
65482 => "0111111111110000",
65483 => "0111111111110000",
65484 => "0111111111110000",
65485 => "0111111111110000",
65486 => "0111111111110000",
65487 => "0111111111110000",
65488 => "0111111111110000",
65489 => "0111111111110000",
65490 => "0111111111110000",
65491 => "0111111111110000",
65492 => "0111111111110000",
65493 => "0111111111110000",
65494 => "0111111111110000",
65495 => "0111111111110000",
65496 => "0111111111110000",
65497 => "0111111111110000",
65498 => "0111111111110000",
65499 => "0111111111110000",
65500 => "0111111111110000",
65501 => "0111111111110000",
65502 => "0111111111110000",
65503 => "0111111111110000",
65504 => "0111111111110000",
65505 => "0111111111110000",
65506 => "0111111111110000",
65507 => "0111111111110000",
65508 => "0111111111110000",
65509 => "0111111111110000",
65510 => "0111111111110000",
65511 => "0111111111110000",
65512 => "0111111111110000",
65513 => "0111111111110000",
65514 => "0111111111110000",
65515 => "0111111111110000",
65516 => "0111111111110000",
65517 => "0111111111110000",
65518 => "0111111111110000",
65519 => "0111111111110000",
65520 => "0111111111110000",
65521 => "0111111111110000",
65522 => "0111111111110000",
65523 => "0111111111110000",
65524 => "0111111111110000",
65525 => "0111111111110000",
65526 => "0111111111110000",
65527 => "0111111111110000",
65528 => "0111111111110000",
65529 => "0111111111110000",
65530 => "0111111111110000",
65531 => "0111111111110000",
65532 => "0111111111110000",
65533 => "0111111111110000",
65534 => "0111111111110000",
65535 => "0111111111110000"

	);

begin
	--data_reg <= lut_data(CounterLUT); -- LUT

-- receive
	receive_proc: process(clk)
	begin 
	if (rising_edge(clk)) then
		if (baudReceive_counter < 5208 ) then -- 9600 baud rate 
			baudReceive_counter <= baud_counter + 1;
		else
			baudReceive_counter <= 0;-- initialise counter again as reached max
			-- check if first bit is 0
			if (rx_counter = 0) then 
				if (rx = '0') then 
				rx_counter <= 1;
				end if;
			elsif (0 < rx_counter and rx_counter < 9) then 
				case (rx_counter) is 
					when 1 => rx_value(0) <= rx;
					when 2 => rx_value(1) <= rx;
					when 3 => rx_value(2) <= rx;
					when 4 => rx_value(3) <= rx;
					when 5 => rx_value(4) <= rx;
					when 6 => rx_value(5) <= rx;
					when 7 => rx_value(6) <= rx;
					when 8 => rx_value(7) <= rx;
					when others => rx_value(7) <= '0';
				end case;
				rx_counter <= rx_counter + 1; -- increment counter
			elsif (rx_counter = 9) then 
				if (rx = '1') then 
					rx_counter <= 0; -- reset the counter -- reached end of recieve
					if (rx_value = "01010011") then 
							flag_receive <= 1; -- S recived correct
					else
							flag_receive <= 0; -- S not recived correctly 
					end if;
				end if;
			end if;	
		end if;
	end if;
	end process receive_proc;
	
-- transmission 
	transmit_proc: process(flag_receive, clk, data_reg, CounterLUT) -- transmission
	begin
		data_reg <= lut_data(CounterLUT);
	if (CounterLUT < 65535) then
		if (rising_edge(clk)) then
			if (baud_counter < 5208 ) then -- 9600 baud rate 
				baud_counter <= baud_counter + 1;
			else
				tx <= '1'; -- assign 1 to tx to keep the line high (<= when assigning to an output pin)
				baud_counter <= 0;-- initialise counter again as reached max
				if (flag_receive = 1) then
					if (tx_counter = 0) then 
						tx <= '0'; -- start bit
						tx_counter <= 1;
					elsif (0 < tx_counter and tx_counter < 9) then
						case (tx_counter) is 
							when 1 => tx <= data_reg(0);
							when 2 => tx <= data_reg(1);
							when 3 => tx <= data_reg(2);
							when 4 => tx <= data_reg(3);
							when 5 => tx <= data_reg(4);
							when 6 => tx <= data_reg(5);
							when 7 => tx <= data_reg(6);
							when 8 => tx <= data_reg(7);
							when others => tx <= '0';
						end case;
						tx_counter <= tx_counter + 1;
					elsif (tx_counter = 9) then 
						tx <= '1'; -- stop bit
						tx_counter <= 10; -- reset counter need a reset somewhere but not sure
					elsif (tx_counter = 10) then 
						tx <= '0'; -- start bit of second byte
						tx_counter <= 11;
					elsif (10 < tx_counter and tx_counter < 19) then 
						case (tx_counter) is 
							when 11 => tx <= data_reg(8);
							when 12 => tx <= data_reg(9);
							when 13 => tx <= data_reg(10);
							when 14 => tx <= data_reg(11);
							when 15 => tx <= data_reg(12);
							when 16 => tx <= data_reg(13);
							when 17 => tx <= data_reg(14);
							when 18 => tx <= data_reg(15);
							when others => tx <= '0';
						end case;
						tx_counter <= tx_counter + 1;
					elsif(tx_counter = 19) then 
						tx <= '1'; -- stop bit
						tx_counter <= 0; -- reset counter
					end if;
				end if;
			end if;
		end if; 
		--CounterLUT <= CounterLUT + 1;
	end if;
	CounterLUT <= CounterLUT + 1;
	end process transmit_proc;
end UART;
